module ibex_core (alert_major_o,
    alert_minor_o,
    clk_i,
    core_sleep_o,
    data_err_i,
    data_gnt_i,
    data_req_o,
    data_rvalid_i,
    data_we_o,
    debug_req_i,
    fetch_enable_i,
    instr_err_i,
    instr_gnt_i,
    instr_req_o,
    instr_rvalid_i,
    irq_external_i,
    irq_nm_i,
    irq_software_i,
    irq_timer_i,
    rst_ni,
    test_en_i,
    boot_addr_i,
    data_addr_o,
    data_be_o,
    data_rdata_i,
    data_wdata_o,
    hart_id_i,
    instr_addr_o,
    instr_rdata_i,
    irq_fast_i);
 output alert_major_o;
 output alert_minor_o;
 input clk_i;
 output core_sleep_o;
 input data_err_i;
 input data_gnt_i;
 output data_req_o;
 input data_rvalid_i;
 output data_we_o;
 input debug_req_i;
 input fetch_enable_i;
 input instr_err_i;
 input instr_gnt_i;
 output instr_req_o;
 input instr_rvalid_i;
 input irq_external_i;
 input irq_nm_i;
 input irq_software_i;
 input irq_timer_i;
 input rst_ni;
 input test_en_i;
 input [31:0] boot_addr_i;
 output [31:0] data_addr_o;
 output [3:0] data_be_o;
 input [31:0] data_rdata_i;
 output [31:0] data_wdata_o;
 input [31:0] hart_id_i;
 output [31:0] instr_addr_o;
 input [31:0] instr_rdata_i;
 input [14:0] irq_fast_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire net1065;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire net1063;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire net1057;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire net1052;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire net1050;
 wire net1049;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire net1048;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire net1047;
 wire net1046;
 wire net1045;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire net1044;
 wire _05541_;
 wire _05542_;
 wire net1042;
 wire _05544_;
 wire net1041;
 wire net1040;
 wire net1039;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire net1038;
 wire _05560_;
 wire net1037;
 wire _05562_;
 wire net1036;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire net1035;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire net1034;
 wire _05584_;
 wire net1033;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire net1032;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire net1031;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire net1030;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire net1029;
 wire net1028;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire net1027;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire net1026;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire net1025;
 wire net1024;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire net1023;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire net1022;
 wire _05743_;
 wire net1021;
 wire _05745_;
 wire net1020;
 wire _05747_;
 wire net1019;
 wire net1018;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire net1017;
 wire _05755_;
 wire net1016;
 wire _05757_;
 wire net1015;
 wire net1014;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire net1013;
 wire _05781_;
 wire _05782_;
 wire net1012;
 wire net1011;
 wire net1010;
 wire _05786_;
 wire net1009;
 wire _05788_;
 wire net1008;
 wire _05790_;
 wire _05791_;
 wire net1007;
 wire net1006;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire net1005;
 wire _05798_;
 wire net1004;
 wire _05800_;
 wire net1003;
 wire _05802_;
 wire _05803_;
 wire net1002;
 wire net1001;
 wire _05806_;
 wire _05807_;
 wire net1000;
 wire net999;
 wire net998;
 wire _05811_;
 wire _05812_;
 wire net997;
 wire _05814_;
 wire _05815_;
 wire net996;
 wire net995;
 wire _05818_;
 wire _05819_;
 wire net994;
 wire _05821_;
 wire _05822_;
 wire net993;
 wire _05824_;
 wire _05825_;
 wire net992;
 wire _05827_;
 wire _05828_;
 wire net991;
 wire net990;
 wire _05831_;
 wire _05832_;
 wire net989;
 wire _05834_;
 wire _05835_;
 wire net988;
 wire net987;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire net986;
 wire _05842_;
 wire _05843_;
 wire net985;
 wire _05845_;
 wire _05846_;
 wire net984;
 wire net983;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire net982;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire net981;
 wire _05857_;
 wire _05858_;
 wire net980;
 wire net979;
 wire net978;
 wire _05862_;
 wire _05863_;
 wire net977;
 wire net976;
 wire _05866_;
 wire _05867_;
 wire net975;
 wire net974;
 wire _05870_;
 wire _05871_;
 wire net973;
 wire net972;
 wire _05874_;
 wire _05875_;
 wire net971;
 wire _05877_;
 wire _05878_;
 wire net970;
 wire net969;
 wire net968;
 wire _05882_;
 wire _05883_;
 wire net967;
 wire net966;
 wire net965;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire net964;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire net963;
 wire net962;
 wire net961;
 wire _05897_;
 wire _05898_;
 wire net960;
 wire _05900_;
 wire _05901_;
 wire net959;
 wire _05903_;
 wire _05904_;
 wire net958;
 wire net957;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire net956;
 wire net954;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire net953;
 wire net952;
 wire _05919_;
 wire _05920_;
 wire net951;
 wire net950;
 wire _05923_;
 wire _05924_;
 wire net949;
 wire net948;
 wire _05927_;
 wire _05928_;
 wire net947;
 wire _05930_;
 wire _05931_;
 wire net946;
 wire net945;
 wire net944;
 wire _05935_;
 wire _05936_;
 wire net943;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire net942;
 wire net941;
 wire net940;
 wire net939;
 wire net938;
 wire net937;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire net936;
 wire _06067_;
 wire _06068_;
 wire net935;
 wire _06070_;
 wire net934;
 wire _06072_;
 wire _06073_;
 wire net933;
 wire net932;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire net931;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire net930;
 wire _06087_;
 wire _06088_;
 wire net929;
 wire _06090_;
 wire _06091_;
 wire net928;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire net927;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire net926;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire net925;
 wire net924;
 wire net923;
 wire net922;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire net921;
 wire net920;
 wire _06257_;
 wire _06258_;
 wire net919;
 wire net918;
 wire net917;
 wire _06262_;
 wire net916;
 wire net915;
 wire net914;
 wire _06266_;
 wire net913;
 wire net912;
 wire net911;
 wire _06270_;
 wire _06271_;
 wire net910;
 wire net909;
 wire net908;
 wire _06275_;
 wire net907;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire net906;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire net905;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire net904;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire net903;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire net902;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire net901;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire net900;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire net899;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire net898;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire net897;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire net896;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire net895;
 wire _06528_;
 wire net894;
 wire net893;
 wire net892;
 wire _06532_;
 wire net891;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire net890;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire net889;
 wire net888;
 wire _06616_;
 wire _06617_;
 wire net887;
 wire _06619_;
 wire net886;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire net885;
 wire net884;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire net883;
 wire net882;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire net881;
 wire net880;
 wire _06669_;
 wire _06670_;
 wire net879;
 wire net878;
 wire _06673_;
 wire _06674_;
 wire net877;
 wire net876;
 wire _06677_;
 wire net875;
 wire net874;
 wire _06680_;
 wire _06681_;
 wire net873;
 wire _06683_;
 wire _06684_;
 wire net872;
 wire net871;
 wire net870;
 wire net869;
 wire net868;
 wire _06690_;
 wire net867;
 wire net866;
 wire net865;
 wire net864;
 wire _06695_;
 wire net863;
 wire _06697_;
 wire net862;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire net861;
 wire net860;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire net859;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire net858;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire net857;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire net856;
 wire net855;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire net854;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire net852;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire net851;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire net850;
 wire _06886_;
 wire net849;
 wire _06888_;
 wire _06889_;
 wire net848;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire net847;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire net846;
 wire net845;
 wire _06927_;
 wire _06928_;
 wire net844;
 wire net843;
 wire _06931_;
 wire _06932_;
 wire net842;
 wire _06934_;
 wire _06935_;
 wire net841;
 wire net840;
 wire _06938_;
 wire _06939_;
 wire net839;
 wire net838;
 wire _06942_;
 wire _06943_;
 wire net837;
 wire net836;
 wire _06946_;
 wire net835;
 wire _06948_;
 wire _06949_;
 wire net834;
 wire net833;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire net832;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire net831;
 wire net830;
 wire _06967_;
 wire _06968_;
 wire net829;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire net828;
 wire net827;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire net826;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire net825;
 wire net824;
 wire net823;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire net822;
 wire _07020_;
 wire _07021_;
 wire net821;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire net820;
 wire net819;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire net818;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire net817;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire net816;
 wire _07073_;
 wire _07074_;
 wire net815;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire net814;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire net813;
 wire net812;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire net811;
 wire _07096_;
 wire _07097_;
 wire net810;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire net809;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire net808;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire net807;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire net806;
 wire _07122_;
 wire net805;
 wire net804;
 wire net803;
 wire net802;
 wire net801;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire net800;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire net799;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire net798;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire net797;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire net796;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire net795;
 wire _07157_;
 wire net794;
 wire _07159_;
 wire net793;
 wire net792;
 wire _07162_;
 wire net791;
 wire net790;
 wire _07165_;
 wire _07166_;
 wire net789;
 wire _07168_;
 wire net788;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire net787;
 wire _07182_;
 wire net786;
 wire _07184_;
 wire net785;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire net784;
 wire _07193_;
 wire _07194_;
 wire net783;
 wire _07196_;
 wire net782;
 wire net781;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire net780;
 wire net779;
 wire _07205_;
 wire _07206_;
 wire net778;
 wire _07208_;
 wire _07209_;
 wire net777;
 wire net776;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire net775;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire net774;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire net773;
 wire net772;
 wire net771;
 wire net770;
 wire net769;
 wire net768;
 wire _07293_;
 wire _07294_;
 wire net767;
 wire _07296_;
 wire _07297_;
 wire net766;
 wire _07299_;
 wire net765;
 wire _07301_;
 wire _07302_;
 wire net764;
 wire net763;
 wire _07305_;
 wire net762;
 wire _07307_;
 wire net761;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire net760;
 wire net759;
 wire _07351_;
 wire net758;
 wire net757;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire net756;
 wire net755;
 wire _07359_;
 wire net754;
 wire net753;
 wire net752;
 wire _07363_;
 wire _07364_;
 wire net751;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire net750;
 wire net749;
 wire _07388_;
 wire net748;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire net747;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire net746;
 wire _07437_;
 wire _07438_;
 wire net745;
 wire net744;
 wire net743;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire net742;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire net741;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire net740;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire net739;
 wire _07507_;
 wire _07508_;
 wire net738;
 wire _07510_;
 wire _07511_;
 wire net737;
 wire _07513_;
 wire net736;
 wire _07515_;
 wire _07516_;
 wire net735;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire net734;
 wire _07526_;
 wire _07527_;
 wire net733;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire net732;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire net731;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire net730;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire net729;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire net728;
 wire net727;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire net726;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire net725;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire net724;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire net723;
 wire net722;
 wire net721;
 wire _07715_;
 wire _07716_;
 wire net720;
 wire _07718_;
 wire _07719_;
 wire net719;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire net718;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire net717;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire net716;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire net715;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire net714;
 wire net713;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire net712;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire net711;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire net710;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire net709;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire net708;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire net707;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire net706;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire net705;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire net704;
 wire net703;
 wire net702;
 wire net701;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire net700;
 wire _08600_;
 wire net699;
 wire net698;
 wire _08603_;
 wire _08604_;
 wire net697;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire net696;
 wire net695;
 wire net694;
 wire _08614_;
 wire net693;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire net692;
 wire net691;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire net690;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire net689;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire net688;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire net687;
 wire _08694_;
 wire _08695_;
 wire net686;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire net685;
 wire net684;
 wire net683;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire net682;
 wire net681;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire net680;
 wire net679;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire net678;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire net677;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire net676;
 wire _08750_;
 wire _08751_;
 wire net675;
 wire net674;
 wire net673;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire net672;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire net671;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire net670;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire net669;
 wire _08788_;
 wire net668;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire net667;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire net666;
 wire net665;
 wire net664;
 wire _09071_;
 wire net663;
 wire net662;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire net661;
 wire net660;
 wire net659;
 wire net658;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire net657;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire net656;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire net655;
 wire net654;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire net653;
 wire _09157_;
 wire _09158_;
 wire net652;
 wire _09160_;
 wire net651;
 wire _09162_;
 wire net650;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire net649;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire net648;
 wire net647;
 wire net646;
 wire _09199_;
 wire _09200_;
 wire net645;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire net644;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire net643;
 wire _09214_;
 wire _09215_;
 wire net642;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire net641;
 wire net640;
 wire net639;
 wire net638;
 wire net637;
 wire _09263_;
 wire net636;
 wire net635;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire net634;
 wire _09270_;
 wire net633;
 wire net632;
 wire net631;
 wire net630;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire net629;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire net628;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire net627;
 wire _09306_;
 wire _09307_;
 wire net626;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire net625;
 wire net624;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire net623;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire net622;
 wire net621;
 wire net620;
 wire net619;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire net618;
 wire net617;
 wire _09370_;
 wire net616;
 wire _09372_;
 wire net615;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire net614;
 wire net613;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire net612;
 wire _09387_;
 wire _09388_;
 wire net611;
 wire _09390_;
 wire _09391_;
 wire net610;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire net609;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire net608;
 wire _09405_;
 wire _09406_;
 wire net607;
 wire _09408_;
 wire net606;
 wire net605;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire net604;
 wire net603;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire net602;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire net601;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire net600;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire net599;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire net598;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire net597;
 wire _09505_;
 wire _09506_;
 wire net596;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire net595;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire net594;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire net593;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire net592;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire net591;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire net590;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire net589;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire net588;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire net587;
 wire _09615_;
 wire net586;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire net585;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire net584;
 wire net583;
 wire net582;
 wire _09669_;
 wire net581;
 wire _09671_;
 wire net580;
 wire _09673_;
 wire net579;
 wire _09675_;
 wire net578;
 wire _09677_;
 wire net577;
 wire _09679_;
 wire net576;
 wire _09681_;
 wire net575;
 wire _09683_;
 wire net574;
 wire net573;
 wire _09686_;
 wire net572;
 wire _09688_;
 wire net571;
 wire net570;
 wire _09691_;
 wire net569;
 wire _09693_;
 wire net568;
 wire _09695_;
 wire net567;
 wire _09697_;
 wire net566;
 wire _09699_;
 wire net565;
 wire _09701_;
 wire net564;
 wire _09703_;
 wire net563;
 wire _09705_;
 wire net562;
 wire net561;
 wire _09708_;
 wire net560;
 wire _09710_;
 wire net559;
 wire net558;
 wire _09713_;
 wire net557;
 wire _09715_;
 wire net556;
 wire _09717_;
 wire net555;
 wire _09719_;
 wire net554;
 wire _09721_;
 wire net553;
 wire _09723_;
 wire net552;
 wire _09725_;
 wire net551;
 wire _09727_;
 wire net550;
 wire _09729_;
 wire net549;
 wire _09731_;
 wire net548;
 wire _09733_;
 wire net547;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire net546;
 wire net545;
 wire net544;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire net543;
 wire _09751_;
 wire _09752_;
 wire net542;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire net541;
 wire _09763_;
 wire _09764_;
 wire net540;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire net539;
 wire net538;
 wire net537;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire net536;
 wire _09793_;
 wire _09794_;
 wire net535;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire net534;
 wire _09805_;
 wire _09806_;
 wire net533;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire net532;
 wire net531;
 wire net530;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire net529;
 wire _09833_;
 wire _09834_;
 wire net528;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire net527;
 wire _09845_;
 wire _09846_;
 wire net526;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire net525;
 wire net524;
 wire net523;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire net522;
 wire _09873_;
 wire _09874_;
 wire net521;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire net520;
 wire _09885_;
 wire _09886_;
 wire net519;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire net518;
 wire net517;
 wire net516;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire net515;
 wire _09913_;
 wire _09914_;
 wire net514;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire net513;
 wire _09925_;
 wire _09926_;
 wire net512;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire net511;
 wire net510;
 wire net509;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire net508;
 wire _09954_;
 wire _09955_;
 wire net507;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire net506;
 wire _09966_;
 wire _09967_;
 wire net505;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire net504;
 wire net503;
 wire net502;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire net501;
 wire _09994_;
 wire _09995_;
 wire net500;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire net499;
 wire _10006_;
 wire _10007_;
 wire net498;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire net497;
 wire net496;
 wire net495;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire net494;
 wire _10034_;
 wire _10035_;
 wire net493;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire net492;
 wire _10046_;
 wire _10047_;
 wire net491;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire net490;
 wire net489;
 wire net488;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire net487;
 wire _10074_;
 wire _10075_;
 wire net486;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire net485;
 wire _10086_;
 wire _10087_;
 wire net484;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire net483;
 wire _10102_;
 wire _10103_;
 wire net482;
 wire net481;
 wire net480;
 wire _10107_;
 wire net479;
 wire _10109_;
 wire net478;
 wire _10111_;
 wire net477;
 wire _10113_;
 wire net476;
 wire _10115_;
 wire net475;
 wire _10117_;
 wire net474;
 wire _10119_;
 wire net473;
 wire _10121_;
 wire net472;
 wire net471;
 wire _10124_;
 wire net470;
 wire _10126_;
 wire net469;
 wire net468;
 wire _10129_;
 wire net467;
 wire _10131_;
 wire net466;
 wire _10133_;
 wire net465;
 wire _10135_;
 wire net464;
 wire _10137_;
 wire net463;
 wire _10139_;
 wire net462;
 wire _10141_;
 wire net461;
 wire _10143_;
 wire net460;
 wire net459;
 wire _10146_;
 wire net458;
 wire _10148_;
 wire net457;
 wire net455;
 wire _10151_;
 wire net454;
 wire _10153_;
 wire net453;
 wire _10155_;
 wire net452;
 wire _10157_;
 wire net451;
 wire _10159_;
 wire net450;
 wire _10161_;
 wire net449;
 wire _10163_;
 wire net448;
 wire _10165_;
 wire net447;
 wire _10167_;
 wire net446;
 wire _10169_;
 wire net445;
 wire _10171_;
 wire net444;
 wire _10173_;
 wire _10174_;
 wire net443;
 wire net442;
 wire net441;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire net440;
 wire _10187_;
 wire _10188_;
 wire net439;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire net438;
 wire _10199_;
 wire _10200_;
 wire net437;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire net436;
 wire net435;
 wire net434;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire net433;
 wire _10227_;
 wire _10228_;
 wire net432;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire net431;
 wire _10239_;
 wire _10240_;
 wire net430;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire net429;
 wire net428;
 wire net427;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire net426;
 wire _10267_;
 wire _10268_;
 wire net425;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire net424;
 wire _10279_;
 wire _10280_;
 wire net423;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire net422;
 wire net421;
 wire net420;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire net419;
 wire _10307_;
 wire _10308_;
 wire net418;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire net417;
 wire _10319_;
 wire _10320_;
 wire net416;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire net415;
 wire _10336_;
 wire net414;
 wire net413;
 wire net412;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire net411;
 wire _10349_;
 wire _10350_;
 wire net410;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire net409;
 wire _10361_;
 wire _10362_;
 wire net408;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire net407;
 wire net406;
 wire net405;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire net404;
 wire _10389_;
 wire _10390_;
 wire net403;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire net402;
 wire _10401_;
 wire _10402_;
 wire net401;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire net400;
 wire net399;
 wire net398;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire net397;
 wire _10429_;
 wire _10430_;
 wire net396;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire net395;
 wire _10441_;
 wire _10442_;
 wire net394;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire net393;
 wire net392;
 wire net391;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire net390;
 wire _10469_;
 wire _10470_;
 wire net389;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire net388;
 wire _10481_;
 wire _10482_;
 wire net387;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire net386;
 wire net385;
 wire net384;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire net383;
 wire _10509_;
 wire _10510_;
 wire net382;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire net381;
 wire _10521_;
 wire _10522_;
 wire net380;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire net379;
 wire _10537_;
 wire net378;
 wire net377;
 wire net376;
 wire _10541_;
 wire net375;
 wire _10543_;
 wire net374;
 wire _10545_;
 wire net373;
 wire _10547_;
 wire net372;
 wire _10549_;
 wire net371;
 wire _10551_;
 wire net370;
 wire _10553_;
 wire net369;
 wire _10555_;
 wire net368;
 wire net367;
 wire _10558_;
 wire net366;
 wire _10560_;
 wire net365;
 wire net364;
 wire _10563_;
 wire net363;
 wire _10565_;
 wire net362;
 wire _10567_;
 wire net361;
 wire _10569_;
 wire net360;
 wire _10571_;
 wire net359;
 wire _10573_;
 wire net358;
 wire _10575_;
 wire net357;
 wire _10577_;
 wire net356;
 wire net355;
 wire _10580_;
 wire net354;
 wire _10582_;
 wire net353;
 wire net352;
 wire _10585_;
 wire net351;
 wire _10587_;
 wire net350;
 wire _10589_;
 wire net349;
 wire _10591_;
 wire net348;
 wire _10593_;
 wire net347;
 wire _10595_;
 wire net346;
 wire _10597_;
 wire net345;
 wire _10599_;
 wire net344;
 wire _10601_;
 wire net343;
 wire _10603_;
 wire net342;
 wire _10605_;
 wire net341;
 wire _10607_;
 wire _10608_;
 wire net340;
 wire net339;
 wire net338;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire net337;
 wire _10621_;
 wire _10622_;
 wire net336;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire net335;
 wire _10633_;
 wire _10634_;
 wire net334;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire net333;
 wire net332;
 wire net331;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire net330;
 wire _10661_;
 wire _10662_;
 wire net329;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire net328;
 wire _10673_;
 wire _10674_;
 wire net327;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire net326;
 wire net325;
 wire net324;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire net323;
 wire _10701_;
 wire _10702_;
 wire net322;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire net321;
 wire _10713_;
 wire _10714_;
 wire net320;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire net319;
 wire net318;
 wire net317;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire net316;
 wire _10741_;
 wire _10742_;
 wire net315;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire net314;
 wire _10753_;
 wire _10754_;
 wire net313;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire net312;
 wire net311;
 wire net310;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire net309;
 wire _10781_;
 wire _10782_;
 wire net308;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire net307;
 wire _10793_;
 wire _10794_;
 wire net306;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire net305;
 wire net304;
 wire net303;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire net302;
 wire _10821_;
 wire _10822_;
 wire net301;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire net300;
 wire _10833_;
 wire _10834_;
 wire net299;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire net298;
 wire net297;
 wire net296;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire net295;
 wire _10861_;
 wire _10862_;
 wire net294;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire net293;
 wire _10873_;
 wire _10874_;
 wire net292;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire net291;
 wire net290;
 wire net289;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire net288;
 wire _10901_;
 wire _10902_;
 wire net287;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire net286;
 wire _10913_;
 wire _10914_;
 wire net285;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire net284;
 wire net283;
 wire net282;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire net281;
 wire _10941_;
 wire _10942_;
 wire net280;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire net279;
 wire _10953_;
 wire _10954_;
 wire net278;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire net277;
 wire _10978_;
 wire net276;
 wire net275;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire net274;
 wire _10988_;
 wire _10989_;
 wire net273;
 wire _10991_;
 wire _10992_;
 wire net272;
 wire net271;
 wire _10995_;
 wire net270;
 wire _10997_;
 wire net269;
 wire net268;
 wire _11000_;
 wire net267;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire net266;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire net265;
 wire net264;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire net263;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire net262;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire net261;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire net260;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire net259;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire net258;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire net257;
 wire _11104_;
 wire _11105_;
 wire net256;
 wire _11107_;
 wire _11108_;
 wire net255;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire net254;
 wire net253;
 wire _11115_;
 wire _11116_;
 wire net252;
 wire net251;
 wire _11119_;
 wire net250;
 wire net249;
 wire net248;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire net247;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire net246;
 wire net245;
 wire _11133_;
 wire _11134_;
 wire net244;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire net243;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire net242;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire net241;
 wire _11228_;
 wire _11229_;
 wire net240;
 wire _11231_;
 wire net239;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire net238;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire net237;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire net236;
 wire net235;
 wire _11255_;
 wire _11256_;
 wire net234;
 wire net233;
 wire _11259_;
 wire net232;
 wire _11261_;
 wire net231;
 wire _11263_;
 wire _11264_;
 wire net230;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire net229;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire net228;
 wire _11293_;
 wire net227;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire net226;
 wire net225;
 wire net224;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire net223;
 wire net222;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire net221;
 wire net220;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire net219;
 wire _11362_;
 wire _11363_;
 wire net218;
 wire _11365_;
 wire net217;
 wire _11367_;
 wire _11368_;
 wire net216;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire net215;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire net214;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire net213;
 wire net212;
 wire net211;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire net210;
 wire _11457_;
 wire _11458_;
 wire net209;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire net208;
 wire _11469_;
 wire _11470_;
 wire net207;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire net206;
 wire net205;
 wire net204;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire net203;
 wire net202;
 wire net201;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire net200;
 wire _11512_;
 wire _11513_;
 wire net199;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire net198;
 wire _11524_;
 wire _11525_;
 wire net197;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire net196;
 wire net195;
 wire net194;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire net193;
 wire net192;
 wire net191;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire net190;
 wire _11603_;
 wire _11604_;
 wire net189;
 wire net188;
 wire _11607_;
 wire _11608_;
 wire net187;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire net186;
 wire _11618_;
 wire net185;
 wire _11620_;
 wire _11621_;
 wire net184;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire net183;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire net182;
 wire _11708_;
 wire net181;
 wire net180;
 wire net179;
 wire net178;
 wire net177;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire net176;
 wire net175;
 wire _11723_;
 wire _11724_;
 wire net174;
 wire _11726_;
 wire net173;
 wire _11728_;
 wire net172;
 wire net171;
 wire net170;
 wire net169;
 wire _11733_;
 wire net168;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire net167;
 wire _11741_;
 wire net166;
 wire net165;
 wire net164;
 wire _11745_;
 wire _11746_;
 wire net163;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire net162;
 wire net161;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire net160;
 wire net159;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire net158;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire net157;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire net156;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire net155;
 wire _11833_;
 wire net154;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire net153;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire net152;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire net151;
 wire net150;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire net149;
 wire _11989_;
 wire net148;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire net147;
 wire _12001_;
 wire net146;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire net145;
 wire _12016_;
 wire net144;
 wire net143;
 wire net142;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire net141;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire net140;
 wire net139;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire net138;
 wire net137;
 wire net136;
 wire _12059_;
 wire _12060_;
 wire net135;
 wire _12062_;
 wire net134;
 wire net133;
 wire _12065_;
 wire _12066_;
 wire net132;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire net131;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire net130;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire net129;
 wire _12169_;
 wire _12170_;
 wire net128;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire net127;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire net126;
 wire _12185_;
 wire _12186_;
 wire net125;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire net124;
 wire net123;
 wire _12216_;
 wire net122;
 wire net121;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire net120;
 wire net119;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire net118;
 wire _12249_;
 wire net117;
 wire net116;
 wire net115;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire net114;
 wire net113;
 wire _12262_;
 wire _12263_;
 wire net112;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire net111;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire net110;
 wire _12301_;
 wire _12302_;
 wire net109;
 wire net108;
 wire net107;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire net106;
 wire net105;
 wire net104;
 wire net103;
 wire net102;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire net101;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire net100;
 wire net99;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire net98;
 wire net97;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire net96;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire net95;
 wire net94;
 wire net93;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire net92;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire net91;
 wire net90;
 wire net89;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire net88;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire net87;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire net86;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire net85;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire net84;
 wire net83;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire net82;
 wire net81;
 wire net80;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire net79;
 wire net78;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire net77;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire net76;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire net75;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire net74;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire net73;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire net72;
 wire _12564_;
 wire net71;
 wire net70;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire net69;
 wire net68;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire net67;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire net66;
 wire net65;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire net64;
 wire net63;
 wire net62;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire net61;
 wire net60;
 wire net59;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire net58;
 wire net57;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire net56;
 wire net55;
 wire _12629_;
 wire net54;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire net53;
 wire _12649_;
 wire net52;
 wire _12651_;
 wire net51;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire net50;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire net49;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire net48;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire net47;
 wire _12709_;
 wire net46;
 wire _12711_;
 wire _12712_;
 wire net45;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire net44;
 wire net43;
 wire _12720_;
 wire net42;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire net41;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire net40;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire net39;
 wire _12755_;
 wire _12756_;
 wire net38;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire net37;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire net36;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire net35;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire net34;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire net33;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire net32;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire net31;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire net30;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire net1632;
 wire net1631;
 wire net1630;
 wire _13122_;
 wire net1629;
 wire _13124_;
 wire net1628;
 wire net1627;
 wire _13127_;
 wire net1626;
 wire net1625;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire net1624;
 wire net1623;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire net1622;
 wire net1621;
 wire net1620;
 wire net1619;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire net1618;
 wire net1617;
 wire _13148_;
 wire net1616;
 wire _13150_;
 wire _13151_;
 wire net1615;
 wire net1614;
 wire _13154_;
 wire net1613;
 wire _13156_;
 wire net1612;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire net1611;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire net1610;
 wire net1609;
 wire net1608;
 wire net1607;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire net1606;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire net1605;
 wire _13179_;
 wire net1604;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire net1603;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire net1602;
 wire _13198_;
 wire net1601;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire net1600;
 wire net1599;
 wire _13208_;
 wire net1598;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire net1597;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire net1596;
 wire net1595;
 wire net1594;
 wire _13227_;
 wire _13228_;
 wire net1593;
 wire _13230_;
 wire net1592;
 wire net1591;
 wire net1590;
 wire _13234_;
 wire _13235_;
 wire net1589;
 wire net1588;
 wire _13238_;
 wire _13239_;
 wire net1587;
 wire net1586;
 wire net1585;
 wire net1584;
 wire net1583;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire net1582;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire net1581;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire net1580;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire net1579;
 wire _13293_;
 wire net1578;
 wire net1577;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire net1575;
 wire net1573;
 wire net1572;
 wire _13306_;
 wire net1571;
 wire net1570;
 wire net1569;
 wire net1568;
 wire _13311_;
 wire net1567;
 wire _13313_;
 wire net1566;
 wire net1565;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire net1564;
 wire net1563;
 wire net1562;
 wire net1561;
 wire _13323_;
 wire net1560;
 wire _13325_;
 wire net1559;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire net1558;
 wire _13332_;
 wire _13333_;
 wire net1557;
 wire _13335_;
 wire _13336_;
 wire net1556;
 wire _13338_;
 wire net1555;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire net1554;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire net1553;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire net1552;
 wire _13389_;
 wire net1551;
 wire net1550;
 wire _13392_;
 wire net1549;
 wire net1548;
 wire net1547;
 wire net1546;
 wire _13397_;
 wire net1545;
 wire net1544;
 wire net1543;
 wire net1542;
 wire net1541;
 wire _13403_;
 wire net1540;
 wire net1539;
 wire net1538;
 wire net1537;
 wire net1536;
 wire net1535;
 wire net1534;
 wire net1533;
 wire net1532;
 wire _13413_;
 wire net1531;
 wire net1530;
 wire net1529;
 wire net1528;
 wire _13418_;
 wire _13419_;
 wire net1527;
 wire net1526;
 wire net1525;
 wire _13423_;
 wire _13424_;
 wire net1524;
 wire net1523;
 wire _13427_;
 wire _13428_;
 wire net1522;
 wire net1521;
 wire net1520;
 wire net1519;
 wire _13433_;
 wire net1518;
 wire net1517;
 wire net1516;
 wire net1515;
 wire net1514;
 wire net1513;
 wire _13440_;
 wire _13441_;
 wire net1512;
 wire net1511;
 wire net1510;
 wire net1509;
 wire net1508;
 wire net1507;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire net1506;
 wire net1505;
 wire net1504;
 wire net1503;
 wire _13456_;
 wire _13457_;
 wire net1502;
 wire net1501;
 wire net1500;
 wire net1499;
 wire net1498;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire net1497;
 wire net1496;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire net1495;
 wire net1494;
 wire net1493;
 wire net1492;
 wire _13477_;
 wire _13478_;
 wire net1491;
 wire net1490;
 wire net1489;
 wire net1488;
 wire net1487;
 wire _13484_;
 wire _13485_;
 wire net1486;
 wire net1485;
 wire net1484;
 wire _13489_;
 wire net1483;
 wire _13491_;
 wire _13492_;
 wire net1482;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire net1481;
 wire net1480;
 wire net1479;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire net1478;
 wire net1477;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire net1476;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire net1475;
 wire net1474;
 wire net1473;
 wire _13527_;
 wire _13528_;
 wire net1472;
 wire _13530_;
 wire net1471;
 wire net1470;
 wire _13533_;
 wire net1469;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire net1468;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire net1467;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire net1466;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire net1465;
 wire _13563_;
 wire net1464;
 wire net1463;
 wire net1462;
 wire _13567_;
 wire net1461;
 wire _13569_;
 wire _13570_;
 wire net1460;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire net1458;
 wire _13576_;
 wire net1457;
 wire net1456;
 wire net1455;
 wire net1454;
 wire net1453;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire net1452;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire net1451;
 wire _13606_;
 wire _13607_;
 wire net1450;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire net1449;
 wire net1448;
 wire net1447;
 wire _13644_;
 wire _13645_;
 wire net1446;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire net1445;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire net1444;
 wire _13658_;
 wire net1443;
 wire net1442;
 wire net1441;
 wire net1439;
 wire net1438;
 wire net1437;
 wire net1435;
 wire net1434;
 wire net1433;
 wire net1432;
 wire net1431;
 wire net1430;
 wire net1429;
 wire net1428;
 wire net1427;
 wire net1426;
 wire _13675_;
 wire _13676_;
 wire net1425;
 wire _13678_;
 wire net1424;
 wire net1423;
 wire net1422;
 wire _13682_;
 wire net1421;
 wire _13684_;
 wire net1420;
 wire net1419;
 wire net1418;
 wire _13688_;
 wire net1417;
 wire _13690_;
 wire net1416;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire net1415;
 wire net1414;
 wire net1413;
 wire net1412;
 wire _13699_;
 wire net1411;
 wire _13701_;
 wire _13702_;
 wire net1410;
 wire _13704_;
 wire _13705_;
 wire net1409;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire net1408;
 wire net1407;
 wire net1406;
 wire _13720_;
 wire net1405;
 wire _13722_;
 wire net1404;
 wire net1403;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire net1402;
 wire net1401;
 wire _13730_;
 wire _13731_;
 wire net1400;
 wire net1399;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire net1398;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire net1397;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire net1396;
 wire _13748_;
 wire net1395;
 wire net1394;
 wire _13751_;
 wire net1393;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire net1392;
 wire net1391;
 wire net1390;
 wire _13762_;
 wire _13763_;
 wire net1389;
 wire _13765_;
 wire _13766_;
 wire net1388;
 wire net1387;
 wire net1386;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire net1385;
 wire net1384;
 wire _13776_;
 wire _13777_;
 wire net1382;
 wire net1381;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire net1379;
 wire net1378;
 wire net1377;
 wire net1376;
 wire net1375;
 wire net1374;
 wire _13789_;
 wire net1373;
 wire _13791_;
 wire _13792_;
 wire net1372;
 wire _13794_;
 wire net1371;
 wire _13796_;
 wire net1370;
 wire net1369;
 wire _13799_;
 wire _13800_;
 wire net1368;
 wire _13802_;
 wire _13803_;
 wire net1367;
 wire _13805_;
 wire net1366;
 wire net1365;
 wire _13808_;
 wire _13809_;
 wire net1364;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire net1363;
 wire net1362;
 wire net1361;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire net1360;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire net1359;
 wire net1358;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire net1357;
 wire _13835_;
 wire net1356;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire net1355;
 wire net1354;
 wire net1353;
 wire net1352;
 wire _13847_;
 wire _13848_;
 wire net1351;
 wire net1350;
 wire _13851_;
 wire _13852_;
 wire net1349;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire net1348;
 wire net1347;
 wire _13860_;
 wire _13861_;
 wire net1346;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire net1345;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire net1344;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire net1343;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire net1342;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire net1341;
 wire _13922_;
 wire _13923_;
 wire net1340;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire net1339;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire net1338;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire net1337;
 wire _13945_;
 wire net1336;
 wire net1335;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire net1334;
 wire net1332;
 wire net1331;
 wire net1330;
 wire net1329;
 wire _13961_;
 wire _13962_;
 wire net1328;
 wire _13964_;
 wire _13965_;
 wire net1327;
 wire _13967_;
 wire _13968_;
 wire net1326;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire net1325;
 wire _13985_;
 wire _13986_;
 wire net1324;
 wire net1323;
 wire _13989_;
 wire _13990_;
 wire net1322;
 wire net1321;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire net1320;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire net1319;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire net1318;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire net1315;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire net1314;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire net1309;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire net1308;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire net1306;
 wire net1305;
 wire _14259_;
 wire net1304;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire net1303;
 wire _14265_;
 wire _14266_;
 wire net1302;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire net1301;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire net1300;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire net1298;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire net1297;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire net1295;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire net1294;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire net1293;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire net1292;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire net1291;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire net1289;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire net1287;
 wire net1286;
 wire net1285;
 wire net1284;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire net1283;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire net1282;
 wire net1281;
 wire _14528_;
 wire net1280;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire net1279;
 wire net1278;
 wire net1277;
 wire _14537_;
 wire _14538_;
 wire net1276;
 wire net1275;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire net1274;
 wire _14545_;
 wire net1273;
 wire _14547_;
 wire net1272;
 wire _14549_;
 wire net1271;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire net1270;
 wire net1269;
 wire net1268;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire net1267;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire net1266;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire net1264;
 wire net1263;
 wire _14580_;
 wire _14581_;
 wire net1262;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire net1261;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire net1260;
 wire _14628_;
 wire net1259;
 wire net1258;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire net1257;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire net1256;
 wire net1255;
 wire net1254;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire net1253;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire net1251;
 wire _14691_;
 wire _14692_;
 wire net1250;
 wire _14694_;
 wire _14695_;
 wire net1249;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire net1248;
 wire _14702_;
 wire net1247;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire net1246;
 wire net1245;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire net1244;
 wire _14717_;
 wire net1243;
 wire _14719_;
 wire _14720_;
 wire net1242;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire net1241;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire net1240;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire net1238;
 wire _14766_;
 wire net1237;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire net1236;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire net1235;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire net1234;
 wire _14794_;
 wire net1233;
 wire _14796_;
 wire net1232;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire net1231;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire net1229;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire net1228;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire net1227;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire net1226;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire net1225;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire net1224;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire net1222;
 wire _14950_;
 wire _14951_;
 wire net1221;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire net1220;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire net1219;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire net1218;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire net1217;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire net1216;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire net1213;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire net1212;
 wire net1211;
 wire net1210;
 wire net1209;
 wire net1208;
 wire net1207;
 wire net1206;
 wire net1205;
 wire net1204;
 wire net1203;
 wire net1202;
 wire net1201;
 wire _15181_;
 wire _15182_;
 wire net1200;
 wire net1199;
 wire net1198;
 wire net1197;
 wire _15187_;
 wire net1196;
 wire net1195;
 wire net1194;
 wire net1193;
 wire net1192;
 wire net1191;
 wire net1190;
 wire _15195_;
 wire net1189;
 wire net1188;
 wire _15198_;
 wire _15199_;
 wire net1187;
 wire _15201_;
 wire _15202_;
 wire net1186;
 wire net1185;
 wire net1184;
 wire _15206_;
 wire net1183;
 wire net1182;
 wire net1181;
 wire net1180;
 wire net1179;
 wire net1178;
 wire _15213_;
 wire _15214_;
 wire net1177;
 wire net1176;
 wire net1175;
 wire _15218_;
 wire net1174;
 wire net1173;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire net1172;
 wire net1171;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire net1170;
 wire net1169;
 wire _15232_;
 wire _15233_;
 wire net1168;
 wire net1167;
 wire _15236_;
 wire _15237_;
 wire net1166;
 wire net1165;
 wire net1164;
 wire _15241_;
 wire net1163;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire net1162;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire net1161;
 wire net1160;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire net1159;
 wire net1158;
 wire net1157;
 wire net1156;
 wire net1155;
 wire _15276_;
 wire net1154;
 wire _15278_;
 wire _15279_;
 wire net1153;
 wire _15281_;
 wire net1152;
 wire net1151;
 wire _15284_;
 wire net1150;
 wire net1149;
 wire _15287_;
 wire _15288_;
 wire net1148;
 wire net1147;
 wire net1146;
 wire _15292_;
 wire _15293_;
 wire net1145;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire net1144;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire net1143;
 wire _15317_;
 wire net1142;
 wire _15319_;
 wire _15320_;
 wire net1141;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire net1140;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire net1139;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire net1138;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire net1137;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire net1136;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire net1134;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire net1133;
 wire net1132;
 wire net1131;
 wire _15421_;
 wire net1130;
 wire _15423_;
 wire net1129;
 wire _15425_;
 wire net1128;
 wire net1127;
 wire _15428_;
 wire _15429_;
 wire net1126;
 wire net1125;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire net1124;
 wire _15437_;
 wire _15438_;
 wire net1123;
 wire _15440_;
 wire _15441_;
 wire net1122;
 wire net1121;
 wire _15444_;
 wire _15445_;
 wire net1120;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire net1119;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire net1118;
 wire _15461_;
 wire _15462_;
 wire net1117;
 wire net1116;
 wire _15465_;
 wire _15466_;
 wire net1115;
 wire _15468_;
 wire _15469_;
 wire net1114;
 wire _15471_;
 wire net1113;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire net1112;
 wire net1111;
 wire _15485_;
 wire net1110;
 wire net1109;
 wire _15488_;
 wire _15489_;
 wire net1108;
 wire net1107;
 wire net1106;
 wire _15493_;
 wire _15494_;
 wire net1105;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire net1104;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire net1103;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire net1101;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire net1099;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire net1097;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire net1096;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire net1095;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire net1093;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire net1091;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire net1090;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire net1089;
 wire _15915_;
 wire _15916_;
 wire net1088;
 wire _15918_;
 wire net1087;
 wire _15920_;
 wire _15921_;
 wire net1086;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire net1085;
 wire _15929_;
 wire net1084;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire net1083;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire net1082;
 wire _15954_;
 wire _15955_;
 wire net1081;
 wire net1080;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire net1079;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire net1078;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire net1076;
 wire _16207_;
 wire net1075;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire net1074;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire net1072;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire net1071;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire net1070;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16331_;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16392_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire net1068;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire net1067;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire _16460_;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire _16468_;
 wire _16469_;
 wire _16470_;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire net1380;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire _16525_;
 wire _16526_;
 wire _16527_;
 wire _16528_;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire _16536_;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire _16552_;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire _16560_;
 wire _16561_;
 wire _16562_;
 wire _16563_;
 wire _16564_;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire _16569_;
 wire _16570_;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire _16624_;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire _16639_;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire _16698_;
 wire _16699_;
 wire _16700_;
 wire _16701_;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire _16707_;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire _16716_;
 wire _16717_;
 wire _16718_;
 wire _16719_;
 wire _16720_;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire _16745_;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire _16754_;
 wire _16755_;
 wire _16756_;
 wire _16757_;
 wire _16758_;
 wire _16759_;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire _16766_;
 wire _16767_;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire _16771_;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire _16776_;
 wire _16777_;
 wire _16778_;
 wire _16779_;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire _16791_;
 wire _16792_;
 wire _16793_;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire _16797_;
 wire _16798_;
 wire _16799_;
 wire _16800_;
 wire _16801_;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire _16805_;
 wire _16806_;
 wire _16807_;
 wire _16808_;
 wire _16809_;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire _16816_;
 wire _16817_;
 wire _16818_;
 wire _16819_;
 wire _16820_;
 wire _16821_;
 wire _16822_;
 wire _16823_;
 wire _16824_;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire _16828_;
 wire _16829_;
 wire _16830_;
 wire _16831_;
 wire _16832_;
 wire _16833_;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire _16837_;
 wire _16838_;
 wire _16839_;
 wire _16840_;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire _16848_;
 wire _16849_;
 wire _16850_;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire _16854_;
 wire _16855_;
 wire _16856_;
 wire _16857_;
 wire _16858_;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire _16862_;
 wire _16863_;
 wire _16864_;
 wire _16865_;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire _16869_;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire _16875_;
 wire _16876_;
 wire _16877_;
 wire _16878_;
 wire _16879_;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire _16884_;
 wire _16885_;
 wire _16886_;
 wire _16887_;
 wire _16888_;
 wire _16889_;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire _16895_;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire _16901_;
 wire _16902_;
 wire net955;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire _16907_;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire _16911_;
 wire _16912_;
 wire _16913_;
 wire _16914_;
 wire _16915_;
 wire _16916_;
 wire _16917_;
 wire _16918_;
 wire _16919_;
 wire _16920_;
 wire _16921_;
 wire _16922_;
 wire _16923_;
 wire _16924_;
 wire _16925_;
 wire _16926_;
 wire _16927_;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire _16936_;
 wire _16937_;
 wire _16938_;
 wire _16939_;
 wire _16940_;
 wire _16941_;
 wire _16942_;
 wire _16943_;
 wire _16944_;
 wire _16945_;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire _16949_;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire _16953_;
 wire _16954_;
 wire _16955_;
 wire _16956_;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire _16962_;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire _16975_;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire _16981_;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire _16985_;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire _16992_;
 wire _16993_;
 wire _16994_;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire _17007_;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire _17032_;
 wire _17033_;
 wire _17034_;
 wire _17035_;
 wire _17036_;
 wire _17037_;
 wire _17038_;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire _17055_;
 wire _17056_;
 wire _17057_;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire _17061_;
 wire _17062_;
 wire _17063_;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire _17067_;
 wire _17068_;
 wire _17069_;
 wire _17070_;
 wire _17071_;
 wire _17072_;
 wire _17073_;
 wire _17074_;
 wire _17075_;
 wire _17076_;
 wire _17077_;
 wire _17078_;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire _17082_;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire _17091_;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire _17095_;
 wire _17096_;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire _17100_;
 wire _17101_;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire _17106_;
 wire _17107_;
 wire _17108_;
 wire _17109_;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire _17121_;
 wire _17122_;
 wire _17123_;
 wire _17124_;
 wire _17125_;
 wire _17126_;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire _17130_;
 wire _17131_;
 wire _17132_;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire _17137_;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire _17141_;
 wire _17142_;
 wire _17143_;
 wire _17144_;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire _17150_;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire _17156_;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire _17160_;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire _17169_;
 wire _17170_;
 wire _17171_;
 wire _17172_;
 wire _17173_;
 wire _17174_;
 wire _17175_;
 wire _17176_;
 wire _17177_;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire _17183_;
 wire _17184_;
 wire _17185_;
 wire _17186_;
 wire _17187_;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire _17196_;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire _17206_;
 wire _17207_;
 wire _17208_;
 wire _17209_;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire _17215_;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire _17228_;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire _17238_;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire _17245_;
 wire _17246_;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire _17259_;
 wire _17260_;
 wire _17261_;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire _17267_;
 wire _17268_;
 wire _17269_;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire _17275_;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire _17280_;
 wire _17281_;
 wire _17282_;
 wire _17283_;
 wire _17284_;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire _17290_;
 wire _17291_;
 wire _17292_;
 wire _17293_;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire _17302_;
 wire _17303_;
 wire _17304_;
 wire _17305_;
 wire _17306_;
 wire _17307_;
 wire _17308_;
 wire _17309_;
 wire _17310_;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire _17317_;
 wire _17318_;
 wire _17319_;
 wire _17320_;
 wire _17321_;
 wire _17322_;
 wire _17323_;
 wire _17324_;
 wire _17325_;
 wire _17326_;
 wire _17327_;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire _17334_;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire _17339_;
 wire _17340_;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire _17350_;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire _17354_;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire _17358_;
 wire _17359_;
 wire _17360_;
 wire _17361_;
 wire _17362_;
 wire _17363_;
 wire _17364_;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire _17372_;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire _17377_;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire _17384_;
 wire _17385_;
 wire _17386_;
 wire _17387_;
 wire _17388_;
 wire _17389_;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire _17397_;
 wire _17398_;
 wire _17399_;
 wire _17400_;
 wire _17401_;
 wire _17402_;
 wire _17403_;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire _17408_;
 wire _17409_;
 wire _17410_;
 wire _17411_;
 wire _17412_;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire _17422_;
 wire _17423_;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire _17432_;
 wire _17433_;
 wire _17434_;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire _17438_;
 wire _17439_;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire _17447_;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire _17451_;
 wire _17452_;
 wire _17453_;
 wire _17454_;
 wire _17455_;
 wire _17456_;
 wire _17457_;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire _17464_;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire _17470_;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire _17474_;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire _17482_;
 wire _17483_;
 wire _17484_;
 wire _17485_;
 wire _17486_;
 wire _17487_;
 wire _17488_;
 wire _17489_;
 wire _17490_;
 wire _17491_;
 wire _17492_;
 wire _17493_;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire _17499_;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire _17504_;
 wire _17505_;
 wire _17506_;
 wire _17507_;
 wire _17508_;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire _17522_;
 wire _17523_;
 wire _17524_;
 wire _17525_;
 wire _17526_;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire _17531_;
 wire _17532_;
 wire _17533_;
 wire _17534_;
 wire _17535_;
 wire _17536_;
 wire _17537_;
 wire _17538_;
 wire _17539_;
 wire _17540_;
 wire _17541_;
 wire _17542_;
 wire _17543_;
 wire _17544_;
 wire _17545_;
 wire _17546_;
 wire _17547_;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire _17552_;
 wire _17553_;
 wire _17554_;
 wire _17555_;
 wire _17556_;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire _17562_;
 wire _17563_;
 wire _17564_;
 wire _17565_;
 wire _17566_;
 wire _17567_;
 wire _17568_;
 wire _17569_;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire _17583_;
 wire _17584_;
 wire _17585_;
 wire _17586_;
 wire _17587_;
 wire _17588_;
 wire net1051;
 wire _17590_;
 wire _17591_;
 wire _17592_;
 wire _17593_;
 wire _17594_;
 wire net853;
 wire net1288;
 wire _17597_;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire _17602_;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire _17606_;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire _17611_;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire _17615_;
 wire _17616_;
 wire _17617_;
 wire _17618_;
 wire _17619_;
 wire _17620_;
 wire _17621_;
 wire _17622_;
 wire _17623_;
 wire _17624_;
 wire _17625_;
 wire _17626_;
 wire _17627_;
 wire _17628_;
 wire _17629_;
 wire _17630_;
 wire _17631_;
 wire _17632_;
 wire _17633_;
 wire _17634_;
 wire _17635_;
 wire _17636_;
 wire _17637_;
 wire _17638_;
 wire _17639_;
 wire _17640_;
 wire _17641_;
 wire _17642_;
 wire _17643_;
 wire _17644_;
 wire _17645_;
 wire _17646_;
 wire _17647_;
 wire _17648_;
 wire _17649_;
 wire _17650_;
 wire _17651_;
 wire _17652_;
 wire _17653_;
 wire _17654_;
 wire _17655_;
 wire _17656_;
 wire _17657_;
 wire _17658_;
 wire _17659_;
 wire _17660_;
 wire _17661_;
 wire _17662_;
 wire _17663_;
 wire _17664_;
 wire _17665_;
 wire _17666_;
 wire _17667_;
 wire _17668_;
 wire _17669_;
 wire _17670_;
 wire _17671_;
 wire _17672_;
 wire _17673_;
 wire _17674_;
 wire _17675_;
 wire _17676_;
 wire _17677_;
 wire _17678_;
 wire _17679_;
 wire _17680_;
 wire _17681_;
 wire _17682_;
 wire _17683_;
 wire _17684_;
 wire _17685_;
 wire _17686_;
 wire _17687_;
 wire _17688_;
 wire _17689_;
 wire _17690_;
 wire _17691_;
 wire _17692_;
 wire _17693_;
 wire _17694_;
 wire _17695_;
 wire _17696_;
 wire _17697_;
 wire _17698_;
 wire _17699_;
 wire _17700_;
 wire _17701_;
 wire _17702_;
 wire _17703_;
 wire _17704_;
 wire _17705_;
 wire _17706_;
 wire _17707_;
 wire _17708_;
 wire _17709_;
 wire _17710_;
 wire _17711_;
 wire _17712_;
 wire _17713_;
 wire _17714_;
 wire _17715_;
 wire _17716_;
 wire _17717_;
 wire _17718_;
 wire _17719_;
 wire _17720_;
 wire _17721_;
 wire _17722_;
 wire _17723_;
 wire _17724_;
 wire _17725_;
 wire _17726_;
 wire _17727_;
 wire _17728_;
 wire _17729_;
 wire _17730_;
 wire _17731_;
 wire _17732_;
 wire _17733_;
 wire _17734_;
 wire _17735_;
 wire _17736_;
 wire _17737_;
 wire _17738_;
 wire _17739_;
 wire _17740_;
 wire _17741_;
 wire _17742_;
 wire _17743_;
 wire _17744_;
 wire _17745_;
 wire _17746_;
 wire _17747_;
 wire _17748_;
 wire _17749_;
 wire _17750_;
 wire _17751_;
 wire _17752_;
 wire _17753_;
 wire _17754_;
 wire _17755_;
 wire _17756_;
 wire _17757_;
 wire _17758_;
 wire _17759_;
 wire _17760_;
 wire _17761_;
 wire _17762_;
 wire _17763_;
 wire _17764_;
 wire _17765_;
 wire _17766_;
 wire _17767_;
 wire _17768_;
 wire _17769_;
 wire _17770_;
 wire _17771_;
 wire _17772_;
 wire _17773_;
 wire _17774_;
 wire _17775_;
 wire _17776_;
 wire _17777_;
 wire _17778_;
 wire _17779_;
 wire _17780_;
 wire _17781_;
 wire _17782_;
 wire _17783_;
 wire _17784_;
 wire _17785_;
 wire _17786_;
 wire _17787_;
 wire _17788_;
 wire _17789_;
 wire _17790_;
 wire _17791_;
 wire _17792_;
 wire _17793_;
 wire _17794_;
 wire _17795_;
 wire _17796_;
 wire _17797_;
 wire _17798_;
 wire _17799_;
 wire _17800_;
 wire _17801_;
 wire _17802_;
 wire _17803_;
 wire _17804_;
 wire _17805_;
 wire _17806_;
 wire _17807_;
 wire _17808_;
 wire _17809_;
 wire _17810_;
 wire _17811_;
 wire _17812_;
 wire _17813_;
 wire _17814_;
 wire _17815_;
 wire _17816_;
 wire _17817_;
 wire _17818_;
 wire _17819_;
 wire _17820_;
 wire _17821_;
 wire _17822_;
 wire _17823_;
 wire _17824_;
 wire _17825_;
 wire _17826_;
 wire _17827_;
 wire _17828_;
 wire _17829_;
 wire _17830_;
 wire _17831_;
 wire _17832_;
 wire _17833_;
 wire _17834_;
 wire _17835_;
 wire _17836_;
 wire _17837_;
 wire _17838_;
 wire _17839_;
 wire _17840_;
 wire _17841_;
 wire _17842_;
 wire _17843_;
 wire _17844_;
 wire _17845_;
 wire _17846_;
 wire _17847_;
 wire _17848_;
 wire _17849_;
 wire _17850_;
 wire _17851_;
 wire _17852_;
 wire _17853_;
 wire _17854_;
 wire _17855_;
 wire _17856_;
 wire _17857_;
 wire _17858_;
 wire _17859_;
 wire _17860_;
 wire _17861_;
 wire _17862_;
 wire _17863_;
 wire _17864_;
 wire _17865_;
 wire _17866_;
 wire _17867_;
 wire _17868_;
 wire _17869_;
 wire _17870_;
 wire _17871_;
 wire _17872_;
 wire _17873_;
 wire _17874_;
 wire _17875_;
 wire _17876_;
 wire _17877_;
 wire _17878_;
 wire _17879_;
 wire _17880_;
 wire _17881_;
 wire _17882_;
 wire _17883_;
 wire _17884_;
 wire _17885_;
 wire _17886_;
 wire _17887_;
 wire _17888_;
 wire _17889_;
 wire _17890_;
 wire _17891_;
 wire _17892_;
 wire _17893_;
 wire _17894_;
 wire _17895_;
 wire _17896_;
 wire _17897_;
 wire _17898_;
 wire _17899_;
 wire _17900_;
 wire _17901_;
 wire _17902_;
 wire _17903_;
 wire _17904_;
 wire _17905_;
 wire _17906_;
 wire _17907_;
 wire _17908_;
 wire _17909_;
 wire _17910_;
 wire _17911_;
 wire _17912_;
 wire _17913_;
 wire _17914_;
 wire _17915_;
 wire _17916_;
 wire _17917_;
 wire _17918_;
 wire _17919_;
 wire _17920_;
 wire _17921_;
 wire _17922_;
 wire _17923_;
 wire _17924_;
 wire _17925_;
 wire _17926_;
 wire _17927_;
 wire _17928_;
 wire _17929_;
 wire _17930_;
 wire _17931_;
 wire _17932_;
 wire _17933_;
 wire _17934_;
 wire _17935_;
 wire _17936_;
 wire _17937_;
 wire _17938_;
 wire _17939_;
 wire _17940_;
 wire _17941_;
 wire _17942_;
 wire _17943_;
 wire _17944_;
 wire _17945_;
 wire _17946_;
 wire _17947_;
 wire _17948_;
 wire _17949_;
 wire _17950_;
 wire _17951_;
 wire _17952_;
 wire _17953_;
 wire _17954_;
 wire _17955_;
 wire _17956_;
 wire _17957_;
 wire _17958_;
 wire _17959_;
 wire _17960_;
 wire _17961_;
 wire _17962_;
 wire _17963_;
 wire _17964_;
 wire _17965_;
 wire _17966_;
 wire _17967_;
 wire _17968_;
 wire _17969_;
 wire _17970_;
 wire _17971_;
 wire _17972_;
 wire _17973_;
 wire _17974_;
 wire _17975_;
 wire _17976_;
 wire _17977_;
 wire _17978_;
 wire _17979_;
 wire _17980_;
 wire _17981_;
 wire _17982_;
 wire _17983_;
 wire _17984_;
 wire _17985_;
 wire _17986_;
 wire _17987_;
 wire _17988_;
 wire _17989_;
 wire _17990_;
 wire _17991_;
 wire _17992_;
 wire _17993_;
 wire _17994_;
 wire _17995_;
 wire _17996_;
 wire _17997_;
 wire _17998_;
 wire _17999_;
 wire _18000_;
 wire _18001_;
 wire _18002_;
 wire _18003_;
 wire _18004_;
 wire _18005_;
 wire _18006_;
 wire _18007_;
 wire _18008_;
 wire _18009_;
 wire _18010_;
 wire _18011_;
 wire _18012_;
 wire _18013_;
 wire _18014_;
 wire _18015_;
 wire _18016_;
 wire _18017_;
 wire _18018_;
 wire _18019_;
 wire _18020_;
 wire _18021_;
 wire _18022_;
 wire _18023_;
 wire _18024_;
 wire _18025_;
 wire _18026_;
 wire _18027_;
 wire _18028_;
 wire _18029_;
 wire _18030_;
 wire _18031_;
 wire _18032_;
 wire _18033_;
 wire _18034_;
 wire _18035_;
 wire _18036_;
 wire _18037_;
 wire _18038_;
 wire _18039_;
 wire _18040_;
 wire _18041_;
 wire _18042_;
 wire _18043_;
 wire _18044_;
 wire _18045_;
 wire _18046_;
 wire _18047_;
 wire _18048_;
 wire _18049_;
 wire _18050_;
 wire _18051_;
 wire _18052_;
 wire _18053_;
 wire _18054_;
 wire _18055_;
 wire _18056_;
 wire _18057_;
 wire _18058_;
 wire _18059_;
 wire _18060_;
 wire _18061_;
 wire _18062_;
 wire _18063_;
 wire _18064_;
 wire _18065_;
 wire _18066_;
 wire _18067_;
 wire _18068_;
 wire _18069_;
 wire _18070_;
 wire _18071_;
 wire _18072_;
 wire _18073_;
 wire _18074_;
 wire _18075_;
 wire _18076_;
 wire _18077_;
 wire _18078_;
 wire _18079_;
 wire _18080_;
 wire _18081_;
 wire _18082_;
 wire _18083_;
 wire _18084_;
 wire _18085_;
 wire _18086_;
 wire _18087_;
 wire _18088_;
 wire _18089_;
 wire _18090_;
 wire _18091_;
 wire _18092_;
 wire _18093_;
 wire _18094_;
 wire _18095_;
 wire _18096_;
 wire _18097_;
 wire _18098_;
 wire _18099_;
 wire _18100_;
 wire _18101_;
 wire _18102_;
 wire _18103_;
 wire net1436;
 wire net1574;
 wire _18106_;
 wire net1333;
 wire _18108_;
 wire net1440;
 wire net1383;
 wire _18111_;
 wire net1459;
 wire net1576;
 wire _18114_;
 wire _18115_;
 wire net1043;
 wire _18117_;
 wire net1252;
 wire _18119_;
 wire net1316;
 wire _18121_;
 wire net1317;
 wire net1239;
 wire _18124_;
 wire net1312;
 wire net1230;
 wire net1313;
 wire _18128_;
 wire _18129_;
 wire net1311;
 wire _18131_;
 wire net1310;
 wire _18133_;
 wire _18134_;
 wire _18135_;
 wire net1223;
 wire _18137_;
 wire _18138_;
 wire _18139_;
 wire net1307;
 wire _18141_;
 wire _18142_;
 wire _18143_;
 wire _18144_;
 wire net1299;
 wire _18146_;
 wire _18147_;
 wire _18148_;
 wire _18149_;
 wire net1296;
 wire net1215;
 wire _18152_;
 wire _18153_;
 wire _18154_;
 wire _18155_;
 wire net1214;
 wire _18157_;
 wire _18158_;
 wire _18159_;
 wire net1290;
 wire net1265;
 wire _18162_;
 wire _18163_;
 wire _18164_;
 wire _18165_;
 wire _18166_;
 wire _18167_;
 wire _18168_;
 wire _18169_;
 wire _18170_;
 wire _18171_;
 wire net1135;
 wire _18173_;
 wire _18174_;
 wire _18175_;
 wire net1102;
 wire _18177_;
 wire _18178_;
 wire _18179_;
 wire net1098;
 wire _18181_;
 wire _18182_;
 wire net1100;
 wire _18184_;
 wire _18185_;
 wire _18186_;
 wire _18187_;
 wire net1094;
 wire _18189_;
 wire _18190_;
 wire net1092;
 wire _18192_;
 wire _18193_;
 wire _18194_;
 wire _18195_;
 wire _18196_;
 wire _18197_;
 wire _18198_;
 wire _18199_;
 wire _18200_;
 wire _18201_;
 wire net1077;
 wire _18203_;
 wire _18204_;
 wire _18205_;
 wire _18206_;
 wire _18207_;
 wire net1073;
 wire _18209_;
 wire net1069;
 wire _18211_;
 wire _18212_;
 wire _18213_;
 wire _18214_;
 wire _18215_;
 wire _18216_;
 wire net1066;
 wire _18218_;
 wire _18219_;
 wire net1064;
 wire _18221_;
 wire _18222_;
 wire _18223_;
 wire _18224_;
 wire _18225_;
 wire _18226_;
 wire _18227_;
 wire net1062;
 wire _18229_;
 wire net1061;
 wire _18231_;
 wire _18232_;
 wire net1060;
 wire _18234_;
 wire _18235_;
 wire _18236_;
 wire _18237_;
 wire _18238_;
 wire _18239_;
 wire net1058;
 wire _18241_;
 wire _18242_;
 wire net1059;
 wire _18244_;
 wire net1056;
 wire _18246_;
 wire _18247_;
 wire _18248_;
 wire _18249_;
 wire net1055;
 wire _18251_;
 wire _18252_;
 wire _18253_;
 wire _18254_;
 wire net1054;
 wire _18256_;
 wire _18257_;
 wire net1053;
 wire _18259_;
 wire _18260_;
 wire _18261_;
 wire _18262_;
 wire _18263_;
 wire _18264_;
 wire _18265_;
 wire _18266_;
 wire _18267_;
 wire _18268_;
 wire _18269_;
 wire _18270_;
 wire _18271_;
 wire _18272_;
 wire _18273_;
 wire _18274_;
 wire _18275_;
 wire _18276_;
 wire _18277_;
 wire _18278_;
 wire _18279_;
 wire _18280_;
 wire _18281_;
 wire _18282_;
 wire _18283_;
 wire _18284_;
 wire _18285_;
 wire _18286_;
 wire _18287_;
 wire _18288_;
 wire _18289_;
 wire _18290_;
 wire _18291_;
 wire _18292_;
 wire _18293_;
 wire _18294_;
 wire _18295_;
 wire _18296_;
 wire _18297_;
 wire _18298_;
 wire _18299_;
 wire _18300_;
 wire _18301_;
 wire _18302_;
 wire _18303_;
 wire _18304_;
 wire _18305_;
 wire _18306_;
 wire _18307_;
 wire _18308_;
 wire _18309_;
 wire _18310_;
 wire _18311_;
 wire _18312_;
 wire _18313_;
 wire _18314_;
 wire _18315_;
 wire _18316_;
 wire _18317_;
 wire _18318_;
 wire _18319_;
 wire _18320_;
 wire _18321_;
 wire _18322_;
 wire _18323_;
 wire _18324_;
 wire _18325_;
 wire _18326_;
 wire _18327_;
 wire _18328_;
 wire _18329_;
 wire _18330_;
 wire _18331_;
 wire _18332_;
 wire _18333_;
 wire _18334_;
 wire _18335_;
 wire _18336_;
 wire _18337_;
 wire _18338_;
 wire _18339_;
 wire _18340_;
 wire _18341_;
 wire _18342_;
 wire _18343_;
 wire _18344_;
 wire _18345_;
 wire _18346_;
 wire _18347_;
 wire _18348_;
 wire _18349_;
 wire _18350_;
 wire _18351_;
 wire _18352_;
 wire _18353_;
 wire _18354_;
 wire _18355_;
 wire _18356_;
 wire _18357_;
 wire _18358_;
 wire _18359_;
 wire _18360_;
 wire _18361_;
 wire _18362_;
 wire _18363_;
 wire _18364_;
 wire _18365_;
 wire _18366_;
 wire _18367_;
 wire _18368_;
 wire _18369_;
 wire _18370_;
 wire _18371_;
 wire _18372_;
 wire _18373_;
 wire _18374_;
 wire _18375_;
 wire _18376_;
 wire _18377_;
 wire _18378_;
 wire _18379_;
 wire _18380_;
 wire _18381_;
 wire _18382_;
 wire _18383_;
 wire _18384_;
 wire _18385_;
 wire _18386_;
 wire _18387_;
 wire clknet_leaf_0_clk_i;
 wire net29;
 wire net456;
 wire core_busy_d;
 wire \core_clock_gate_i.clk_o ;
 wire \core_clock_gate_i.en_latch ;
 wire \cs_registers_i.mcycle_counter_i.counter[0] ;
 wire \cs_registers_i.mcycle_counter_i.counter[10] ;
 wire \cs_registers_i.mcycle_counter_i.counter[12] ;
 wire \cs_registers_i.mcycle_counter_i.counter[14] ;
 wire \cs_registers_i.mcycle_counter_i.counter[16] ;
 wire \cs_registers_i.mcycle_counter_i.counter[18] ;
 wire \cs_registers_i.mcycle_counter_i.counter[1] ;
 wire \cs_registers_i.mcycle_counter_i.counter[20] ;
 wire \cs_registers_i.mcycle_counter_i.counter[22] ;
 wire \cs_registers_i.mcycle_counter_i.counter[24] ;
 wire \cs_registers_i.mcycle_counter_i.counter[26] ;
 wire \cs_registers_i.mcycle_counter_i.counter[28] ;
 wire \cs_registers_i.mcycle_counter_i.counter[2] ;
 wire \cs_registers_i.mcycle_counter_i.counter[30] ;
 wire \cs_registers_i.mcycle_counter_i.counter[32] ;
 wire \cs_registers_i.mcycle_counter_i.counter[34] ;
 wire \cs_registers_i.mcycle_counter_i.counter[36] ;
 wire \cs_registers_i.mcycle_counter_i.counter[38] ;
 wire \cs_registers_i.mcycle_counter_i.counter[40] ;
 wire \cs_registers_i.mcycle_counter_i.counter[42] ;
 wire \cs_registers_i.mcycle_counter_i.counter[44] ;
 wire \cs_registers_i.mcycle_counter_i.counter[46] ;
 wire \cs_registers_i.mcycle_counter_i.counter[48] ;
 wire \cs_registers_i.mcycle_counter_i.counter[4] ;
 wire \cs_registers_i.mcycle_counter_i.counter[50] ;
 wire \cs_registers_i.mcycle_counter_i.counter[52] ;
 wire \cs_registers_i.mcycle_counter_i.counter[54] ;
 wire \cs_registers_i.mcycle_counter_i.counter[56] ;
 wire \cs_registers_i.mcycle_counter_i.counter[58] ;
 wire \cs_registers_i.mcycle_counter_i.counter[60] ;
 wire \cs_registers_i.mcycle_counter_i.counter[62] ;
 wire \cs_registers_i.mcycle_counter_i.counter[6] ;
 wire \cs_registers_i.mcycle_counter_i.counter[8] ;
 wire \cs_registers_i.mhpmcounter[2][0] ;
 wire \cs_registers_i.mhpmcounter[2][10] ;
 wire \cs_registers_i.mhpmcounter[2][12] ;
 wire \cs_registers_i.mhpmcounter[2][14] ;
 wire \cs_registers_i.mhpmcounter[2][16] ;
 wire \cs_registers_i.mhpmcounter[2][18] ;
 wire \cs_registers_i.mhpmcounter[2][1] ;
 wire \cs_registers_i.mhpmcounter[2][20] ;
 wire \cs_registers_i.mhpmcounter[2][22] ;
 wire \cs_registers_i.mhpmcounter[2][24] ;
 wire \cs_registers_i.mhpmcounter[2][26] ;
 wire \cs_registers_i.mhpmcounter[2][28] ;
 wire \cs_registers_i.mhpmcounter[2][2] ;
 wire \cs_registers_i.mhpmcounter[2][30] ;
 wire \cs_registers_i.mhpmcounter[2][32] ;
 wire \cs_registers_i.mhpmcounter[2][34] ;
 wire \cs_registers_i.mhpmcounter[2][36] ;
 wire \cs_registers_i.mhpmcounter[2][38] ;
 wire \cs_registers_i.mhpmcounter[2][40] ;
 wire \cs_registers_i.mhpmcounter[2][42] ;
 wire \cs_registers_i.mhpmcounter[2][44] ;
 wire \cs_registers_i.mhpmcounter[2][46] ;
 wire \cs_registers_i.mhpmcounter[2][48] ;
 wire \cs_registers_i.mhpmcounter[2][4] ;
 wire \cs_registers_i.mhpmcounter[2][50] ;
 wire \cs_registers_i.mhpmcounter[2][52] ;
 wire \cs_registers_i.mhpmcounter[2][54] ;
 wire \cs_registers_i.mhpmcounter[2][56] ;
 wire \cs_registers_i.mhpmcounter[2][58] ;
 wire \cs_registers_i.mhpmcounter[2][60] ;
 wire \cs_registers_i.mhpmcounter[2][62] ;
 wire \cs_registers_i.mhpmcounter[2][6] ;
 wire \cs_registers_i.mhpmcounter[2][8] ;
 wire \cs_registers_i.pc_id_i[11] ;
 wire \cs_registers_i.pc_id_i[13] ;
 wire \cs_registers_i.pc_id_i[15] ;
 wire \cs_registers_i.pc_id_i[17] ;
 wire \cs_registers_i.pc_id_i[19] ;
 wire \cs_registers_i.pc_id_i[1] ;
 wire \cs_registers_i.pc_id_i[21] ;
 wire \cs_registers_i.pc_id_i[23] ;
 wire \cs_registers_i.pc_id_i[25] ;
 wire \cs_registers_i.pc_id_i[27] ;
 wire \cs_registers_i.pc_id_i[29] ;
 wire \cs_registers_i.pc_id_i[2] ;
 wire \cs_registers_i.pc_id_i[3] ;
 wire \cs_registers_i.pc_id_i[5] ;
 wire \cs_registers_i.pc_id_i[7] ;
 wire \cs_registers_i.pc_id_i[9] ;
 wire \cs_registers_i.pc_if_i[11] ;
 wire \cs_registers_i.pc_if_i[13] ;
 wire \cs_registers_i.pc_if_i[15] ;
 wire \cs_registers_i.pc_if_i[17] ;
 wire \cs_registers_i.pc_if_i[19] ;
 wire \cs_registers_i.pc_if_i[21] ;
 wire \cs_registers_i.pc_if_i[23] ;
 wire \cs_registers_i.pc_if_i[25] ;
 wire \cs_registers_i.pc_if_i[27] ;
 wire \cs_registers_i.pc_if_i[29] ;
 wire \cs_registers_i.pc_if_i[2] ;
 wire \cs_registers_i.pc_if_i[3] ;
 wire \cs_registers_i.pc_if_i[5] ;
 wire \cs_registers_i.pc_if_i[7] ;
 wire \cs_registers_i.pc_if_i[9] ;
 wire \cs_registers_i.priv_lvl_q[0] ;
 wire \ex_block_i.alu_adder_result_ex_o[0] ;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire net11;
 wire \ex_block_i.alu_adder_result_ex_o[1] ;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ;
 wire \id_stage_i.branch_set_d ;
 wire \id_stage_i.controller_i.exc_req_d ;
 wire \id_stage_i.controller_i.illegal_insn_d ;
 wire \id_stage_i.controller_i.load_err_d ;
 wire \id_stage_i.controller_i.store_err_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ;
 wire \if_stage_i.instr_valid_id_d ;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_2_clk_i;
 wire clknet_leaf_3_clk_i;
 wire clknet_leaf_4_clk_i;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_6_clk_i;
 wire clknet_leaf_7_clk_i;
 wire clknet_leaf_8_clk_i;
 wire clknet_leaf_9_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_leaf_12_clk_i;
 wire clknet_leaf_13_clk_i;
 wire clknet_leaf_14_clk_i;
 wire clknet_leaf_15_clk_i;
 wire clknet_leaf_16_clk_i;
 wire clknet_leaf_17_clk_i;
 wire clknet_leaf_18_clk_i;
 wire clknet_leaf_19_clk_i;
 wire clknet_leaf_20_clk_i;
 wire clknet_leaf_21_clk_i;
 wire clknet_leaf_22_clk_i;
 wire clknet_leaf_23_clk_i;
 wire clknet_leaf_24_clk_i;
 wire clknet_leaf_25_clk_i;
 wire clknet_leaf_26_clk_i;
 wire clknet_leaf_27_clk_i;
 wire clknet_leaf_28_clk_i;
 wire clknet_leaf_29_clk_i;
 wire clknet_leaf_30_clk_i;
 wire clknet_leaf_31_clk_i;
 wire clknet_leaf_32_clk_i;
 wire clknet_leaf_33_clk_i;
 wire clknet_0_clk_i;
 wire clknet_2_0__leaf_clk_i;
 wire clknet_2_1__leaf_clk_i;
 wire clknet_2_2__leaf_clk_i;
 wire clknet_2_3__leaf_clk_i;
 wire clknet_level_0_1_10_clk_i;
 wire clknet_level_1_1_11_clk_i;
 wire clknet_level_2_1_12_clk_i;
 wire clknet_level_3_1_13_clk_i;
 wire clknet_level_0_1_24_clk_i;
 wire clknet_level_1_1_25_clk_i;
 wire clknet_level_2_1_26_clk_i;
 wire clknet_level_3_1_27_clk_i;
 wire clknet_level_0_1_38_clk_i;
 wire clknet_level_1_1_39_clk_i;
 wire clknet_level_2_1_310_clk_i;
 wire clknet_level_3_1_311_clk_i;
 wire clknet_level_0_1_412_clk_i;
 wire clknet_level_1_1_413_clk_i;
 wire clknet_level_2_1_414_clk_i;
 wire clknet_level_3_1_415_clk_i;
 wire clknet_level_0_1_516_clk_i;
 wire clknet_level_1_1_517_clk_i;
 wire clknet_level_2_1_518_clk_i;
 wire clknet_level_3_1_519_clk_i;
 wire clknet_level_0_1_620_clk_i;
 wire clknet_level_1_1_621_clk_i;
 wire clknet_level_2_1_622_clk_i;
 wire clknet_level_3_1_623_clk_i;
 wire clknet_level_0_1_724_clk_i;
 wire clknet_level_1_1_725_clk_i;
 wire clknet_level_2_1_726_clk_i;
 wire clknet_level_3_1_727_clk_i;
 wire clknet_level_0_1_828_clk_i;
 wire clknet_level_1_1_829_clk_i;
 wire clknet_level_2_1_830_clk_i;
 wire clknet_level_3_1_831_clk_i;
 wire clknet_level_0_1_932_clk_i;
 wire clknet_level_1_1_933_clk_i;
 wire clknet_level_2_1_934_clk_i;
 wire clknet_level_3_1_935_clk_i;
 wire clknet_level_0_1_1036_clk_i;
 wire clknet_level_1_1_1037_clk_i;
 wire clknet_level_2_1_1038_clk_i;
 wire clknet_level_3_1_1039_clk_i;
 wire clknet_level_0_1_1140_clk_i;
 wire clknet_level_1_1_1141_clk_i;
 wire clknet_level_2_1_1142_clk_i;
 wire clknet_level_3_1_1143_clk_i;
 wire clknet_level_0_1_1244_clk_i;
 wire clknet_level_1_1_1245_clk_i;
 wire clknet_level_2_1_1246_clk_i;
 wire clknet_level_3_1_1247_clk_i;
 wire clknet_level_0_1_1348_clk_i;
 wire clknet_level_1_1_1349_clk_i;
 wire clknet_level_2_1_1350_clk_i;
 wire clknet_level_3_1_1351_clk_i;
 wire clknet_level_0_1_1452_clk_i;
 wire clknet_level_1_1_1453_clk_i;
 wire clknet_level_2_1_1454_clk_i;
 wire clknet_level_3_1_1455_clk_i;
 wire clknet_level_0_1_1556_clk_i;
 wire clknet_level_1_1_1557_clk_i;
 wire clknet_level_2_1_1558_clk_i;
 wire clknet_level_3_1_1559_clk_i;
 wire clknet_level_0_1_1660_clk_i;
 wire clknet_level_1_1_1661_clk_i;
 wire clknet_level_2_1_1662_clk_i;
 wire clknet_level_3_1_1663_clk_i;
 wire clknet_level_0_1_1764_clk_i;
 wire clknet_level_1_1_1765_clk_i;
 wire clknet_level_2_1_1766_clk_i;
 wire clknet_level_3_1_1767_clk_i;
 wire clknet_level_0_1_1868_clk_i;
 wire clknet_level_1_1_1869_clk_i;
 wire clknet_level_2_1_1870_clk_i;
 wire clknet_level_3_1_1871_clk_i;
 wire clknet_level_0_1_1972_clk_i;
 wire clknet_level_1_1_1973_clk_i;
 wire clknet_level_2_1_1974_clk_i;
 wire clknet_level_3_1_1975_clk_i;
 wire clknet_level_0_1_2076_clk_i;
 wire clknet_level_1_1_2077_clk_i;
 wire clknet_level_2_1_2078_clk_i;
 wire clknet_level_3_1_2079_clk_i;
 wire clknet_level_0_1_2180_clk_i;
 wire clknet_level_1_1_2181_clk_i;
 wire clknet_level_2_1_2182_clk_i;
 wire clknet_level_3_1_2183_clk_i;
 wire clknet_level_0_1_2284_clk_i;
 wire clknet_level_1_1_2285_clk_i;
 wire clknet_level_2_1_2286_clk_i;
 wire clknet_level_3_1_2287_clk_i;
 wire clknet_level_0_1_2388_clk_i;
 wire clknet_level_1_1_2389_clk_i;
 wire clknet_level_2_1_2390_clk_i;
 wire clknet_level_3_1_2391_clk_i;
 wire clknet_level_0_1_2492_clk_i;
 wire clknet_level_1_1_2493_clk_i;
 wire clknet_level_2_1_2494_clk_i;
 wire clknet_level_3_1_2495_clk_i;
 wire clknet_level_0_1_2596_clk_i;
 wire clknet_level_1_1_2597_clk_i;
 wire clknet_level_2_1_2598_clk_i;
 wire clknet_level_3_1_2599_clk_i;
 wire clknet_level_0_1_26100_clk_i;
 wire clknet_level_1_1_26101_clk_i;
 wire clknet_level_2_1_26102_clk_i;
 wire clknet_level_3_1_26103_clk_i;
 wire clknet_level_0_1_27104_clk_i;
 wire clknet_level_1_1_27105_clk_i;
 wire clknet_level_2_1_27106_clk_i;
 wire clknet_level_3_1_27107_clk_i;
 wire clknet_level_0_1_28108_clk_i;
 wire clknet_level_1_1_28109_clk_i;
 wire clknet_level_2_1_28110_clk_i;
 wire clknet_level_3_1_28111_clk_i;
 wire clknet_level_0_1_29112_clk_i;
 wire clknet_level_1_1_29113_clk_i;
 wire clknet_level_2_1_29114_clk_i;
 wire clknet_level_3_1_29115_clk_i;
 wire clknet_level_0_1_30116_clk_i;
 wire clknet_level_1_1_30117_clk_i;
 wire clknet_level_2_1_30118_clk_i;
 wire clknet_level_3_1_30119_clk_i;
 wire clknet_level_0_1_31120_clk_i;
 wire clknet_level_1_1_31121_clk_i;
 wire clknet_level_2_1_31122_clk_i;
 wire clknet_level_3_1_31123_clk_i;
 wire clknet_level_0_1_32124_clk_i;
 wire clknet_level_1_1_32125_clk_i;
 wire clknet_level_2_1_32126_clk_i;
 wire clknet_level_3_1_32127_clk_i;
 wire clknet_level_0_1_33128_clk_i;
 wire clknet_level_1_1_33129_clk_i;
 wire clknet_level_2_1_33130_clk_i;
 wire clknet_level_3_1_33131_clk_i;
 wire clknet_level_0_1_34132_clk_i;
 wire clknet_level_1_1_34133_clk_i;
 wire clknet_level_2_1_34134_clk_i;
 wire clknet_level_3_1_34135_clk_i;
 wire \clknet_leaf_0_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_1_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_2_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_3_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_4_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_5_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_6_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_7_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_8_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_9_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_10_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_11_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_12_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_13_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_14_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_15_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_16_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_17_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_18_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_19_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_20_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_21_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_22_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_23_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_24_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_25_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_26_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_27_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_28_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_29_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_30_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_31_core_clock_gate_i.clk_o ;
 wire \clknet_0_core_clock_gate_i.clk_o ;
 wire \clknet_2_0__leaf_core_clock_gate_i.clk_o ;
 wire \clknet_2_1__leaf_core_clock_gate_i.clk_o ;
 wire \clknet_2_2__leaf_core_clock_gate_i.clk_o ;
 wire \clknet_2_3__leaf_core_clock_gate_i.clk_o ;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;

 TIEHIx1_ASAP7_75t_R _34856__807 (.H(net807));
 TIEHIx1_ASAP7_75t_R _34855__806 (.H(net806));
 TIEHIx1_ASAP7_75t_R _34854__805 (.H(net805));
 NAND2x1_ASAP7_75t_R _18393_ (.A(net317),
    .B(net314),
    .Y(_13122_));
 TIEHIx1_ASAP7_75t_R _34853__804 (.H(net804));
 NOR2x2_ASAP7_75t_R _18395_ (.A(net354),
    .B(net322),
    .Y(_13124_));
 TIEHIx1_ASAP7_75t_R _34852__803 (.H(net803));
 TIEHIx1_ASAP7_75t_R _34851__802 (.H(net802));
 INVx11_ASAP7_75t_R _18398_ (.A(net351),
    .Y(_13127_));
 TIEHIx1_ASAP7_75t_R _34850__801 (.H(net801));
 TIEHIx1_ASAP7_75t_R _34849__800 (.H(net800));
 AND2x2_ASAP7_75t_R _18401_ (.A(net348),
    .B(_00250_),
    .Y(_13130_));
 AO21x1_ASAP7_75t_R _18402_ (.A1(net312),
    .A2(_00252_),
    .B(_13130_),
    .Y(_13131_));
 CKINVDCx20_ASAP7_75t_R _18403_ (.A(net324),
    .Y(_13132_));
 AND2x6_ASAP7_75t_R _18404_ (.A(_00246_),
    .B(_13132_),
    .Y(_13133_));
 TIEHIx1_ASAP7_75t_R _34848__799 (.H(net799));
 TIEHIx1_ASAP7_75t_R _34847__798 (.H(net798));
 AND2x2_ASAP7_75t_R _18407_ (.A(net348),
    .B(_00249_),
    .Y(_13136_));
 AO21x1_ASAP7_75t_R _18408_ (.A1(net312),
    .A2(_00251_),
    .B(_13136_),
    .Y(_13137_));
 AO22x1_ASAP7_75t_R _18409_ (.A1(_13124_),
    .A2(_13131_),
    .B1(_13133_),
    .B2(_13137_),
    .Y(_13138_));
 TIEHIx1_ASAP7_75t_R _34846__797 (.H(net797));
 TIEHIx1_ASAP7_75t_R _34845__796 (.H(net796));
 TIEHIx1_ASAP7_75t_R _34844__795 (.H(net795));
 TIEHIx1_ASAP7_75t_R _34843__794 (.H(net794));
 AND2x2_ASAP7_75t_R _18414_ (.A(net348),
    .B(_01708_),
    .Y(_13143_));
 AO21x1_ASAP7_75t_R _18415_ (.A1(_00248_),
    .A2(net312),
    .B(_13143_),
    .Y(_13144_));
 CKINVDCx16_ASAP7_75t_R _18416_ (.A(net355),
    .Y(_13145_));
 TIEHIx1_ASAP7_75t_R _34842__793 (.H(net793));
 TIEHIx1_ASAP7_75t_R _34841__792 (.H(net792));
 OR3x1_ASAP7_75t_R _18419_ (.A(_00247_),
    .B(net311),
    .C(net348),
    .Y(_13148_));
 TIEHIx1_ASAP7_75t_R _34840__791 (.H(net791));
 OA211x2_ASAP7_75t_R _18421_ (.A1(net361),
    .A2(_13144_),
    .B(_13148_),
    .C(net323),
    .Y(_13150_));
 OR3x4_ASAP7_75t_R _18422_ (.A(_13122_),
    .B(_13138_),
    .C(_13150_),
    .Y(_13151_));
 TIEHIx1_ASAP7_75t_R _34839__790 (.H(net790));
 TIEHIx1_ASAP7_75t_R _34838__789 (.H(net789));
 INVx1_ASAP7_75t_R _18425_ (.A(_00263_),
    .Y(_13154_));
 TIEHIx1_ASAP7_75t_R _34837__788 (.H(net788));
 NAND2x1_ASAP7_75t_R _18427_ (.A(net348),
    .B(_00261_),
    .Y(_13156_));
 TIEHIx1_ASAP7_75t_R _34836__787 (.H(net787));
 OA211x2_ASAP7_75t_R _18429_ (.A1(net348),
    .A2(_13154_),
    .B(_13156_),
    .C(net323),
    .Y(_13158_));
 INVx1_ASAP7_75t_R _18430_ (.A(_00267_),
    .Y(_13159_));
 NAND2x1_ASAP7_75t_R _18431_ (.A(net348),
    .B(_00265_),
    .Y(_13160_));
 TIEHIx1_ASAP7_75t_R _34835__786 (.H(net786));
 OA211x2_ASAP7_75t_R _18433_ (.A1(net348),
    .A2(_13159_),
    .B(_13160_),
    .C(_13132_),
    .Y(_13162_));
 OR3x1_ASAP7_75t_R _18434_ (.A(net311),
    .B(_13158_),
    .C(_13162_),
    .Y(_13163_));
 AND2x6_ASAP7_75t_R _18435_ (.A(net311),
    .B(net322),
    .Y(_13164_));
 TIEHIx1_ASAP7_75t_R _34834__785 (.H(net785));
 TIEHIx1_ASAP7_75t_R _34833__784 (.H(net784));
 TIEHIx1_ASAP7_75t_R _34832__783 (.H(net783));
 TIEHIx1_ASAP7_75t_R _34831__782 (.H(net782));
 AND2x2_ASAP7_75t_R _18440_ (.A(net348),
    .B(_00262_),
    .Y(_13169_));
 AO21x1_ASAP7_75t_R _18441_ (.A1(net312),
    .A2(_00264_),
    .B(_13169_),
    .Y(_13170_));
 AND2x2_ASAP7_75t_R _18442_ (.A(net348),
    .B(_00266_),
    .Y(_13171_));
 AO21x1_ASAP7_75t_R _18443_ (.A1(net312),
    .A2(_00268_),
    .B(_13171_),
    .Y(_13172_));
 TIEHIx1_ASAP7_75t_R _34830__781 (.H(net781));
 CKINVDCx20_ASAP7_75t_R _18445_ (.A(_00244_),
    .Y(_13174_));
 NAND2x2_ASAP7_75t_R _18446_ (.A(net317),
    .B(_13174_),
    .Y(_13175_));
 AOI221x1_ASAP7_75t_R _18447_ (.A1(_13164_),
    .A2(_13170_),
    .B1(_13172_),
    .B2(_13124_),
    .C(_13175_),
    .Y(_13176_));
 NAND2x2_ASAP7_75t_R _18448_ (.A(_13163_),
    .B(_13176_),
    .Y(_13177_));
 TIEHIx1_ASAP7_75t_R _34829__780 (.H(net780));
 INVx1_ASAP7_75t_R _18450_ (.A(_00254_),
    .Y(_13179_));
 TIEHIx1_ASAP7_75t_R _34828__779 (.H(net779));
 NOR2x1_ASAP7_75t_R _18452_ (.A(net349),
    .B(_00256_),
    .Y(_13181_));
 AO21x1_ASAP7_75t_R _18453_ (.A1(net349),
    .A2(_13179_),
    .B(_13181_),
    .Y(_13182_));
 INVx1_ASAP7_75t_R _18454_ (.A(_00255_),
    .Y(_13183_));
 AND2x6_ASAP7_75t_R _18455_ (.A(net354),
    .B(net323),
    .Y(_13184_));
 NAND2x1_ASAP7_75t_R _18456_ (.A(net349),
    .B(_00253_),
    .Y(_13185_));
 OA211x2_ASAP7_75t_R _18457_ (.A1(net349),
    .A2(_13183_),
    .B(_13184_),
    .C(_13185_),
    .Y(_13186_));
 AOI21x1_ASAP7_75t_R _18458_ (.A1(_13164_),
    .A2(_13182_),
    .B(_13186_),
    .Y(_13187_));
 TIEHIx1_ASAP7_75t_R _34827__778 (.H(net778));
 AND3x1_ASAP7_75t_R _18460_ (.A(net361),
    .B(net349),
    .C(_00257_),
    .Y(_13189_));
 AND2x6_ASAP7_75t_R _18461_ (.A(net355),
    .B(net313),
    .Y(_13190_));
 OR3x1_ASAP7_75t_R _18462_ (.A(net323),
    .B(net317),
    .C(_13174_),
    .Y(_13191_));
 AO21x1_ASAP7_75t_R _18463_ (.A1(_00259_),
    .A2(_13190_),
    .B(_13191_),
    .Y(_13192_));
 AND2x2_ASAP7_75t_R _18464_ (.A(net349),
    .B(_00258_),
    .Y(_13193_));
 AO21x1_ASAP7_75t_R _18465_ (.A1(net312),
    .A2(_00260_),
    .B(_13193_),
    .Y(_13194_));
 AND2x2_ASAP7_75t_R _18466_ (.A(net311),
    .B(_13194_),
    .Y(_13195_));
 OA33x2_ASAP7_75t_R _18467_ (.A1(net317),
    .A2(_13174_),
    .A3(_13187_),
    .B1(_13189_),
    .B2(_13192_),
    .B3(_13195_),
    .Y(_13196_));
 TIEHIx1_ASAP7_75t_R _34826__777 (.H(net777));
 INVx1_ASAP7_75t_R _18469_ (.A(_00270_),
    .Y(_13198_));
 TIEHIx1_ASAP7_75t_R _34825__776 (.H(net776));
 NOR2x1_ASAP7_75t_R _18471_ (.A(net349),
    .B(_00272_),
    .Y(_13200_));
 AO21x1_ASAP7_75t_R _18472_ (.A1(net349),
    .A2(_13198_),
    .B(_13200_),
    .Y(_13201_));
 INVx1_ASAP7_75t_R _18473_ (.A(_00276_),
    .Y(_13202_));
 NAND2x1_ASAP7_75t_R _18474_ (.A(net349),
    .B(_00274_),
    .Y(_13203_));
 OA211x2_ASAP7_75t_R _18475_ (.A1(net349),
    .A2(_13202_),
    .B(_13124_),
    .C(_13203_),
    .Y(_13204_));
 AO21x1_ASAP7_75t_R _18476_ (.A1(_13164_),
    .A2(_13201_),
    .B(_13204_),
    .Y(_13205_));
 TIEHIx1_ASAP7_75t_R _34824__775 (.H(net775));
 TIEHIx1_ASAP7_75t_R _34823__774 (.H(net774));
 NAND2x1_ASAP7_75t_R _18479_ (.A(net349),
    .B(_00273_),
    .Y(_13208_));
 TIEHIx1_ASAP7_75t_R _34822__773 (.H(net773));
 NAND2x1_ASAP7_75t_R _18481_ (.A(net312),
    .B(_00275_),
    .Y(_13210_));
 NAND2x1_ASAP7_75t_R _18482_ (.A(net349),
    .B(_00269_),
    .Y(_13211_));
 NAND2x1_ASAP7_75t_R _18483_ (.A(net312),
    .B(_00271_),
    .Y(_13212_));
 TIEHIx1_ASAP7_75t_R _34821__772 (.H(net772));
 AO33x2_ASAP7_75t_R _18485_ (.A1(_13133_),
    .A2(_13208_),
    .A3(_13210_),
    .B1(_13211_),
    .B2(_13212_),
    .B3(_13184_),
    .Y(_13214_));
 NOR2x2_ASAP7_75t_R _18486_ (.A(net317),
    .B(net314),
    .Y(_13215_));
 OAI21x1_ASAP7_75t_R _18487_ (.A1(_13205_),
    .A2(_13214_),
    .B(_13215_),
    .Y(_13216_));
 AND4x2_ASAP7_75t_R _18488_ (.A(_13151_),
    .B(_13177_),
    .C(_13196_),
    .D(_13216_),
    .Y(_13217_));
 NAND2x2_ASAP7_75t_R _18489_ (.A(_01608_),
    .B(_01609_),
    .Y(_13218_));
 OR2x4_ASAP7_75t_R _18490_ (.A(_00277_),
    .B(_13218_),
    .Y(_13219_));
 INVx1_ASAP7_75t_R _18491_ (.A(_01609_),
    .Y(_13220_));
 INVx1_ASAP7_75t_R _18492_ (.A(_00277_),
    .Y(_13221_));
 AO211x2_ASAP7_75t_R _18493_ (.A1(_18336_),
    .A2(_13220_),
    .B(_01608_),
    .C(_13221_),
    .Y(_13222_));
 AND2x6_ASAP7_75t_R _18494_ (.A(_13219_),
    .B(_13222_),
    .Y(_13223_));
 TIEHIx1_ASAP7_75t_R _34820__771 (.H(net771));
 TIEHIx1_ASAP7_75t_R _34819__770 (.H(net770));
 TIEHIx1_ASAP7_75t_R _34818__769 (.H(net769));
 CKINVDCx6p67_ASAP7_75t_R _18498_ (.A(_01317_),
    .Y(_13227_));
 NAND2x2_ASAP7_75t_R _18499_ (.A(_01713_),
    .B(_13227_),
    .Y(_13228_));
 TIEHIx1_ASAP7_75t_R _34817__768 (.H(net768));
 CKINVDCx5p33_ASAP7_75t_R _18501_ (.A(_01746_),
    .Y(_13230_));
 TIEHIx1_ASAP7_75t_R _34816__767 (.H(net767));
 TIEHIx1_ASAP7_75t_R _34815__766 (.H(net766));
 TIEHIx1_ASAP7_75t_R _34814__765 (.H(net765));
 NOR3x2_ASAP7_75t_R _18505_ (.B(_00163_),
    .C(_00175_),
    .Y(_13234_),
    .A(_00278_));
 AND3x4_ASAP7_75t_R _18506_ (.A(_00172_),
    .B(_13230_),
    .C(_13234_),
    .Y(_13235_));
 TIEHIx1_ASAP7_75t_R _34813__764 (.H(net764));
 TIEHIx1_ASAP7_75t_R _34812__763 (.H(net763));
 INVx5_ASAP7_75t_R _18509_ (.A(_00175_),
    .Y(_13238_));
 AND4x2_ASAP7_75t_R _18510_ (.A(_00278_),
    .B(_00279_),
    .C(_00172_),
    .D(_13238_),
    .Y(_13239_));
 TIEHIx1_ASAP7_75t_R _34811__762 (.H(net762));
 TIEHIx1_ASAP7_75t_R _34810__761 (.H(net761));
 TIEHIx1_ASAP7_75t_R _34809__760 (.H(net760));
 TIEHIx1_ASAP7_75t_R _34808__759 (.H(net759));
 TIEHIx1_ASAP7_75t_R _34807__758 (.H(net758));
 NAND2x2_ASAP7_75t_R _18516_ (.A(_00165_),
    .B(_00168_),
    .Y(_13245_));
 NOR2x1_ASAP7_75t_R _18517_ (.A(_00278_),
    .B(_00172_),
    .Y(_13246_));
 OR5x2_ASAP7_75t_R _18518_ (.A(_00163_),
    .B(_00175_),
    .C(_01746_),
    .D(_13245_),
    .E(_13246_),
    .Y(_13247_));
 AOI211x1_ASAP7_75t_R _18519_ (.A1(_13228_),
    .A2(_13235_),
    .B(_13239_),
    .C(_13247_),
    .Y(_13248_));
 AOI21x1_ASAP7_75t_R _18520_ (.A1(_01713_),
    .A2(_13227_),
    .B(_00165_),
    .Y(_13249_));
 NAND2x1_ASAP7_75t_R _18521_ (.A(_13235_),
    .B(_13249_),
    .Y(_13250_));
 TIEHIx1_ASAP7_75t_R _34806__757 (.H(net757));
 AND2x6_ASAP7_75t_R _18523_ (.A(_00165_),
    .B(_00168_),
    .Y(_13252_));
 AND4x2_ASAP7_75t_R _18524_ (.A(_00172_),
    .B(_13230_),
    .C(_13234_),
    .D(_13252_),
    .Y(_13253_));
 NAND2x1_ASAP7_75t_R _18525_ (.A(_13228_),
    .B(_13253_),
    .Y(_13254_));
 INVx2_ASAP7_75t_R _18526_ (.A(_00278_),
    .Y(_13255_));
 INVx3_ASAP7_75t_R _18527_ (.A(_00168_),
    .Y(_13256_));
 OR5x1_ASAP7_75t_R _18528_ (.A(_13255_),
    .B(_00163_),
    .C(_13256_),
    .D(_00172_),
    .E(_01746_),
    .Y(_13257_));
 OA211x2_ASAP7_75t_R _18529_ (.A1(_00165_),
    .A2(_13257_),
    .B(_13222_),
    .C(_13219_),
    .Y(_13258_));
 NOR2x2_ASAP7_75t_R _18530_ (.A(_00163_),
    .B(_01746_),
    .Y(_13259_));
 AND2x2_ASAP7_75t_R _18531_ (.A(_13252_),
    .B(_13259_),
    .Y(_13260_));
 CKINVDCx9p33_ASAP7_75t_R _18532_ (.A(_00281_),
    .Y(_13261_));
 TIEHIx1_ASAP7_75t_R _34805__756 (.H(net756));
 AND2x4_ASAP7_75t_R _18534_ (.A(_00279_),
    .B(_00282_),
    .Y(_13263_));
 AND2x2_ASAP7_75t_R _18535_ (.A(_13261_),
    .B(_13263_),
    .Y(_13264_));
 NOR2x2_ASAP7_75t_R _18536_ (.A(_00163_),
    .B(_00165_),
    .Y(_13265_));
 AND2x2_ASAP7_75t_R _18537_ (.A(_00278_),
    .B(_00175_),
    .Y(_13266_));
 AND5x2_ASAP7_75t_R _18538_ (.A(_13256_),
    .B(_00172_),
    .C(_13230_),
    .D(_13265_),
    .E(_13266_),
    .Y(_13267_));
 AOI22x1_ASAP7_75t_R _18539_ (.A1(_13239_),
    .A2(_13260_),
    .B1(_13264_),
    .B2(_13267_),
    .Y(_13268_));
 AND4x2_ASAP7_75t_R _18540_ (.A(_13250_),
    .B(_13254_),
    .C(_13258_),
    .D(_13268_),
    .Y(_13269_));
 NAND2x2_ASAP7_75t_R _18541_ (.A(_13219_),
    .B(_13222_),
    .Y(_13270_));
 INVx3_ASAP7_75t_R _18542_ (.A(_00165_),
    .Y(_13271_));
 INVx2_ASAP7_75t_R _18543_ (.A(_00163_),
    .Y(_13272_));
 INVx5_ASAP7_75t_R _18544_ (.A(_00172_),
    .Y(_13273_));
 AND5x2_ASAP7_75t_R _18545_ (.A(_00278_),
    .B(_13272_),
    .C(_00168_),
    .D(_13273_),
    .E(_13230_),
    .Y(_13274_));
 AND2x2_ASAP7_75t_R _18546_ (.A(_13271_),
    .B(_13274_),
    .Y(_13275_));
 TIEHIx1_ASAP7_75t_R _34804__755 (.H(net755));
 AND3x1_ASAP7_75t_R _18548_ (.A(_00172_),
    .B(_13230_),
    .C(_13265_),
    .Y(_13277_));
 NOR2x1_ASAP7_75t_R _18549_ (.A(_00278_),
    .B(_00175_),
    .Y(_13278_));
 AO31x2_ASAP7_75t_R _18550_ (.A1(_13261_),
    .A2(_13263_),
    .A3(_13266_),
    .B(_13278_),
    .Y(_13279_));
 AND4x2_ASAP7_75t_R _18551_ (.A(_00168_),
    .B(_00172_),
    .C(_13230_),
    .D(_13234_),
    .Y(_13280_));
 AO32x2_ASAP7_75t_R _18552_ (.A1(_13256_),
    .A2(_13277_),
    .A3(_13279_),
    .B1(_13280_),
    .B2(_13249_),
    .Y(_13281_));
 OR3x1_ASAP7_75t_R _18553_ (.A(_13270_),
    .B(_13275_),
    .C(_13281_),
    .Y(_13282_));
 INVx3_ASAP7_75t_R _18554_ (.A(_18336_),
    .Y(_13283_));
 INVx1_ASAP7_75t_R _18555_ (.A(_01608_),
    .Y(_13284_));
 OA211x2_ASAP7_75t_R _18556_ (.A1(_13283_),
    .A2(_01609_),
    .B(_13284_),
    .C(_00277_),
    .Y(_13285_));
 NOR2x1_ASAP7_75t_R _18557_ (.A(_00277_),
    .B(_13218_),
    .Y(_13286_));
 AO211x2_ASAP7_75t_R _18558_ (.A1(_13271_),
    .A2(_13274_),
    .B(_13285_),
    .C(_13286_),
    .Y(_13287_));
 AND2x2_ASAP7_75t_R _18559_ (.A(_13228_),
    .B(_13253_),
    .Y(_13288_));
 AO211x2_ASAP7_75t_R _18560_ (.A1(_13250_),
    .A2(_13268_),
    .B(_13287_),
    .C(_13288_),
    .Y(_13289_));
 AND4x1_ASAP7_75t_R _18561_ (.A(_13256_),
    .B(_00172_),
    .C(_13230_),
    .D(_13265_),
    .Y(_13290_));
 AOI22x1_ASAP7_75t_R _18562_ (.A1(_13279_),
    .A2(_13290_),
    .B1(_13280_),
    .B2(_13249_),
    .Y(_13291_));
 TIEHIx1_ASAP7_75t_R _34803__754 (.H(net754));
 OA33x2_ASAP7_75t_R _18564_ (.A1(_00184_),
    .A2(_13269_),
    .A3(_13282_),
    .B1(_13289_),
    .B2(_13291_),
    .B3(_00385_),
    .Y(_13293_));
 TIEHIx1_ASAP7_75t_R _34802__753 (.H(net753));
 TIEHIx1_ASAP7_75t_R _34801__752 (.H(net752));
 AND2x2_ASAP7_75t_R _18567_ (.A(_13235_),
    .B(_13249_),
    .Y(_13296_));
 AO32x1_ASAP7_75t_R _18568_ (.A1(_13239_),
    .A2(_13252_),
    .A3(_13259_),
    .B1(_13264_),
    .B2(_13267_),
    .Y(_13297_));
 OR4x2_ASAP7_75t_R _18569_ (.A(_13296_),
    .B(_13288_),
    .C(_13287_),
    .D(_13297_),
    .Y(_13298_));
 NAND2x2_ASAP7_75t_R _18570_ (.A(_13223_),
    .B(_13248_),
    .Y(_13299_));
 OA21x2_ASAP7_75t_R _18571_ (.A1(_01745_),
    .A2(_13298_),
    .B(_13299_),
    .Y(_13300_));
 AO32x2_ASAP7_75t_R _18572_ (.A1(_13217_),
    .A2(_13223_),
    .A3(_13248_),
    .B1(_13293_),
    .B2(_13300_),
    .Y(_13301_));
 CKINVDCx10_ASAP7_75t_R _18573_ (.A(_13301_),
    .Y(_13302_));
 TIEHIx1_ASAP7_75t_R _34800__751 (.H(net751));
 TIEHIx1_ASAP7_75t_R _34799__750 (.H(net750));
 TIEHIx1_ASAP7_75t_R _34798__749 (.H(net749));
 TIEHIx1_ASAP7_75t_R _34797__748 (.H(net748));
 TIEHIx1_ASAP7_75t_R _34796__747 (.H(net747));
 INVx2_ASAP7_75t_R _18579_ (.A(_01743_),
    .Y(_13306_));
 TIEHIx1_ASAP7_75t_R _34795__746 (.H(net746));
 TIEHIx1_ASAP7_75t_R _34794__745 (.H(net745));
 TIEHIx1_ASAP7_75t_R _34793__744 (.H(net744));
 TIEHIx1_ASAP7_75t_R _34792__743 (.H(net743));
 AND4x2_ASAP7_75t_R _18584_ (.A(_00280_),
    .B(_01740_),
    .C(_01741_),
    .D(_01742_),
    .Y(_13311_));
 TIEHIx1_ASAP7_75t_R _34791__742 (.H(net742));
 AND4x2_ASAP7_75t_R _18586_ (.A(_00283_),
    .B(_01739_),
    .C(_13306_),
    .D(_13311_),
    .Y(_13313_));
 TIEHIx1_ASAP7_75t_R _34790__741 (.H(net741));
 TIEHIx1_ASAP7_75t_R _34789__740 (.H(net740));
 AND5x2_ASAP7_75t_R _18589_ (.A(_00278_),
    .B(_13272_),
    .C(_13273_),
    .D(_13230_),
    .E(_13252_),
    .Y(_13316_));
 AND2x6_ASAP7_75t_R _18590_ (.A(_13238_),
    .B(_13316_),
    .Y(_13317_));
 NAND2x2_ASAP7_75t_R _18591_ (.A(_13313_),
    .B(_13317_),
    .Y(_13318_));
 TIEHIx1_ASAP7_75t_R _34788__739 (.H(net739));
 TIEHIx1_ASAP7_75t_R _34787__738 (.H(net738));
 TIEHIx1_ASAP7_75t_R _34786__737 (.H(net737));
 TIEHIx1_ASAP7_75t_R _34785__736 (.H(net736));
 CKINVDCx6p67_ASAP7_75t_R _18596_ (.A(_00282_),
    .Y(_13323_));
 TIEHIx1_ASAP7_75t_R _34784__735 (.H(net735));
 CKINVDCx9p33_ASAP7_75t_R _18598_ (.A(_00279_),
    .Y(_13325_));
 TIEHIx1_ASAP7_75t_R _34783__734 (.H(net734));
 NAND2x2_ASAP7_75t_R _18600_ (.A(_13325_),
    .B(_00281_),
    .Y(_13327_));
 AND2x4_ASAP7_75t_R _18601_ (.A(_01713_),
    .B(_13227_),
    .Y(_13328_));
 AND2x6_ASAP7_75t_R _18602_ (.A(_13328_),
    .B(_13253_),
    .Y(_13329_));
 OA21x2_ASAP7_75t_R _18603_ (.A1(_13323_),
    .A2(_13327_),
    .B(_13329_),
    .Y(_13330_));
 TIEHIx1_ASAP7_75t_R _34782__733 (.H(net733));
 AND2x2_ASAP7_75t_R _18605_ (.A(_00283_),
    .B(_01743_),
    .Y(_13332_));
 AND4x1_ASAP7_75t_R _18606_ (.A(_13325_),
    .B(_01739_),
    .C(_13311_),
    .D(_13332_),
    .Y(_13333_));
 TIEHIx1_ASAP7_75t_R _34781__732 (.H(net732));
 NOR2x2_ASAP7_75t_R _18608_ (.A(_00281_),
    .B(_00282_),
    .Y(_13335_));
 OA211x2_ASAP7_75t_R _18609_ (.A1(_00175_),
    .A2(_13333_),
    .B(_13335_),
    .C(_13316_),
    .Y(_13336_));
 TIEHIx1_ASAP7_75t_R _34780__731 (.H(net731));
 OA211x2_ASAP7_75t_R _18611_ (.A1(_13325_),
    .A2(_01739_),
    .B(_13311_),
    .C(_13332_),
    .Y(_13338_));
 TIEHIx1_ASAP7_75t_R _34779__730 (.H(net730));
 OA21x2_ASAP7_75t_R _18613_ (.A1(_00279_),
    .A2(_13311_),
    .B(_00175_),
    .Y(_13340_));
 AO21x1_ASAP7_75t_R _18614_ (.A1(_13238_),
    .A2(_13338_),
    .B(_13340_),
    .Y(_13341_));
 AND4x2_ASAP7_75t_R _18615_ (.A(_13261_),
    .B(_00282_),
    .C(_13316_),
    .D(_13341_),
    .Y(_13342_));
 OR3x1_ASAP7_75t_R _18616_ (.A(_13330_),
    .B(_13336_),
    .C(_13342_),
    .Y(_13343_));
 NAND2x2_ASAP7_75t_R _18617_ (.A(_00279_),
    .B(_00282_),
    .Y(_13344_));
 NAND2x2_ASAP7_75t_R _18618_ (.A(_13344_),
    .B(_13267_),
    .Y(_13345_));
 OA21x2_ASAP7_75t_R _18619_ (.A1(_00278_),
    .A2(_13238_),
    .B(_00172_),
    .Y(_13346_));
 AO21x1_ASAP7_75t_R _18620_ (.A1(_13256_),
    .A2(_13266_),
    .B(_13278_),
    .Y(_13347_));
 AO221x1_ASAP7_75t_R _18621_ (.A1(_13260_),
    .A2(_13346_),
    .B1(_13347_),
    .B2(_13277_),
    .C(_13274_),
    .Y(_13348_));
 NAND2x2_ASAP7_75t_R _18622_ (.A(_13345_),
    .B(_13348_),
    .Y(_13349_));
 NAND2x2_ASAP7_75t_R _18623_ (.A(_13261_),
    .B(_00282_),
    .Y(_13350_));
 OA21x2_ASAP7_75t_R _18624_ (.A1(_00282_),
    .A2(_13327_),
    .B(_13350_),
    .Y(_13351_));
 NAND2x1_ASAP7_75t_R _18625_ (.A(_00279_),
    .B(_00281_),
    .Y(_13352_));
 NOR2x1_ASAP7_75t_R _18626_ (.A(_00279_),
    .B(_00281_),
    .Y(_13353_));
 OAI21x1_ASAP7_75t_R _18627_ (.A1(_13323_),
    .A2(_13311_),
    .B(_13353_),
    .Y(_13354_));
 AND4x1_ASAP7_75t_R _18628_ (.A(_00175_),
    .B(_13316_),
    .C(_13352_),
    .D(_13354_),
    .Y(_13355_));
 AO21x2_ASAP7_75t_R _18629_ (.A1(_13329_),
    .A2(_13351_),
    .B(_13355_),
    .Y(_13356_));
 TIEHIx1_ASAP7_75t_R _34778__729 (.H(net729));
 NAND2x1_ASAP7_75t_R _18631_ (.A(_00283_),
    .B(_13311_),
    .Y(_13358_));
 XOR2x1_ASAP7_75t_R _18632_ (.A(_00279_),
    .Y(_13359_),
    .B(_00281_));
 AND2x2_ASAP7_75t_R _18633_ (.A(_00282_),
    .B(_01743_),
    .Y(_13360_));
 NOR2x1_ASAP7_75t_R _18634_ (.A(_01739_),
    .B(_13360_),
    .Y(_13361_));
 AO21x1_ASAP7_75t_R _18635_ (.A1(_01743_),
    .A2(_13359_),
    .B(_13361_),
    .Y(_13362_));
 OA21x2_ASAP7_75t_R _18636_ (.A1(_13358_),
    .A2(_13362_),
    .B(_13317_),
    .Y(_13363_));
 OR3x4_ASAP7_75t_R _18637_ (.A(_13349_),
    .B(_13356_),
    .C(_13363_),
    .Y(_13364_));
 TIEHIx1_ASAP7_75t_R _34777__728 (.H(net728));
 OA21x2_ASAP7_75t_R _18639_ (.A1(_13325_),
    .A2(_00281_),
    .B(_00282_),
    .Y(_13366_));
 AND3x1_ASAP7_75t_R _18640_ (.A(_00282_),
    .B(_01739_),
    .C(_13353_),
    .Y(_13367_));
 AND2x2_ASAP7_75t_R _18641_ (.A(_13323_),
    .B(_01739_),
    .Y(_13368_));
 INVx3_ASAP7_75t_R _18642_ (.A(_01739_),
    .Y(_13369_));
 AND2x2_ASAP7_75t_R _18643_ (.A(_13369_),
    .B(_13263_),
    .Y(_13370_));
 OA21x2_ASAP7_75t_R _18644_ (.A1(_13368_),
    .A2(_13370_),
    .B(_00281_),
    .Y(_13371_));
 AND2x2_ASAP7_75t_R _18645_ (.A(_13311_),
    .B(_13332_),
    .Y(_13372_));
 OA211x2_ASAP7_75t_R _18646_ (.A1(_13367_),
    .A2(_13371_),
    .B(_13317_),
    .C(_13372_),
    .Y(_13373_));
 AO22x1_ASAP7_75t_R _18647_ (.A1(_00281_),
    .A2(_13323_),
    .B1(_13311_),
    .B2(_13367_),
    .Y(_13374_));
 AND3x1_ASAP7_75t_R _18648_ (.A(_00175_),
    .B(_13316_),
    .C(_13374_),
    .Y(_13375_));
 AOI211x1_ASAP7_75t_R _18649_ (.A1(_13329_),
    .A2(_13366_),
    .B(_13373_),
    .C(_13375_),
    .Y(_13376_));
 AO22x1_ASAP7_75t_R _18650_ (.A1(_13261_),
    .A2(_13369_),
    .B1(_01743_),
    .B2(_13323_),
    .Y(_13377_));
 AND2x2_ASAP7_75t_R _18651_ (.A(_00279_),
    .B(_13377_),
    .Y(_13378_));
 AOI21x1_ASAP7_75t_R _18652_ (.A1(_13327_),
    .A2(_13360_),
    .B(_01739_),
    .Y(_13379_));
 OA31x2_ASAP7_75t_R _18653_ (.A1(_13358_),
    .A2(_13378_),
    .A3(_13379_),
    .B1(_13317_),
    .Y(_13380_));
 AND2x2_ASAP7_75t_R _18654_ (.A(_00279_),
    .B(_13323_),
    .Y(_13381_));
 OR2x2_ASAP7_75t_R _18655_ (.A(_00279_),
    .B(_00281_),
    .Y(_13382_));
 NOR3x1_ASAP7_75t_R _18656_ (.A(_13323_),
    .B(_13311_),
    .C(_13382_),
    .Y(_13383_));
 OA211x2_ASAP7_75t_R _18657_ (.A1(_13381_),
    .A2(_13383_),
    .B(_00175_),
    .C(_13316_),
    .Y(_13384_));
 OR2x2_ASAP7_75t_R _18658_ (.A(_13384_),
    .B(_13329_),
    .Y(_13385_));
 NOR3x2_ASAP7_75t_R _18659_ (.B(_13380_),
    .C(_13385_),
    .Y(_13386_),
    .A(_13349_));
 OA31x2_ASAP7_75t_R _18660_ (.A1(_13343_),
    .A2(_13364_),
    .A3(_13376_),
    .B1(_13386_),
    .Y(_13387_));
 TIEHIx1_ASAP7_75t_R _34776__727 (.H(net727));
 XNOR2x1_ASAP7_75t_R _18662_ (.B(_13387_),
    .Y(_13389_),
    .A(_13301_));
 TIEHIx1_ASAP7_75t_R _34775__726 (.H(net726));
 TIEHIx1_ASAP7_75t_R _34774__725 (.H(net725));
 CKINVDCx20_ASAP7_75t_R _18665_ (.A(net364),
    .Y(_13392_));
 TIEHIx1_ASAP7_75t_R _34773__724 (.H(net724));
 TIEHIx1_ASAP7_75t_R _34772__723 (.H(net723));
 TIEHIx1_ASAP7_75t_R _34771__722 (.H(net722));
 TIEHIx1_ASAP7_75t_R _34770__721 (.H(net721));
 CKINVDCx20_ASAP7_75t_R _18670_ (.A(net370),
    .Y(_13397_));
 TIEHIx1_ASAP7_75t_R _34769__720 (.H(net720));
 TIEHIx1_ASAP7_75t_R _34768__719 (.H(net719));
 TIEHIx1_ASAP7_75t_R _34767__718 (.H(net718));
 TIEHIx1_ASAP7_75t_R _34766__717 (.H(net717));
 TIEHIx1_ASAP7_75t_R _34765__716 (.H(net716));
 INVx1_ASAP7_75t_R _18676_ (.A(_00259_),
    .Y(_13403_));
 TIEHIx1_ASAP7_75t_R _34764__715 (.H(net715));
 TIEHIx1_ASAP7_75t_R _34763__714 (.H(net714));
 TIEHIx1_ASAP7_75t_R _34762__713 (.H(net713));
 TIEHIx1_ASAP7_75t_R _34761__712 (.H(net712));
 TIEHIx1_ASAP7_75t_R _34760__711 (.H(net711));
 TIEHIx1_ASAP7_75t_R _34759__710 (.H(net710));
 TIEHIx1_ASAP7_75t_R _34758__709 (.H(net709));
 TIEHIx1_ASAP7_75t_R _34757__708 (.H(net708));
 TIEHIx1_ASAP7_75t_R _34756__707 (.H(net707));
 NAND2x1_ASAP7_75t_R _18686_ (.A(_00257_),
    .B(net382),
    .Y(_13413_));
 TIEHIx1_ASAP7_75t_R _34755__706 (.H(net706));
 TIEHIx1_ASAP7_75t_R _34754__705 (.H(net705));
 TIEHIx1_ASAP7_75t_R _34753__704 (.H(net704));
 TIEHIx1_ASAP7_75t_R _34752__703 (.H(net703));
 OA211x2_ASAP7_75t_R _18691_ (.A1(_13403_),
    .A2(net382),
    .B(_13413_),
    .C(net404),
    .Y(_13418_));
 INVx1_ASAP7_75t_R _18692_ (.A(_00260_),
    .Y(_13419_));
 TIEHIx1_ASAP7_75t_R _34751__702 (.H(net702));
 TIEHIx1_ASAP7_75t_R _34750__701 (.H(net701));
 TIEHIx1_ASAP7_75t_R _34749__700 (.H(net700));
 NAND2x1_ASAP7_75t_R _18696_ (.A(_00258_),
    .B(net382),
    .Y(_13423_));
 INVx13_ASAP7_75t_R _18697_ (.A(net407),
    .Y(_13424_));
 TIEHIx1_ASAP7_75t_R _34748__699 (.H(net699));
 TIEHIx1_ASAP7_75t_R _34747__698 (.H(net698));
 OA211x2_ASAP7_75t_R _18700_ (.A1(_13419_),
    .A2(net382),
    .B(_13423_),
    .C(net305),
    .Y(_13427_));
 OR3x1_ASAP7_75t_R _18701_ (.A(net368),
    .B(_13418_),
    .C(_13427_),
    .Y(_13428_));
 TIEHIx1_ASAP7_75t_R _34746__697 (.H(net697));
 TIEHIx1_ASAP7_75t_R _34745__696 (.H(net696));
 TIEHIx1_ASAP7_75t_R _34744__695 (.H(net695));
 TIEHIx1_ASAP7_75t_R _34743__694 (.H(net694));
 INVx13_ASAP7_75t_R _18706_ (.A(net377),
    .Y(_13433_));
 TIEHIx1_ASAP7_75t_R _34742__693 (.H(net693));
 TIEHIx1_ASAP7_75t_R _34741__692 (.H(net692));
 TIEHIx1_ASAP7_75t_R _34740__691 (.H(net691));
 TIEHIx1_ASAP7_75t_R _34739__690 (.H(net690));
 TIEHIx1_ASAP7_75t_R _34738__689 (.H(net689));
 TIEHIx1_ASAP7_75t_R _34737__688 (.H(net688));
 AND2x2_ASAP7_75t_R _18713_ (.A(_00249_),
    .B(net382),
    .Y(_13440_));
 AO21x1_ASAP7_75t_R _18714_ (.A1(_00251_),
    .A2(net303),
    .B(_13440_),
    .Y(_13441_));
 TIEHIx1_ASAP7_75t_R _34736__687 (.H(net687));
 TIEHIx1_ASAP7_75t_R _34735__686 (.H(net686));
 TIEHIx1_ASAP7_75t_R _34734__685 (.H(net685));
 TIEHIx1_ASAP7_75t_R _34733__684 (.H(net684));
 TIEHIx1_ASAP7_75t_R _34702__683 (.H(net683));
 TIEHIx1_ASAP7_75t_R _34701__682 (.H(net682));
 AND2x2_ASAP7_75t_R _18721_ (.A(_00250_),
    .B(net382),
    .Y(_13448_));
 AO21x1_ASAP7_75t_R _18722_ (.A1(_00252_),
    .A2(net303),
    .B(_13448_),
    .Y(_13449_));
 OA21x2_ASAP7_75t_R _18723_ (.A1(net404),
    .A2(_13449_),
    .B(net368),
    .Y(_13450_));
 OAI21x1_ASAP7_75t_R _18724_ (.A1(net305),
    .A2(_13441_),
    .B(_13450_),
    .Y(_13451_));
 TIEHIx1_ASAP7_75t_R _34700__681 (.H(net681));
 TIEHIx1_ASAP7_75t_R _34699__680 (.H(net680));
 TIEHIx1_ASAP7_75t_R _34698__679 (.H(net679));
 TIEHIx1_ASAP7_75t_R _34697__678 (.H(net678));
 NAND2x1_ASAP7_75t_R _18729_ (.A(_00256_),
    .B(net305),
    .Y(_13456_));
 OA211x2_ASAP7_75t_R _18730_ (.A1(_13183_),
    .A2(net305),
    .B(net303),
    .C(_13456_),
    .Y(_13457_));
 TIEHIx1_ASAP7_75t_R _34696__677 (.H(net677));
 TIEHIx1_ASAP7_75t_R _34695__676 (.H(net676));
 TIEHIx1_ASAP7_75t_R _34694__675 (.H(net675));
 TIEHIx1_ASAP7_75t_R _34693__674 (.H(net674));
 TIEHIx1_ASAP7_75t_R _34692__673 (.H(net673));
 NAND2x1_ASAP7_75t_R _18736_ (.A(_00253_),
    .B(net404),
    .Y(_13463_));
 OA211x2_ASAP7_75t_R _18737_ (.A1(_13179_),
    .A2(net404),
    .B(net382),
    .C(_13463_),
    .Y(_13464_));
 OR3x1_ASAP7_75t_R _18738_ (.A(net368),
    .B(_13457_),
    .C(_13464_),
    .Y(_13465_));
 INVx1_ASAP7_75t_R _18739_ (.A(_00248_),
    .Y(_13466_));
 TIEHIx1_ASAP7_75t_R _34691__672 (.H(net672));
 TIEHIx1_ASAP7_75t_R _34690__671 (.H(net671));
 NAND2x1_ASAP7_75t_R _18742_ (.A(net382),
    .B(_01708_),
    .Y(_13469_));
 OA211x2_ASAP7_75t_R _18743_ (.A1(_13466_),
    .A2(net382),
    .B(_13469_),
    .C(net305),
    .Y(_13470_));
 NAND2x2_ASAP7_75t_R _18744_ (.A(net409),
    .B(net303),
    .Y(_13471_));
 OAI21x1_ASAP7_75t_R _18745_ (.A1(_00247_),
    .A2(_13471_),
    .B(net368),
    .Y(_13472_));
 TIEHIx1_ASAP7_75t_R _34689__670 (.H(net670));
 TIEHIx1_ASAP7_75t_R _34688__669 (.H(net669));
 TIEHIx1_ASAP7_75t_R _34687__668 (.H(net668));
 TIEHIx1_ASAP7_75t_R _34686__667 (.H(net667));
 OA21x2_ASAP7_75t_R _18750_ (.A1(_13470_),
    .A2(_13472_),
    .B(net369),
    .Y(_13477_));
 AO32x1_ASAP7_75t_R _18751_ (.A1(_13397_),
    .A2(_13428_),
    .A3(_13451_),
    .B1(_13465_),
    .B2(_13477_),
    .Y(_13478_));
 TIEHIx1_ASAP7_75t_R _34685__666 (.H(net666));
 TIEHIx1_ASAP7_75t_R _34684__665 (.H(net665));
 TIEHIx1_ASAP7_75t_R _34683__664 (.H(net664));
 TIEHIx1_ASAP7_75t_R _34682__663 (.H(net663));
 TIEHIx1_ASAP7_75t_R _34681__662 (.H(net662));
 CKINVDCx20_ASAP7_75t_R _18757_ (.A(net365),
    .Y(_13484_));
 INVx1_ASAP7_75t_R _18758_ (.A(_00268_),
    .Y(_13485_));
 TIEHIx1_ASAP7_75t_R _34680__661 (.H(net661));
 TIEHIx1_ASAP7_75t_R _34679__660 (.H(net660));
 TIEHIx1_ASAP7_75t_R _34678__659 (.H(net659));
 NAND2x1_ASAP7_75t_R _18762_ (.A(_00266_),
    .B(net386),
    .Y(_13489_));
 TIEHIx1_ASAP7_75t_R _34677__658 (.H(net658));
 OA211x2_ASAP7_75t_R _18764_ (.A1(_13485_),
    .A2(net386),
    .B(_13489_),
    .C(net304),
    .Y(_13491_));
 NAND2x1_ASAP7_75t_R _18765_ (.A(_00265_),
    .B(net386),
    .Y(_13492_));
 TIEHIx1_ASAP7_75t_R _34676__657 (.H(net657));
 OA211x2_ASAP7_75t_R _18767_ (.A1(_13159_),
    .A2(net386),
    .B(_13492_),
    .C(net404),
    .Y(_13494_));
 OR3x1_ASAP7_75t_R _18768_ (.A(_13484_),
    .B(_13491_),
    .C(_13494_),
    .Y(_13495_));
 INVx1_ASAP7_75t_R _18769_ (.A(_00274_),
    .Y(_13496_));
 TIEHIx1_ASAP7_75t_R _34675__656 (.H(net656));
 TIEHIx1_ASAP7_75t_R _34674__655 (.H(net655));
 TIEHIx1_ASAP7_75t_R _34673__654 (.H(net654));
 NAND2x1_ASAP7_75t_R _18773_ (.A(_00273_),
    .B(net404),
    .Y(_13500_));
 OA211x2_ASAP7_75t_R _18774_ (.A1(_13496_),
    .A2(net404),
    .B(net382),
    .C(_13500_),
    .Y(_13501_));
 NAND2x1_ASAP7_75t_R _18775_ (.A(_00275_),
    .B(net404),
    .Y(_13502_));
 OA211x2_ASAP7_75t_R _18776_ (.A1(_13202_),
    .A2(net404),
    .B(net303),
    .C(_13502_),
    .Y(_13503_));
 OR3x1_ASAP7_75t_R _18777_ (.A(net368),
    .B(_13501_),
    .C(_13503_),
    .Y(_13504_));
 AND3x1_ASAP7_75t_R _18778_ (.A(_13397_),
    .B(_13495_),
    .C(_13504_),
    .Y(_13505_));
 INVx1_ASAP7_75t_R _18779_ (.A(_00264_),
    .Y(_13506_));
 NAND2x1_ASAP7_75t_R _18780_ (.A(_00262_),
    .B(net386),
    .Y(_13507_));
 OA211x2_ASAP7_75t_R _18781_ (.A1(_13506_),
    .A2(net386),
    .B(_13507_),
    .C(net305),
    .Y(_13508_));
 TIEHIx1_ASAP7_75t_R _34672__653 (.H(net653));
 TIEHIx1_ASAP7_75t_R _34671__652 (.H(net652));
 NAND2x1_ASAP7_75t_R _18784_ (.A(_00261_),
    .B(net386),
    .Y(_13511_));
 OA211x2_ASAP7_75t_R _18785_ (.A1(_13154_),
    .A2(net386),
    .B(_13511_),
    .C(net404),
    .Y(_13512_));
 OR3x1_ASAP7_75t_R _18786_ (.A(_13484_),
    .B(_13508_),
    .C(_13512_),
    .Y(_13513_));
 TIEHIx1_ASAP7_75t_R _34670__651 (.H(net651));
 NAND2x1_ASAP7_75t_R _18788_ (.A(_00269_),
    .B(net404),
    .Y(_13515_));
 OA211x2_ASAP7_75t_R _18789_ (.A1(_13198_),
    .A2(net404),
    .B(net382),
    .C(_13515_),
    .Y(_13516_));
 INVx1_ASAP7_75t_R _18790_ (.A(_00272_),
    .Y(_13517_));
 NAND2x1_ASAP7_75t_R _18791_ (.A(_00271_),
    .B(net404),
    .Y(_13518_));
 OA211x2_ASAP7_75t_R _18792_ (.A1(_13517_),
    .A2(net404),
    .B(net303),
    .C(_13518_),
    .Y(_13519_));
 OR3x1_ASAP7_75t_R _18793_ (.A(net368),
    .B(_13516_),
    .C(_13519_),
    .Y(_13520_));
 AND3x1_ASAP7_75t_R _18794_ (.A(net369),
    .B(_13513_),
    .C(_13520_),
    .Y(_13521_));
 OR3x1_ASAP7_75t_R _18795_ (.A(net363),
    .B(_13505_),
    .C(_13521_),
    .Y(_13522_));
 OA21x2_ASAP7_75t_R _18796_ (.A1(_13392_),
    .A2(_13478_),
    .B(_13522_),
    .Y(_13523_));
 TIEHIx1_ASAP7_75t_R _34638__650 (.H(net650));
 TIEHIx1_ASAP7_75t_R _34637__649 (.H(net649));
 TIEHIx1_ASAP7_75t_R _34636__648 (.H(net648));
 AND3x4_ASAP7_75t_R _18800_ (.A(_00285_),
    .B(_01357_),
    .C(_01727_),
    .Y(_13527_));
 AND2x6_ASAP7_75t_R _18801_ (.A(_00284_),
    .B(_13527_),
    .Y(_13528_));
 TIEHIx1_ASAP7_75t_R _34635__647 (.H(net647));
 CKINVDCx20_ASAP7_75t_R _18803_ (.A(_00285_),
    .Y(_13530_));
 TIEHIx1_ASAP7_75t_R _34634__646 (.H(net646));
 TIEHIx1_ASAP7_75t_R _34633__645 (.H(net645));
 NAND2x2_ASAP7_75t_R _18806_ (.A(_01357_),
    .B(_01727_),
    .Y(_13533_));
 TIEHIx1_ASAP7_75t_R _34632__644 (.H(net644));
 AO221x1_ASAP7_75t_R _18808_ (.A1(_13530_),
    .A2(_00291_),
    .B1(_01451_),
    .B2(_13533_),
    .C(net295),
    .Y(_13535_));
 AOI21x1_ASAP7_75t_R _18809_ (.A1(_13217_),
    .A2(_13528_),
    .B(_13535_),
    .Y(_13536_));
 OA21x2_ASAP7_75t_R _18810_ (.A1(_00284_),
    .A2(_13523_),
    .B(_13536_),
    .Y(_13537_));
 AOI21x1_ASAP7_75t_R _18811_ (.A1(net294),
    .A2(_13389_),
    .B(_13537_),
    .Y(_17537_));
 INVx1_ASAP7_75t_R _18812_ (.A(_17537_),
    .Y(_16497_));
 INVx1_ASAP7_75t_R _18813_ (.A(_01720_),
    .Y(\cs_registers_i.pc_id_i[1] ));
 INVx1_ASAP7_75t_R _18814_ (.A(_01640_),
    .Y(_13538_));
 TIEHIx1_ASAP7_75t_R _34631__643 (.H(net643));
 OR2x2_ASAP7_75t_R _18816_ (.A(_00163_),
    .B(_00165_),
    .Y(_13540_));
 NAND2x1_ASAP7_75t_R _18817_ (.A(_00278_),
    .B(_00175_),
    .Y(_13541_));
 OR5x2_ASAP7_75t_R _18818_ (.A(_00168_),
    .B(_13273_),
    .C(_01746_),
    .D(_13540_),
    .E(_13541_),
    .Y(_13542_));
 OR3x1_ASAP7_75t_R _18819_ (.A(_00278_),
    .B(_00163_),
    .C(_00175_),
    .Y(_13543_));
 OR4x1_ASAP7_75t_R _18820_ (.A(_13256_),
    .B(_13273_),
    .C(_01746_),
    .D(_13543_),
    .Y(_13544_));
 OR4x1_ASAP7_75t_R _18821_ (.A(_13255_),
    .B(_00163_),
    .C(_01746_),
    .D(_13245_),
    .Y(_13545_));
 OR4x1_ASAP7_75t_R _18822_ (.A(_00278_),
    .B(_00163_),
    .C(_00175_),
    .D(_01746_),
    .Y(_13546_));
 OR3x4_ASAP7_75t_R _18823_ (.A(_00172_),
    .B(_13245_),
    .C(_13546_),
    .Y(_13547_));
 TIEHIx1_ASAP7_75t_R _34630__642 (.H(net642));
 AND4x2_ASAP7_75t_R _18825_ (.A(_13542_),
    .B(_13544_),
    .C(_13545_),
    .D(_13547_),
    .Y(_13549_));
 NAND3x2_ASAP7_75t_R _18826_ (.B(_00281_),
    .C(_00282_),
    .Y(_13550_),
    .A(_00279_));
 AND5x2_ASAP7_75t_R _18827_ (.A(_13325_),
    .B(_13273_),
    .C(_13230_),
    .D(_13234_),
    .E(_13252_),
    .Y(_13551_));
 AO221x2_ASAP7_75t_R _18828_ (.A1(_13228_),
    .A2(_13280_),
    .B1(_13550_),
    .B2(_13267_),
    .C(_13551_),
    .Y(_13552_));
 OA21x2_ASAP7_75t_R _18829_ (.A1(_13549_),
    .A2(_13552_),
    .B(_13223_),
    .Y(_13553_));
 TIEHIx1_ASAP7_75t_R _34629__641 (.H(net641));
 NAND2x1_ASAP7_75t_R _18831_ (.A(_13542_),
    .B(_13547_),
    .Y(_13555_));
 OR4x1_ASAP7_75t_R _18832_ (.A(_00278_),
    .B(_00168_),
    .C(_13273_),
    .D(_00175_),
    .Y(_13556_));
 OR3x1_ASAP7_75t_R _18833_ (.A(_13256_),
    .B(_00172_),
    .C(_13541_),
    .Y(_13557_));
 OR3x1_ASAP7_75t_R _18834_ (.A(_00163_),
    .B(_00165_),
    .C(_01746_),
    .Y(_13558_));
 AO21x1_ASAP7_75t_R _18835_ (.A1(_13556_),
    .A2(_13557_),
    .B(_13558_),
    .Y(_13559_));
 AO211x2_ASAP7_75t_R _18836_ (.A1(_13323_),
    .A2(_13267_),
    .B(_13285_),
    .C(_13286_),
    .Y(_13560_));
 AO221x2_ASAP7_75t_R _18837_ (.A1(_13325_),
    .A2(_13555_),
    .B1(_13549_),
    .B2(_13559_),
    .C(_13560_),
    .Y(_13561_));
 TIEHIx1_ASAP7_75t_R _34628__640 (.H(net640));
 NOR2x2_ASAP7_75t_R _18839_ (.A(_13553_),
    .B(_13561_),
    .Y(_13563_));
 TIEHIx1_ASAP7_75t_R _34627__639 (.H(net639));
 TIEHIx1_ASAP7_75t_R _34626__638 (.H(net638));
 TIEHIx1_ASAP7_75t_R _34625__637 (.H(net637));
 AND5x2_ASAP7_75t_R _18843_ (.A(_13273_),
    .B(_13230_),
    .C(_13234_),
    .D(_13252_),
    .E(_13550_),
    .Y(_13567_));
 TIEHIx1_ASAP7_75t_R _34624__636 (.H(net636));
 AND3x1_ASAP7_75t_R _18845_ (.A(_13433_),
    .B(_13567_),
    .C(_13561_),
    .Y(_13569_));
 NOR2x1_ASAP7_75t_R _18846_ (.A(_01720_),
    .B(_13561_),
    .Y(_13570_));
 TIEHIx1_ASAP7_75t_R _34623__635 (.H(net635));
 OA21x2_ASAP7_75t_R _18848_ (.A1(_13569_),
    .A2(_13570_),
    .B(_13553_),
    .Y(_13572_));
 AO221x2_ASAP7_75t_R _18849_ (.A1(_13538_),
    .A2(_13270_),
    .B1(_13523_),
    .B2(_13563_),
    .C(_13572_),
    .Y(_13573_));
 TIEHIx1_ASAP7_75t_R _34622__634 (.H(net634));
 INVx3_ASAP7_75t_R _18851_ (.A(_13573_),
    .Y(_18114_));
 AND2x6_ASAP7_75t_R _18852_ (.A(_01357_),
    .B(_01727_),
    .Y(_13574_));
 TIEHIx1_ASAP7_75t_R _34621__633 (.H(net633));
 AND3x4_ASAP7_75t_R _18854_ (.A(_13238_),
    .B(_13313_),
    .C(_13316_),
    .Y(_13576_));
 TIEHIx1_ASAP7_75t_R _34620__632 (.H(net632));
 TIEHIx1_ASAP7_75t_R _34619__631 (.H(net631));
 TIEHIx1_ASAP7_75t_R _34618__630 (.H(net630));
 TIEHIx1_ASAP7_75t_R _34617__629 (.H(net629));
 TIEHIx1_ASAP7_75t_R _34616__628 (.H(net628));
 OA21x2_ASAP7_75t_R _18860_ (.A1(_00291_),
    .A2(_13574_),
    .B(_13576_),
    .Y(_13582_));
 AOI21x1_ASAP7_75t_R _18861_ (.A1(net294),
    .A2(_18114_),
    .B(_13582_),
    .Y(_17538_));
 INVx1_ASAP7_75t_R _18862_ (.A(_17538_),
    .Y(_16498_));
 AND2x6_ASAP7_75t_R _18863_ (.A(_13223_),
    .B(_13248_),
    .Y(_13583_));
 NAND2x2_ASAP7_75t_R _18864_ (.A(net322),
    .B(net321),
    .Y(_13584_));
 TIEHIx1_ASAP7_75t_R _34615__627 (.H(net627));
 NAND2x2_ASAP7_75t_R _18866_ (.A(net356),
    .B(net312),
    .Y(_13586_));
 AND2x2_ASAP7_75t_R _18867_ (.A(net327),
    .B(_01709_),
    .Y(_13587_));
 AO21x1_ASAP7_75t_R _18868_ (.A1(net312),
    .A2(_00294_),
    .B(_13587_),
    .Y(_13588_));
 OAI22x1_ASAP7_75t_R _18869_ (.A1(_00293_),
    .A2(_13586_),
    .B1(_13588_),
    .B2(net354),
    .Y(_13589_));
 INVx1_ASAP7_75t_R _18870_ (.A(_00306_),
    .Y(_13590_));
 NAND2x1_ASAP7_75t_R _18871_ (.A(net329),
    .B(_00304_),
    .Y(_13591_));
 OA211x2_ASAP7_75t_R _18872_ (.A1(net329),
    .A2(_13590_),
    .B(_13591_),
    .C(net310),
    .Y(_13592_));
 INVx1_ASAP7_75t_R _18873_ (.A(_00305_),
    .Y(_13593_));
 NAND2x1_ASAP7_75t_R _18874_ (.A(net329),
    .B(_00303_),
    .Y(_13594_));
 OA211x2_ASAP7_75t_R _18875_ (.A1(net329),
    .A2(_13593_),
    .B(_13594_),
    .C(net354),
    .Y(_13595_));
 OR4x1_ASAP7_75t_R _18876_ (.A(net322),
    .B(net321),
    .C(_13592_),
    .D(_13595_),
    .Y(_13596_));
 OA211x2_ASAP7_75t_R _18877_ (.A1(_13584_),
    .A2(_13589_),
    .B(_13596_),
    .C(net316),
    .Y(_13597_));
 CKINVDCx20_ASAP7_75t_R _18878_ (.A(net320),
    .Y(_13598_));
 AND2x2_ASAP7_75t_R _18879_ (.A(net327),
    .B(_00295_),
    .Y(_13599_));
 AO21x1_ASAP7_75t_R _18880_ (.A1(net312),
    .A2(_00297_),
    .B(_13599_),
    .Y(_13600_));
 AND2x2_ASAP7_75t_R _18881_ (.A(net327),
    .B(_00296_),
    .Y(_13601_));
 AO21x1_ASAP7_75t_R _18882_ (.A1(net312),
    .A2(_00298_),
    .B(_13601_),
    .Y(_13602_));
 AOI22x1_ASAP7_75t_R _18883_ (.A1(_13133_),
    .A2(_13600_),
    .B1(_13602_),
    .B2(_13124_),
    .Y(_13603_));
 INVx1_ASAP7_75t_R _18884_ (.A(_00301_),
    .Y(_13604_));
 TIEHIx1_ASAP7_75t_R _34614__626 (.H(net626));
 NAND2x1_ASAP7_75t_R _18886_ (.A(net327),
    .B(_00299_),
    .Y(_13606_));
 OA211x2_ASAP7_75t_R _18887_ (.A1(net327),
    .A2(_13604_),
    .B(_13606_),
    .C(net354),
    .Y(_13607_));
 TIEHIx1_ASAP7_75t_R _34613__625 (.H(net625));
 INVx1_ASAP7_75t_R _18889_ (.A(_00302_),
    .Y(_13609_));
 NAND2x1_ASAP7_75t_R _18890_ (.A(net327),
    .B(_00300_),
    .Y(_13610_));
 OA211x2_ASAP7_75t_R _18891_ (.A1(net327),
    .A2(_13609_),
    .B(_13610_),
    .C(net310),
    .Y(_13611_));
 OR4x1_ASAP7_75t_R _18892_ (.A(_13132_),
    .B(net321),
    .C(_13607_),
    .D(_13611_),
    .Y(_13612_));
 OA21x2_ASAP7_75t_R _18893_ (.A1(_13598_),
    .A2(_13603_),
    .B(_13612_),
    .Y(_13613_));
 AND2x6_ASAP7_75t_R _18894_ (.A(net321),
    .B(_13174_),
    .Y(_13614_));
 INVx1_ASAP7_75t_R _18895_ (.A(_00310_),
    .Y(_13615_));
 NAND2x1_ASAP7_75t_R _18896_ (.A(net328),
    .B(_00308_),
    .Y(_13616_));
 OA211x2_ASAP7_75t_R _18897_ (.A1(net328),
    .A2(_13615_),
    .B(_13616_),
    .C(net322),
    .Y(_13617_));
 INVx1_ASAP7_75t_R _18898_ (.A(_00314_),
    .Y(_13618_));
 NAND2x1_ASAP7_75t_R _18899_ (.A(net328),
    .B(_00312_),
    .Y(_13619_));
 OA211x2_ASAP7_75t_R _18900_ (.A1(net328),
    .A2(_13618_),
    .B(_13619_),
    .C(_13132_),
    .Y(_13620_));
 OR3x1_ASAP7_75t_R _18901_ (.A(net354),
    .B(_13617_),
    .C(_13620_),
    .Y(_13621_));
 AND2x2_ASAP7_75t_R _18902_ (.A(net329),
    .B(_00307_),
    .Y(_13622_));
 AO21x1_ASAP7_75t_R _18903_ (.A1(net312),
    .A2(_00309_),
    .B(_13622_),
    .Y(_13623_));
 AND2x2_ASAP7_75t_R _18904_ (.A(net329),
    .B(_00311_),
    .Y(_13624_));
 AO21x1_ASAP7_75t_R _18905_ (.A1(net312),
    .A2(_00313_),
    .B(_13624_),
    .Y(_13625_));
 AOI22x1_ASAP7_75t_R _18906_ (.A1(_13184_),
    .A2(_13623_),
    .B1(_13625_),
    .B2(_13133_),
    .Y(_13626_));
 INVx1_ASAP7_75t_R _18907_ (.A(_00322_),
    .Y(_13627_));
 NAND2x1_ASAP7_75t_R _18908_ (.A(net328),
    .B(_00320_),
    .Y(_13628_));
 OA211x2_ASAP7_75t_R _18909_ (.A1(net328),
    .A2(_13627_),
    .B(_13628_),
    .C(_13132_),
    .Y(_13629_));
 INVx1_ASAP7_75t_R _18910_ (.A(_00318_),
    .Y(_13630_));
 NAND2x1_ASAP7_75t_R _18911_ (.A(net328),
    .B(_00316_),
    .Y(_13631_));
 OA211x2_ASAP7_75t_R _18912_ (.A1(net328),
    .A2(_13630_),
    .B(_13631_),
    .C(net322),
    .Y(_13632_));
 OR3x1_ASAP7_75t_R _18913_ (.A(net354),
    .B(_13629_),
    .C(_13632_),
    .Y(_13633_));
 AND2x2_ASAP7_75t_R _18914_ (.A(net329),
    .B(_00315_),
    .Y(_13634_));
 AO21x1_ASAP7_75t_R _18915_ (.A1(net312),
    .A2(_00317_),
    .B(_13634_),
    .Y(_13635_));
 AND2x2_ASAP7_75t_R _18916_ (.A(net328),
    .B(_00319_),
    .Y(_13636_));
 AO21x1_ASAP7_75t_R _18917_ (.A1(net312),
    .A2(_00321_),
    .B(_13636_),
    .Y(_13637_));
 AOI22x1_ASAP7_75t_R _18918_ (.A1(_13184_),
    .A2(_13635_),
    .B1(_13637_),
    .B2(_13133_),
    .Y(_13638_));
 AO33x2_ASAP7_75t_R _18919_ (.A1(_13614_),
    .A2(_13621_),
    .A3(_13626_),
    .B1(_13633_),
    .B2(_13638_),
    .B3(_13215_),
    .Y(_13639_));
 AO21x2_ASAP7_75t_R _18920_ (.A1(_13597_),
    .A2(_13613_),
    .B(_13639_),
    .Y(_13640_));
 TIEHIx1_ASAP7_75t_R _34612__624 (.H(net624));
 TIEHIx1_ASAP7_75t_R _34611__623 (.H(net623));
 TIEHIx1_ASAP7_75t_R _34610__622 (.H(net622));
 NOR2x1_ASAP7_75t_R _18924_ (.A(_18336_),
    .B(_01608_),
    .Y(_13644_));
 XOR2x2_ASAP7_75t_R _18925_ (.A(_00277_),
    .B(_01608_),
    .Y(_13645_));
 TIEHIx1_ASAP7_75t_R _34609__621 (.H(net621));
 AO221x1_ASAP7_75t_R _18927_ (.A1(_00277_),
    .A2(_13644_),
    .B1(_13645_),
    .B2(_01609_),
    .C(net360),
    .Y(_13647_));
 AO221x1_ASAP7_75t_R _18928_ (.A1(_13279_),
    .A2(_13290_),
    .B1(_13280_),
    .B2(_13249_),
    .C(_13647_),
    .Y(_13648_));
 NOR2x1_ASAP7_75t_R _18929_ (.A(_13298_),
    .B(_13648_),
    .Y(_13649_));
 AO211x2_ASAP7_75t_R _18930_ (.A1(_13228_),
    .A2(_13235_),
    .B(_13239_),
    .C(_13247_),
    .Y(_13650_));
 TIEHIx1_ASAP7_75t_R _34608__620 (.H(net620));
 INVx2_ASAP7_75t_R _18932_ (.A(_00323_),
    .Y(_13652_));
 AND2x4_ASAP7_75t_R _18933_ (.A(_13223_),
    .B(_13291_),
    .Y(_13653_));
 OA211x2_ASAP7_75t_R _18934_ (.A1(_13296_),
    .A2(_13297_),
    .B(_13258_),
    .C(_13254_),
    .Y(_13654_));
 AND3x1_ASAP7_75t_R _18935_ (.A(_13652_),
    .B(_13653_),
    .C(_13654_),
    .Y(_13655_));
 AOI221x1_ASAP7_75t_R _18936_ (.A1(_13583_),
    .A2(_13640_),
    .B1(_13649_),
    .B2(_13650_),
    .C(_13655_),
    .Y(_13656_));
 TIEHIx1_ASAP7_75t_R _34607__619 (.H(net619));
 CKINVDCx20_ASAP7_75t_R _18938_ (.A(net289),
    .Y(_13658_));
 TIEHIx1_ASAP7_75t_R _34606__618 (.H(net618));
 TIEHIx1_ASAP7_75t_R _34605__617 (.H(net617));
 TIEHIx1_ASAP7_75t_R _34604__616 (.H(net616));
 TIEHIx1_ASAP7_75t_R _34603__615 (.H(net615));
 TIEHIx1_ASAP7_75t_R _34602__614 (.H(net614));
 TIEHIx1_ASAP7_75t_R _34601__613 (.H(net613));
 TIEHIx1_ASAP7_75t_R _34600__612 (.H(net612));
 TIEHIx1_ASAP7_75t_R _34599__611 (.H(net611));
 TIEHIx1_ASAP7_75t_R _34598__610 (.H(net610));
 TIEHIx1_ASAP7_75t_R _34597__609 (.H(net609));
 TIEHIx1_ASAP7_75t_R _34596__608 (.H(net608));
 TIEHIx1_ASAP7_75t_R _34595__607 (.H(net607));
 TIEHIx1_ASAP7_75t_R _34594__606 (.H(net606));
 TIEHIx1_ASAP7_75t_R _34593__605 (.H(net605));
 TIEHIx1_ASAP7_75t_R _34592__604 (.H(net604));
 TIEHIx1_ASAP7_75t_R _34591__603 (.H(net603));
 TIEHIx1_ASAP7_75t_R _34590__602 (.H(net602));
 TIEHIx1_ASAP7_75t_R _34589__601 (.H(net601));
 AND2x2_ASAP7_75t_R _18957_ (.A(net381),
    .B(_01709_),
    .Y(_13675_));
 AO21x1_ASAP7_75t_R _18958_ (.A1(net303),
    .A2(_00294_),
    .B(_13675_),
    .Y(_13676_));
 TIEHIx1_ASAP7_75t_R _34588__600 (.H(net600));
 OAI22x1_ASAP7_75t_R _18960_ (.A1(_00293_),
    .A2(_13471_),
    .B1(_13676_),
    .B2(net406),
    .Y(_13678_));
 TIEHIx1_ASAP7_75t_R _34587__599 (.H(net599));
 TIEHIx1_ASAP7_75t_R _34586__598 (.H(net598));
 TIEHIx1_ASAP7_75t_R _34585__597 (.H(net597));
 NAND2x1_ASAP7_75t_R _18964_ (.A(net380),
    .B(_00308_),
    .Y(_13682_));
 TIEHIx1_ASAP7_75t_R _34584__596 (.H(net596));
 OA211x2_ASAP7_75t_R _18966_ (.A1(net380),
    .A2(_13615_),
    .B(_13682_),
    .C(net305),
    .Y(_13684_));
 TIEHIx1_ASAP7_75t_R _34583__595 (.H(net595));
 TIEHIx1_ASAP7_75t_R _34582__594 (.H(net594));
 TIEHIx1_ASAP7_75t_R _34581__593 (.H(net593));
 INVx1_ASAP7_75t_R _18970_ (.A(_00309_),
    .Y(_13688_));
 TIEHIx1_ASAP7_75t_R _34580__592 (.H(net592));
 NAND2x1_ASAP7_75t_R _18972_ (.A(net381),
    .B(_00307_),
    .Y(_13690_));
 TIEHIx1_ASAP7_75t_R _34579__591 (.H(net591));
 OA211x2_ASAP7_75t_R _18974_ (.A1(net381),
    .A2(_13688_),
    .B(_13690_),
    .C(net406),
    .Y(_13692_));
 OR3x1_ASAP7_75t_R _18975_ (.A(net363),
    .B(_13684_),
    .C(_13692_),
    .Y(_13693_));
 OA21x2_ASAP7_75t_R _18976_ (.A1(_13392_),
    .A2(_13678_),
    .B(_13693_),
    .Y(_13694_));
 TIEHIx1_ASAP7_75t_R _34578__590 (.H(net590));
 TIEHIx1_ASAP7_75t_R _34577__589 (.H(net589));
 TIEHIx1_ASAP7_75t_R _34576__588 (.H(net588));
 TIEHIx1_ASAP7_75t_R _34575__587 (.H(net587));
 INVx1_ASAP7_75t_R _18981_ (.A(_00298_),
    .Y(_13699_));
 TIEHIx1_ASAP7_75t_R _34574__586 (.H(net586));
 NAND2x1_ASAP7_75t_R _18983_ (.A(net381),
    .B(_00296_),
    .Y(_13701_));
 OA211x2_ASAP7_75t_R _18984_ (.A1(net381),
    .A2(_13699_),
    .B(_13701_),
    .C(net304),
    .Y(_13702_));
 TIEHIx1_ASAP7_75t_R _34573__585 (.H(net585));
 INVx1_ASAP7_75t_R _18986_ (.A(_00297_),
    .Y(_13704_));
 NAND2x1_ASAP7_75t_R _18987_ (.A(net381),
    .B(_00295_),
    .Y(_13705_));
 TIEHIx1_ASAP7_75t_R _34572__584 (.H(net584));
 OA211x2_ASAP7_75t_R _18989_ (.A1(net381),
    .A2(_13704_),
    .B(_13705_),
    .C(net406),
    .Y(_13707_));
 OR3x1_ASAP7_75t_R _18990_ (.A(_13392_),
    .B(_13702_),
    .C(_13707_),
    .Y(_13708_));
 NAND2x1_ASAP7_75t_R _18991_ (.A(net380),
    .B(_00312_),
    .Y(_13709_));
 OA211x2_ASAP7_75t_R _18992_ (.A1(net380),
    .A2(_13618_),
    .B(_13709_),
    .C(net305),
    .Y(_13710_));
 INVx1_ASAP7_75t_R _18993_ (.A(_00313_),
    .Y(_13711_));
 NAND2x1_ASAP7_75t_R _18994_ (.A(net381),
    .B(_00311_),
    .Y(_13712_));
 OA211x2_ASAP7_75t_R _18995_ (.A1(net381),
    .A2(_13711_),
    .B(_13712_),
    .C(net406),
    .Y(_13713_));
 OR3x1_ASAP7_75t_R _18996_ (.A(net363),
    .B(_13710_),
    .C(_13713_),
    .Y(_13714_));
 AND3x1_ASAP7_75t_R _18997_ (.A(_13397_),
    .B(_13708_),
    .C(_13714_),
    .Y(_13715_));
 AO21x1_ASAP7_75t_R _18998_ (.A1(net375),
    .A2(_13694_),
    .B(_13715_),
    .Y(_13716_));
 TIEHIx1_ASAP7_75t_R _34571__583 (.H(net583));
 TIEHIx1_ASAP7_75t_R _34570__582 (.H(net582));
 TIEHIx1_ASAP7_75t_R _34569__581 (.H(net581));
 NAND2x1_ASAP7_75t_R _19002_ (.A(net381),
    .B(_00300_),
    .Y(_13720_));
 TIEHIx1_ASAP7_75t_R _34568__580 (.H(net580));
 OA211x2_ASAP7_75t_R _19004_ (.A1(net381),
    .A2(_13609_),
    .B(_13720_),
    .C(net304),
    .Y(_13722_));
 TIEHIx1_ASAP7_75t_R _34567__579 (.H(net579));
 TIEHIx1_ASAP7_75t_R _34566__578 (.H(net578));
 NAND2x1_ASAP7_75t_R _19007_ (.A(net381),
    .B(_00299_),
    .Y(_13725_));
 OA211x2_ASAP7_75t_R _19008_ (.A1(net381),
    .A2(_13604_),
    .B(_13725_),
    .C(net406),
    .Y(_13726_));
 OR3x1_ASAP7_75t_R _19009_ (.A(_13397_),
    .B(_13722_),
    .C(_13726_),
    .Y(_13727_));
 TIEHIx1_ASAP7_75t_R _34565__577 (.H(net577));
 TIEHIx1_ASAP7_75t_R _34564__576 (.H(net576));
 NAND2x1_ASAP7_75t_R _19012_ (.A(net381),
    .B(_00304_),
    .Y(_13730_));
 OA211x2_ASAP7_75t_R _19013_ (.A1(net381),
    .A2(_13590_),
    .B(_13730_),
    .C(net304),
    .Y(_13731_));
 TIEHIx1_ASAP7_75t_R _34563__575 (.H(net575));
 TIEHIx1_ASAP7_75t_R _34562__574 (.H(net574));
 NAND2x1_ASAP7_75t_R _19016_ (.A(net381),
    .B(_00303_),
    .Y(_13734_));
 OA211x2_ASAP7_75t_R _19017_ (.A1(net381),
    .A2(_13593_),
    .B(_13734_),
    .C(net406),
    .Y(_13735_));
 OR3x1_ASAP7_75t_R _19018_ (.A(net375),
    .B(_13731_),
    .C(_13735_),
    .Y(_13736_));
 AND3x1_ASAP7_75t_R _19019_ (.A(net363),
    .B(_13727_),
    .C(_13736_),
    .Y(_13737_));
 TIEHIx1_ASAP7_75t_R _34561__573 (.H(net573));
 NAND2x1_ASAP7_75t_R _19021_ (.A(net380),
    .B(_00316_),
    .Y(_13739_));
 OA211x2_ASAP7_75t_R _19022_ (.A1(net380),
    .A2(_13630_),
    .B(_13739_),
    .C(net305),
    .Y(_13740_));
 INVx1_ASAP7_75t_R _19023_ (.A(_00317_),
    .Y(_13741_));
 NAND2x1_ASAP7_75t_R _19024_ (.A(net380),
    .B(_00315_),
    .Y(_13742_));
 TIEHIx1_ASAP7_75t_R _34560__572 (.H(net572));
 OA211x2_ASAP7_75t_R _19026_ (.A1(net380),
    .A2(_13741_),
    .B(_13742_),
    .C(net406),
    .Y(_13744_));
 OR3x1_ASAP7_75t_R _19027_ (.A(_13397_),
    .B(_13740_),
    .C(_13744_),
    .Y(_13745_));
 NAND2x1_ASAP7_75t_R _19028_ (.A(net380),
    .B(_00320_),
    .Y(_13746_));
 TIEHIx1_ASAP7_75t_R _34559__571 (.H(net571));
 OA211x2_ASAP7_75t_R _19030_ (.A1(net380),
    .A2(_13627_),
    .B(_13746_),
    .C(net305),
    .Y(_13748_));
 TIEHIx1_ASAP7_75t_R _34558__570 (.H(net570));
 TIEHIx1_ASAP7_75t_R _34557__569 (.H(net569));
 INVx1_ASAP7_75t_R _19033_ (.A(_00321_),
    .Y(_13751_));
 TIEHIx1_ASAP7_75t_R _34556__568 (.H(net568));
 NAND2x1_ASAP7_75t_R _19035_ (.A(net380),
    .B(_00319_),
    .Y(_13753_));
 OA211x2_ASAP7_75t_R _19036_ (.A1(net380),
    .A2(_13751_),
    .B(_13753_),
    .C(net406),
    .Y(_13754_));
 OR3x1_ASAP7_75t_R _19037_ (.A(net375),
    .B(_13748_),
    .C(_13754_),
    .Y(_13755_));
 AND3x1_ASAP7_75t_R _19038_ (.A(_13392_),
    .B(_13745_),
    .C(_13755_),
    .Y(_13756_));
 OR3x1_ASAP7_75t_R _19039_ (.A(net368),
    .B(_13737_),
    .C(_13756_),
    .Y(_13757_));
 OA21x2_ASAP7_75t_R _19040_ (.A1(_13484_),
    .A2(_13716_),
    .B(_13757_),
    .Y(_13758_));
 TIEHIx1_ASAP7_75t_R _34555__567 (.H(net567));
 TIEHIx1_ASAP7_75t_R _34554__566 (.H(net566));
 TIEHIx1_ASAP7_75t_R _34553__565 (.H(net565));
 AOI22x1_ASAP7_75t_R _19044_ (.A1(_13530_),
    .A2(_00324_),
    .B1(_01452_),
    .B2(_13533_),
    .Y(_13762_));
 NAND2x2_ASAP7_75t_R _19045_ (.A(_00284_),
    .B(_13527_),
    .Y(_13763_));
 TIEHIx1_ASAP7_75t_R _34552__564 (.H(net564));
 OA211x2_ASAP7_75t_R _19047_ (.A1(_00284_),
    .A2(_13758_),
    .B(_13762_),
    .C(_13763_),
    .Y(_13765_));
 AO21x1_ASAP7_75t_R _19048_ (.A1(_13528_),
    .A2(_13640_),
    .B(_13765_),
    .Y(_13766_));
 TIEHIx1_ASAP7_75t_R _34551__563 (.H(net563));
 TIEHIx1_ASAP7_75t_R _34550__562 (.H(net562));
 TIEHIx1_ASAP7_75t_R _34549__561 (.H(net561));
 XNOR2x1_ASAP7_75t_R _19052_ (.B(net288),
    .Y(_13770_),
    .A(_13387_));
 AND2x2_ASAP7_75t_R _19053_ (.A(net294),
    .B(_13770_),
    .Y(_13771_));
 AO21x1_ASAP7_75t_R _19054_ (.A1(_13576_),
    .A2(_13766_),
    .B(_13771_),
    .Y(_16500_));
 AND4x2_ASAP7_75t_R _19055_ (.A(_13273_),
    .B(_13230_),
    .C(_13234_),
    .D(_13252_),
    .Y(_13772_));
 AND2x2_ASAP7_75t_R _19056_ (.A(net305),
    .B(_13772_),
    .Y(_13773_));
 TIEHIx1_ASAP7_75t_R _34548__560 (.H(net560));
 TIEHIx1_ASAP7_75t_R _34547__559 (.H(net559));
 NOR2x1_ASAP7_75t_R _19059_ (.A(_01641_),
    .B(_13223_),
    .Y(_13776_));
 AO221x2_ASAP7_75t_R _19060_ (.A1(_13563_),
    .A2(_13758_),
    .B1(_13773_),
    .B2(_13553_),
    .C(_13776_),
    .Y(_13777_));
 TIEHIx1_ASAP7_75t_R _34546__558 (.H(net558));
 INVx2_ASAP7_75t_R _19062_ (.A(_13777_),
    .Y(_18108_));
 TIEHIx1_ASAP7_75t_R _34545__557 (.H(net557));
 TIEHIx1_ASAP7_75t_R _34544__556 (.H(net556));
 OA21x2_ASAP7_75t_R _19065_ (.A1(_00324_),
    .A2(_13574_),
    .B(_13576_),
    .Y(_13780_));
 AO21x1_ASAP7_75t_R _19066_ (.A1(net294),
    .A2(_18108_),
    .B(_13780_),
    .Y(_16501_));
 AND2x6_ASAP7_75t_R _19067_ (.A(net294),
    .B(_13387_),
    .Y(_13781_));
 TIEHIx1_ASAP7_75t_R _34543__555 (.H(net555));
 OR2x6_ASAP7_75t_R _19069_ (.A(_13553_),
    .B(_13561_),
    .Y(_13782_));
 TIEHIx1_ASAP7_75t_R _34542__554 (.H(net554));
 TIEHIx1_ASAP7_75t_R _34541__553 (.H(net553));
 TIEHIx1_ASAP7_75t_R _34540__552 (.H(net552));
 TIEHIx1_ASAP7_75t_R _34539__551 (.H(net551));
 TIEHIx1_ASAP7_75t_R _34538__550 (.H(net550));
 TIEHIx1_ASAP7_75t_R _34537__549 (.H(net549));
 INVx1_ASAP7_75t_R _19076_ (.A(_00335_),
    .Y(_13789_));
 TIEHIx1_ASAP7_75t_R _34536__548 (.H(net548));
 NOR2x1_ASAP7_75t_R _19078_ (.A(net380),
    .B(_00337_),
    .Y(_13791_));
 AO21x1_ASAP7_75t_R _19079_ (.A1(net380),
    .A2(_13789_),
    .B(_13791_),
    .Y(_13792_));
 TIEHIx1_ASAP7_75t_R _34535__547 (.H(net547));
 INVx1_ASAP7_75t_R _19081_ (.A(_00338_),
    .Y(_13794_));
 TIEHIx1_ASAP7_75t_R _34534__546 (.H(net546));
 NAND2x1_ASAP7_75t_R _19083_ (.A(net380),
    .B(_00336_),
    .Y(_13796_));
 TIEHIx1_ASAP7_75t_R _34533__545 (.H(net545));
 TIEHIx1_ASAP7_75t_R _34532__544 (.H(net544));
 OA211x2_ASAP7_75t_R _19086_ (.A1(net380),
    .A2(_13794_),
    .B(_13796_),
    .C(net305),
    .Y(_13799_));
 AO21x1_ASAP7_75t_R _19087_ (.A1(net406),
    .A2(_13792_),
    .B(_13799_),
    .Y(_13800_));
 TIEHIx1_ASAP7_75t_R _34531__543 (.H(net543));
 INVx1_ASAP7_75t_R _19089_ (.A(_00334_),
    .Y(_13802_));
 NAND2x1_ASAP7_75t_R _19090_ (.A(net381),
    .B(_00332_),
    .Y(_13803_));
 TIEHIx1_ASAP7_75t_R _34530__542 (.H(net542));
 OA211x2_ASAP7_75t_R _19092_ (.A1(net381),
    .A2(_13802_),
    .B(_13803_),
    .C(net305),
    .Y(_13805_));
 TIEHIx1_ASAP7_75t_R _34529__541 (.H(net541));
 TIEHIx1_ASAP7_75t_R _34528__540 (.H(net540));
 INVx1_ASAP7_75t_R _19095_ (.A(_00333_),
    .Y(_13808_));
 NAND2x1_ASAP7_75t_R _19096_ (.A(net381),
    .B(_00331_),
    .Y(_13809_));
 TIEHIx1_ASAP7_75t_R _34527__539 (.H(net539));
 OA211x2_ASAP7_75t_R _19098_ (.A1(net381),
    .A2(_13808_),
    .B(_13809_),
    .C(net404),
    .Y(_13811_));
 OR3x1_ASAP7_75t_R _19099_ (.A(_13397_),
    .B(_13805_),
    .C(_13811_),
    .Y(_13812_));
 OA21x2_ASAP7_75t_R _19100_ (.A1(net369),
    .A2(_13800_),
    .B(_13812_),
    .Y(_13813_));
 NAND2x2_ASAP7_75t_R _19101_ (.A(_13397_),
    .B(net366),
    .Y(_13814_));
 TIEHIx1_ASAP7_75t_R _34526__538 (.H(net538));
 TIEHIx1_ASAP7_75t_R _34525__537 (.H(net537));
 TIEHIx1_ASAP7_75t_R _34524__536 (.H(net536));
 INVx1_ASAP7_75t_R _19105_ (.A(_00329_),
    .Y(_13818_));
 NAND2x1_ASAP7_75t_R _19106_ (.A(net381),
    .B(_00327_),
    .Y(_13819_));
 OA211x2_ASAP7_75t_R _19107_ (.A1(net381),
    .A2(_13818_),
    .B(_13819_),
    .C(net406),
    .Y(_13820_));
 INVx1_ASAP7_75t_R _19108_ (.A(_00330_),
    .Y(_13821_));
 NAND2x1_ASAP7_75t_R _19109_ (.A(net381),
    .B(_00328_),
    .Y(_13822_));
 TIEHIx1_ASAP7_75t_R _34523__535 (.H(net535));
 OA211x2_ASAP7_75t_R _19111_ (.A1(net381),
    .A2(_13821_),
    .B(_13822_),
    .C(net305),
    .Y(_13824_));
 INVx1_ASAP7_75t_R _19112_ (.A(_00326_),
    .Y(_13825_));
 NAND2x1_ASAP7_75t_R _19113_ (.A(net381),
    .B(_01697_),
    .Y(_13826_));
 OA211x2_ASAP7_75t_R _19114_ (.A1(net381),
    .A2(_13825_),
    .B(_13826_),
    .C(net305),
    .Y(_13827_));
 NAND2x2_ASAP7_75t_R _19115_ (.A(net370),
    .B(net366),
    .Y(_13828_));
 TIEHIx1_ASAP7_75t_R _34522__534 (.H(net534));
 TIEHIx1_ASAP7_75t_R _34521__533 (.H(net533));
 NOR2x1_ASAP7_75t_R _19118_ (.A(_00325_),
    .B(_13471_),
    .Y(_13831_));
 OA33x2_ASAP7_75t_R _19119_ (.A1(net298),
    .A2(_13820_),
    .A3(_13824_),
    .B1(_13827_),
    .B2(net301),
    .B3(_13831_),
    .Y(_13832_));
 OAI21x1_ASAP7_75t_R _19120_ (.A1(net368),
    .A2(_13813_),
    .B(_13832_),
    .Y(_13833_));
 TIEHIx1_ASAP7_75t_R _34520__532 (.H(net532));
 INVx1_ASAP7_75t_R _19122_ (.A(_00341_),
    .Y(_13835_));
 TIEHIx1_ASAP7_75t_R _34519__531 (.H(net531));
 NAND2x1_ASAP7_75t_R _19124_ (.A(net380),
    .B(_00339_),
    .Y(_13837_));
 OA211x2_ASAP7_75t_R _19125_ (.A1(net380),
    .A2(_13835_),
    .B(_13837_),
    .C(net375),
    .Y(_13838_));
 INVx1_ASAP7_75t_R _19126_ (.A(_00345_),
    .Y(_13839_));
 NAND2x1_ASAP7_75t_R _19127_ (.A(net380),
    .B(_00343_),
    .Y(_13840_));
 OA211x2_ASAP7_75t_R _19128_ (.A1(net380),
    .A2(_13839_),
    .B(_13840_),
    .C(_13397_),
    .Y(_13841_));
 OR3x1_ASAP7_75t_R _19129_ (.A(net305),
    .B(_13838_),
    .C(_13841_),
    .Y(_13842_));
 TIEHIx1_ASAP7_75t_R _34518__530 (.H(net530));
 TIEHIx1_ASAP7_75t_R _34517__529 (.H(net529));
 TIEHIx1_ASAP7_75t_R _34516__528 (.H(net528));
 TIEHIx1_ASAP7_75t_R _34515__527 (.H(net527));
 INVx1_ASAP7_75t_R _19134_ (.A(_00342_),
    .Y(_13847_));
 NAND2x1_ASAP7_75t_R _19135_ (.A(net380),
    .B(_00340_),
    .Y(_13848_));
 TIEHIx1_ASAP7_75t_R _34514__526 (.H(net526));
 TIEHIx1_ASAP7_75t_R _34513__525 (.H(net525));
 OA211x2_ASAP7_75t_R _19138_ (.A1(net380),
    .A2(_13847_),
    .B(_13848_),
    .C(net375),
    .Y(_13851_));
 INVx1_ASAP7_75t_R _19139_ (.A(_00346_),
    .Y(_13852_));
 TIEHIx1_ASAP7_75t_R _34512__524 (.H(net524));
 NAND2x1_ASAP7_75t_R _19141_ (.A(net380),
    .B(_00344_),
    .Y(_13854_));
 OA211x2_ASAP7_75t_R _19142_ (.A1(net380),
    .A2(_13852_),
    .B(_13854_),
    .C(_13397_),
    .Y(_13855_));
 OR3x1_ASAP7_75t_R _19143_ (.A(net406),
    .B(_13851_),
    .C(_13855_),
    .Y(_13856_));
 NAND2x1_ASAP7_75t_R _19144_ (.A(_13842_),
    .B(_13856_),
    .Y(_13857_));
 TIEHIx1_ASAP7_75t_R _34511__523 (.H(net523));
 TIEHIx1_ASAP7_75t_R _34510__522 (.H(net522));
 INVx1_ASAP7_75t_R _19147_ (.A(_00349_),
    .Y(_13860_));
 NAND2x1_ASAP7_75t_R _19148_ (.A(net380),
    .B(_00347_),
    .Y(_13861_));
 TIEHIx1_ASAP7_75t_R _34509__521 (.H(net521));
 OA211x2_ASAP7_75t_R _19150_ (.A1(net380),
    .A2(_13860_),
    .B(_13861_),
    .C(net375),
    .Y(_13863_));
 INVx1_ASAP7_75t_R _19151_ (.A(_00353_),
    .Y(_13864_));
 NAND2x1_ASAP7_75t_R _19152_ (.A(net380),
    .B(_00351_),
    .Y(_13865_));
 OA211x2_ASAP7_75t_R _19153_ (.A1(net380),
    .A2(_13864_),
    .B(_13865_),
    .C(_13397_),
    .Y(_13866_));
 OR3x1_ASAP7_75t_R _19154_ (.A(net305),
    .B(_13863_),
    .C(_13866_),
    .Y(_13867_));
 INVx1_ASAP7_75t_R _19155_ (.A(_00350_),
    .Y(_13868_));
 NAND2x1_ASAP7_75t_R _19156_ (.A(net380),
    .B(_00348_),
    .Y(_13869_));
 TIEHIx1_ASAP7_75t_R _34508__520 (.H(net520));
 OA211x2_ASAP7_75t_R _19158_ (.A1(net380),
    .A2(_13868_),
    .B(_13869_),
    .C(net375),
    .Y(_13871_));
 INVx1_ASAP7_75t_R _19159_ (.A(_00354_),
    .Y(_13872_));
 NAND2x1_ASAP7_75t_R _19160_ (.A(net380),
    .B(_00352_),
    .Y(_13873_));
 OA211x2_ASAP7_75t_R _19161_ (.A1(net380),
    .A2(_13872_),
    .B(_13873_),
    .C(_13397_),
    .Y(_13874_));
 OR3x1_ASAP7_75t_R _19162_ (.A(net406),
    .B(_13871_),
    .C(_13874_),
    .Y(_13875_));
 NAND3x1_ASAP7_75t_R _19163_ (.A(_13484_),
    .B(_13867_),
    .C(_13875_),
    .Y(_13876_));
 OA211x2_ASAP7_75t_R _19164_ (.A1(_13484_),
    .A2(_13857_),
    .B(_13876_),
    .C(_13392_),
    .Y(_13877_));
 AO21x2_ASAP7_75t_R _19165_ (.A1(net363),
    .A2(_13833_),
    .B(_13877_),
    .Y(_13878_));
 OAI21x1_ASAP7_75t_R _19166_ (.A1(_13549_),
    .A2(_13552_),
    .B(_13223_),
    .Y(_13879_));
 OR2x6_ASAP7_75t_R _19167_ (.A(_13879_),
    .B(_13561_),
    .Y(_13880_));
 TIEHIx1_ASAP7_75t_R _34507__519 (.H(net519));
 OA22x2_ASAP7_75t_R _19169_ (.A1(_01629_),
    .A2(_13223_),
    .B1(_13880_),
    .B2(_00199_),
    .Y(_13882_));
 OAI21x1_ASAP7_75t_R _19170_ (.A1(_13782_),
    .A2(_13878_),
    .B(_13882_),
    .Y(_18165_));
 INVx6_ASAP7_75t_R _19171_ (.A(_18165_),
    .Y(_18167_));
 INVx1_ASAP7_75t_R _19172_ (.A(_00375_),
    .Y(_13883_));
 NAND2x1_ASAP7_75t_R _19173_ (.A(net341),
    .B(_00373_),
    .Y(_13884_));
 OA211x2_ASAP7_75t_R _19174_ (.A1(net341),
    .A2(_13883_),
    .B(_13133_),
    .C(_13884_),
    .Y(_13885_));
 TIEHIx1_ASAP7_75t_R _34506__518 (.H(net518));
 INVx1_ASAP7_75t_R _19176_ (.A(_00376_),
    .Y(_13887_));
 NAND2x1_ASAP7_75t_R _19177_ (.A(net341),
    .B(_00374_),
    .Y(_13888_));
 OA211x2_ASAP7_75t_R _19178_ (.A1(net341),
    .A2(_13887_),
    .B(_13124_),
    .C(_13888_),
    .Y(_13889_));
 INVx1_ASAP7_75t_R _19179_ (.A(_00372_),
    .Y(_13890_));
 NAND2x1_ASAP7_75t_R _19180_ (.A(net341),
    .B(_00370_),
    .Y(_13891_));
 OA211x2_ASAP7_75t_R _19181_ (.A1(net341),
    .A2(_13890_),
    .B(_13164_),
    .C(_13891_),
    .Y(_13892_));
 INVx1_ASAP7_75t_R _19182_ (.A(_00371_),
    .Y(_13893_));
 NAND2x1_ASAP7_75t_R _19183_ (.A(net341),
    .B(_00369_),
    .Y(_13894_));
 OA211x2_ASAP7_75t_R _19184_ (.A1(net341),
    .A2(_13893_),
    .B(_13184_),
    .C(_13894_),
    .Y(_13895_));
 OR4x1_ASAP7_75t_R _19185_ (.A(_13885_),
    .B(_13889_),
    .C(_13892_),
    .D(_13895_),
    .Y(_13896_));
 INVx1_ASAP7_75t_R _19186_ (.A(_00363_),
    .Y(_13897_));
 NAND2x1_ASAP7_75t_R _19187_ (.A(net350),
    .B(_00361_),
    .Y(_13898_));
 OA21x2_ASAP7_75t_R _19188_ (.A1(net350),
    .A2(_13897_),
    .B(_13898_),
    .Y(_13899_));
 INVx1_ASAP7_75t_R _19189_ (.A(_00367_),
    .Y(_13900_));
 NAND2x1_ASAP7_75t_R _19190_ (.A(net350),
    .B(_00365_),
    .Y(_13901_));
 OA21x2_ASAP7_75t_R _19191_ (.A1(net350),
    .A2(_13900_),
    .B(_13901_),
    .Y(_13902_));
 INVx1_ASAP7_75t_R _19192_ (.A(_00368_),
    .Y(_13903_));
 NAND2x1_ASAP7_75t_R _19193_ (.A(net350),
    .B(_00366_),
    .Y(_13904_));
 OA211x2_ASAP7_75t_R _19194_ (.A1(net350),
    .A2(_13903_),
    .B(_13124_),
    .C(_13904_),
    .Y(_13905_));
 AO221x1_ASAP7_75t_R _19195_ (.A1(_13184_),
    .A2(_13899_),
    .B1(_13902_),
    .B2(_13133_),
    .C(_13905_),
    .Y(_13906_));
 TIEHIx1_ASAP7_75t_R _34505__517 (.H(net517));
 INVx1_ASAP7_75t_R _19197_ (.A(_00364_),
    .Y(_13908_));
 NAND2x1_ASAP7_75t_R _19198_ (.A(net350),
    .B(_00362_),
    .Y(_13909_));
 OA21x2_ASAP7_75t_R _19199_ (.A1(net350),
    .A2(_13908_),
    .B(_13909_),
    .Y(_13910_));
 AO21x1_ASAP7_75t_R _19200_ (.A1(_13164_),
    .A2(_13910_),
    .B(net320),
    .Y(_13911_));
 AND2x2_ASAP7_75t_R _19201_ (.A(net341),
    .B(_00357_),
    .Y(_13912_));
 AO21x1_ASAP7_75t_R _19202_ (.A1(net313),
    .A2(_00359_),
    .B(_13912_),
    .Y(_13913_));
 AND2x2_ASAP7_75t_R _19203_ (.A(net341),
    .B(_00358_),
    .Y(_13914_));
 AO21x1_ASAP7_75t_R _19204_ (.A1(net313),
    .A2(_00360_),
    .B(_13914_),
    .Y(_13915_));
 AOI22x1_ASAP7_75t_R _19205_ (.A1(_13133_),
    .A2(_13913_),
    .B1(_13915_),
    .B2(_13124_),
    .Y(_13916_));
 INVx1_ASAP7_75t_R _19206_ (.A(_00355_),
    .Y(_13917_));
 INVx1_ASAP7_75t_R _19207_ (.A(_01707_),
    .Y(_13918_));
 NOR2x1_ASAP7_75t_R _19208_ (.A(net341),
    .B(_00356_),
    .Y(_13919_));
 AO21x1_ASAP7_75t_R _19209_ (.A1(net341),
    .A2(_13918_),
    .B(_13919_),
    .Y(_13920_));
 TIEHIx1_ASAP7_75t_R _34504__516 (.H(net516));
 AO221x1_ASAP7_75t_R _19211_ (.A1(_13917_),
    .A2(_13190_),
    .B1(_13920_),
    .B2(net309),
    .C(_13584_),
    .Y(_13922_));
 OA221x2_ASAP7_75t_R _19212_ (.A1(_13906_),
    .A2(_13911_),
    .B1(_13916_),
    .B2(_13598_),
    .C(_13922_),
    .Y(_13923_));
 TIEHIx1_ASAP7_75t_R _34503__515 (.H(net515));
 INVx1_ASAP7_75t_R _19214_ (.A(_00381_),
    .Y(_13925_));
 NOR2x1_ASAP7_75t_R _19215_ (.A(net350),
    .B(_00383_),
    .Y(_13926_));
 AO21x1_ASAP7_75t_R _19216_ (.A1(net350),
    .A2(_13925_),
    .B(_13926_),
    .Y(_13927_));
 TIEHIx1_ASAP7_75t_R _34502__514 (.H(net514));
 INVx1_ASAP7_75t_R _19218_ (.A(_00384_),
    .Y(_13929_));
 NAND2x1_ASAP7_75t_R _19219_ (.A(net350),
    .B(_00382_),
    .Y(_13930_));
 OA211x2_ASAP7_75t_R _19220_ (.A1(net350),
    .A2(_13929_),
    .B(_13124_),
    .C(_13930_),
    .Y(_13931_));
 AO21x1_ASAP7_75t_R _19221_ (.A1(_13133_),
    .A2(_13927_),
    .B(_13931_),
    .Y(_13932_));
 AND2x6_ASAP7_75t_R _19222_ (.A(net349),
    .B(net323),
    .Y(_13933_));
 NAND2x1_ASAP7_75t_R _19223_ (.A(net309),
    .B(_00378_),
    .Y(_13934_));
 TIEHIx1_ASAP7_75t_R _34501__513 (.H(net513));
 NAND2x1_ASAP7_75t_R _19225_ (.A(net359),
    .B(_00377_),
    .Y(_13936_));
 INVx1_ASAP7_75t_R _19226_ (.A(_00379_),
    .Y(_13937_));
 NOR2x1_ASAP7_75t_R _19227_ (.A(net359),
    .B(_00380_),
    .Y(_13938_));
 AO21x1_ASAP7_75t_R _19228_ (.A1(net359),
    .A2(_13937_),
    .B(_13938_),
    .Y(_13939_));
 AND2x4_ASAP7_75t_R _19229_ (.A(net313),
    .B(net323),
    .Y(_13940_));
 AO32x1_ASAP7_75t_R _19230_ (.A1(_13933_),
    .A2(_13934_),
    .A3(_13936_),
    .B1(_13939_),
    .B2(_13940_),
    .Y(_13941_));
 OA21x2_ASAP7_75t_R _19231_ (.A1(_13932_),
    .A2(_13941_),
    .B(_13215_),
    .Y(_13942_));
 AO221x2_ASAP7_75t_R _19232_ (.A1(_13614_),
    .A2(_13896_),
    .B1(_13923_),
    .B2(net314),
    .C(_13942_),
    .Y(_13943_));
 TIEHIx1_ASAP7_75t_R _34500__512 (.H(net512));
 AND3x1_ASAP7_75t_R _19234_ (.A(_00385_),
    .B(_13281_),
    .C(_13654_),
    .Y(_13945_));
 TIEHIx1_ASAP7_75t_R _34499__511 (.H(net511));
 TIEHIx1_ASAP7_75t_R _34498__510 (.H(net510));
 AND2x2_ASAP7_75t_R _19237_ (.A(_13223_),
    .B(_13650_),
    .Y(_13948_));
 OAI21x1_ASAP7_75t_R _19238_ (.A1(_01744_),
    .A2(_13298_),
    .B(_13948_),
    .Y(_13949_));
 INVx2_ASAP7_75t_R _19239_ (.A(_00187_),
    .Y(_13950_));
 NAND2x2_ASAP7_75t_R _19240_ (.A(_13271_),
    .B(_13274_),
    .Y(_13951_));
 AND3x2_ASAP7_75t_R _19241_ (.A(_13223_),
    .B(_13951_),
    .C(_13291_),
    .Y(_13952_));
 AND3x1_ASAP7_75t_R _19242_ (.A(_13950_),
    .B(_13298_),
    .C(_13952_),
    .Y(_13953_));
 OA33x2_ASAP7_75t_R _19243_ (.A1(_13270_),
    .A2(_13650_),
    .A3(_13943_),
    .B1(_13945_),
    .B2(_13949_),
    .B3(_13953_),
    .Y(_13954_));
 CKINVDCx14_ASAP7_75t_R _19244_ (.A(_13954_),
    .Y(_13955_));
 TIEHIx1_ASAP7_75t_R _34497__509 (.H(net509));
 TIEHIx1_ASAP7_75t_R _34496__508 (.H(net508));
 TIEHIx1_ASAP7_75t_R _34495__507 (.H(net507));
 TIEHIx1_ASAP7_75t_R _34494__506 (.H(net506));
 TIEHIx1_ASAP7_75t_R _34493__505 (.H(net505));
 TIEHIx1_ASAP7_75t_R _34492__504 (.H(net504));
 AND2x2_ASAP7_75t_R _19251_ (.A(net349),
    .B(_00408_),
    .Y(_13961_));
 AO21x1_ASAP7_75t_R _19252_ (.A1(net312),
    .A2(_00410_),
    .B(_13961_),
    .Y(_13962_));
 TIEHIx1_ASAP7_75t_R _34491__503 (.H(net503));
 AND2x2_ASAP7_75t_R _19254_ (.A(net349),
    .B(_00412_),
    .Y(_13964_));
 AO21x1_ASAP7_75t_R _19255_ (.A1(net312),
    .A2(_00414_),
    .B(_13964_),
    .Y(_13965_));
 TIEHIx1_ASAP7_75t_R _34490__502 (.H(net502));
 AOI22x1_ASAP7_75t_R _19257_ (.A1(_13184_),
    .A2(_13962_),
    .B1(_13965_),
    .B2(_13133_),
    .Y(_13967_));
 INVx1_ASAP7_75t_R _19258_ (.A(_00415_),
    .Y(_13968_));
 TIEHIx1_ASAP7_75t_R _34489__501 (.H(net501));
 NAND2x1_ASAP7_75t_R _19260_ (.A(net349),
    .B(_00413_),
    .Y(_13970_));
 OA211x2_ASAP7_75t_R _19261_ (.A1(net349),
    .A2(_13968_),
    .B(_13970_),
    .C(_13132_),
    .Y(_13971_));
 INVx1_ASAP7_75t_R _19262_ (.A(_00411_),
    .Y(_13972_));
 NAND2x1_ASAP7_75t_R _19263_ (.A(net349),
    .B(_00409_),
    .Y(_13973_));
 OA211x2_ASAP7_75t_R _19264_ (.A1(net349),
    .A2(_13972_),
    .B(_13973_),
    .C(net323),
    .Y(_13974_));
 OR3x1_ASAP7_75t_R _19265_ (.A(net354),
    .B(_13971_),
    .C(_13974_),
    .Y(_13975_));
 OR2x4_ASAP7_75t_R _19266_ (.A(net317),
    .B(net314),
    .Y(_13976_));
 AO21x1_ASAP7_75t_R _19267_ (.A1(_13967_),
    .A2(_13975_),
    .B(_13976_),
    .Y(_13977_));
 AND2x2_ASAP7_75t_R _19268_ (.A(net347),
    .B(_00388_),
    .Y(_13978_));
 AO21x1_ASAP7_75t_R _19269_ (.A1(net312),
    .A2(_00390_),
    .B(_13978_),
    .Y(_13979_));
 AND2x2_ASAP7_75t_R _19270_ (.A(net347),
    .B(_00389_),
    .Y(_13980_));
 AO21x1_ASAP7_75t_R _19271_ (.A1(net312),
    .A2(_00391_),
    .B(_13980_),
    .Y(_13981_));
 AOI22x1_ASAP7_75t_R _19272_ (.A1(_13133_),
    .A2(_13979_),
    .B1(_13981_),
    .B2(_13124_),
    .Y(_13982_));
 INVx1_ASAP7_75t_R _19273_ (.A(_00386_),
    .Y(_13983_));
 TIEHIx1_ASAP7_75t_R _34488__500 (.H(net500));
 AND2x2_ASAP7_75t_R _19275_ (.A(net347),
    .B(_01706_),
    .Y(_13985_));
 AOI21x1_ASAP7_75t_R _19276_ (.A1(net312),
    .A2(_00387_),
    .B(_13985_),
    .Y(_13986_));
 TIEHIx1_ASAP7_75t_R _34487__499 (.H(net499));
 TIEHIx1_ASAP7_75t_R _34486__498 (.H(net498));
 AO221x1_ASAP7_75t_R _19279_ (.A1(_13983_),
    .A2(_13190_),
    .B1(_13986_),
    .B2(net311),
    .C(_13132_),
    .Y(_13989_));
 AO21x1_ASAP7_75t_R _19280_ (.A1(_13982_),
    .A2(_13989_),
    .B(_13122_),
    .Y(_13990_));
 TIEHIx1_ASAP7_75t_R _34485__497 (.H(net497));
 TIEHIx1_ASAP7_75t_R _34484__496 (.H(net496));
 INVx1_ASAP7_75t_R _19283_ (.A(_00403_),
    .Y(_13993_));
 NAND2x1_ASAP7_75t_R _19284_ (.A(net348),
    .B(_00401_),
    .Y(_13994_));
 OA211x2_ASAP7_75t_R _19285_ (.A1(net348),
    .A2(_13993_),
    .B(_13164_),
    .C(_13994_),
    .Y(_13995_));
 INVx1_ASAP7_75t_R _19286_ (.A(_00402_),
    .Y(_13996_));
 NAND2x1_ASAP7_75t_R _19287_ (.A(net348),
    .B(_00400_),
    .Y(_13997_));
 OA211x2_ASAP7_75t_R _19288_ (.A1(net348),
    .A2(_13996_),
    .B(_13184_),
    .C(_13997_),
    .Y(_13998_));
 NAND2x1_ASAP7_75t_R _19289_ (.A(net343),
    .B(_00405_),
    .Y(_13999_));
 NAND2x1_ASAP7_75t_R _19290_ (.A(net312),
    .B(_00407_),
    .Y(_14000_));
 NAND2x1_ASAP7_75t_R _19291_ (.A(net343),
    .B(_00404_),
    .Y(_14001_));
 NAND2x1_ASAP7_75t_R _19292_ (.A(net312),
    .B(_00406_),
    .Y(_14002_));
 AO33x2_ASAP7_75t_R _19293_ (.A1(_13124_),
    .A2(_13999_),
    .A3(_14000_),
    .B1(_14001_),
    .B2(_14002_),
    .B3(_13133_),
    .Y(_14003_));
 OR4x1_ASAP7_75t_R _19294_ (.A(_13175_),
    .B(_13995_),
    .C(_13998_),
    .D(_14003_),
    .Y(_14004_));
 TIEHIx1_ASAP7_75t_R _34483__495 (.H(net495));
 INVx1_ASAP7_75t_R _19296_ (.A(_00399_),
    .Y(_14006_));
 NAND2x1_ASAP7_75t_R _19297_ (.A(net349),
    .B(_00397_),
    .Y(_14007_));
 OA211x2_ASAP7_75t_R _19298_ (.A1(net349),
    .A2(_14006_),
    .B(_13124_),
    .C(_14007_),
    .Y(_14008_));
 NAND2x1_ASAP7_75t_R _19299_ (.A(net348),
    .B(_00392_),
    .Y(_14009_));
 NAND2x1_ASAP7_75t_R _19300_ (.A(net312),
    .B(_00394_),
    .Y(_14010_));
 NAND2x1_ASAP7_75t_R _19301_ (.A(net348),
    .B(_00393_),
    .Y(_14011_));
 NAND2x1_ASAP7_75t_R _19302_ (.A(net312),
    .B(_00395_),
    .Y(_14012_));
 AO33x2_ASAP7_75t_R _19303_ (.A1(_13184_),
    .A2(_14009_),
    .A3(_14010_),
    .B1(_14011_),
    .B2(_14012_),
    .B3(_13164_),
    .Y(_14013_));
 TIEHIx1_ASAP7_75t_R _34482__494 (.H(net494));
 INVx1_ASAP7_75t_R _19305_ (.A(_00398_),
    .Y(_14015_));
 NAND2x1_ASAP7_75t_R _19306_ (.A(net349),
    .B(_00396_),
    .Y(_14016_));
 OA211x2_ASAP7_75t_R _19307_ (.A1(net349),
    .A2(_14015_),
    .B(_13133_),
    .C(_14016_),
    .Y(_14017_));
 OR5x1_ASAP7_75t_R _19308_ (.A(net317),
    .B(_13174_),
    .C(_14008_),
    .D(_14013_),
    .E(_14017_),
    .Y(_14018_));
 AND4x2_ASAP7_75t_R _19309_ (.A(_13977_),
    .B(_13990_),
    .C(_14004_),
    .D(_14018_),
    .Y(_14019_));
 TIEHIx1_ASAP7_75t_R _34481__493 (.H(net493));
 INVx2_ASAP7_75t_R _19311_ (.A(_00191_),
    .Y(_14021_));
 AND3x1_ASAP7_75t_R _19312_ (.A(_14021_),
    .B(_13298_),
    .C(_13952_),
    .Y(_14022_));
 NAND2x2_ASAP7_75t_R _19313_ (.A(_13598_),
    .B(_13650_),
    .Y(_14023_));
 NOR2x2_ASAP7_75t_R _19314_ (.A(_13298_),
    .B(_14023_),
    .Y(_14024_));
 AOI211x1_ASAP7_75t_R _19315_ (.A1(_13583_),
    .A2(_14019_),
    .B(_14022_),
    .C(_14024_),
    .Y(_14025_));
 CKINVDCx9p33_ASAP7_75t_R _19316_ (.A(_14025_),
    .Y(_14026_));
 TIEHIx1_ASAP7_75t_R _34480__492 (.H(net492));
 TIEHIx1_ASAP7_75t_R _34479__491 (.H(net491));
 INVx3_ASAP7_75t_R _19319_ (.A(_00194_),
    .Y(_14027_));
 AND2x2_ASAP7_75t_R _19320_ (.A(_13298_),
    .B(_13952_),
    .Y(_14028_));
 INVx1_ASAP7_75t_R _19321_ (.A(_00440_),
    .Y(_14029_));
 NAND2x1_ASAP7_75t_R _19322_ (.A(net310),
    .B(_00441_),
    .Y(_14030_));
 OA211x2_ASAP7_75t_R _19323_ (.A1(net310),
    .A2(_14029_),
    .B(_13940_),
    .C(_14030_),
    .Y(_14031_));
 INVx1_ASAP7_75t_R _19324_ (.A(_00439_),
    .Y(_14032_));
 NAND2x1_ASAP7_75t_R _19325_ (.A(net354),
    .B(_00438_),
    .Y(_14033_));
 OA211x2_ASAP7_75t_R _19326_ (.A1(net354),
    .A2(_14032_),
    .B(_13933_),
    .C(_14033_),
    .Y(_14034_));
 INVx1_ASAP7_75t_R _19327_ (.A(_00444_),
    .Y(_14035_));
 NAND2x1_ASAP7_75t_R _19328_ (.A(net329),
    .B(_00442_),
    .Y(_14036_));
 OA211x2_ASAP7_75t_R _19329_ (.A1(net329),
    .A2(_14035_),
    .B(_13133_),
    .C(_14036_),
    .Y(_14037_));
 INVx1_ASAP7_75t_R _19330_ (.A(_00445_),
    .Y(_14038_));
 NAND2x1_ASAP7_75t_R _19331_ (.A(net329),
    .B(_00443_),
    .Y(_14039_));
 OA211x2_ASAP7_75t_R _19332_ (.A1(net329),
    .A2(_14038_),
    .B(_13124_),
    .C(_14039_),
    .Y(_14040_));
 OR4x1_ASAP7_75t_R _19333_ (.A(_14031_),
    .B(_14034_),
    .C(_14037_),
    .D(_14040_),
    .Y(_14041_));
 INVx1_ASAP7_75t_R _19334_ (.A(_00428_),
    .Y(_14042_));
 NAND2x1_ASAP7_75t_R _19335_ (.A(net326),
    .B(_00426_),
    .Y(_14043_));
 OA211x2_ASAP7_75t_R _19336_ (.A1(net326),
    .A2(_14042_),
    .B(_13133_),
    .C(_14043_),
    .Y(_14044_));
 TIEHIx1_ASAP7_75t_R _34478__490 (.H(net490));
 AND2x2_ASAP7_75t_R _19338_ (.A(net326),
    .B(_00422_),
    .Y(_14046_));
 AO21x1_ASAP7_75t_R _19339_ (.A1(net313),
    .A2(_00424_),
    .B(_14046_),
    .Y(_14047_));
 OR2x2_ASAP7_75t_R _19340_ (.A(net326),
    .B(_00425_),
    .Y(_14048_));
 OA211x2_ASAP7_75t_R _19341_ (.A1(net313),
    .A2(_00423_),
    .B(_14048_),
    .C(net310),
    .Y(_14049_));
 AOI211x1_ASAP7_75t_R _19342_ (.A1(_00246_),
    .A2(_14047_),
    .B(_14049_),
    .C(_13132_),
    .Y(_14050_));
 INVx1_ASAP7_75t_R _19343_ (.A(_00429_),
    .Y(_14051_));
 NAND2x1_ASAP7_75t_R _19344_ (.A(net326),
    .B(_00427_),
    .Y(_14052_));
 OA211x2_ASAP7_75t_R _19345_ (.A1(net326),
    .A2(_14051_),
    .B(_13124_),
    .C(_14052_),
    .Y(_14053_));
 OR4x1_ASAP7_75t_R _19346_ (.A(net321),
    .B(_14044_),
    .C(_14050_),
    .D(_14053_),
    .Y(_14054_));
 AND2x2_ASAP7_75t_R _19347_ (.A(net326),
    .B(_00418_),
    .Y(_14055_));
 AO21x1_ASAP7_75t_R _19348_ (.A1(net313),
    .A2(_00420_),
    .B(_14055_),
    .Y(_14056_));
 AND2x2_ASAP7_75t_R _19349_ (.A(net326),
    .B(_00419_),
    .Y(_14057_));
 AO21x1_ASAP7_75t_R _19350_ (.A1(net313),
    .A2(_00421_),
    .B(_14057_),
    .Y(_14058_));
 AOI22x1_ASAP7_75t_R _19351_ (.A1(_13133_),
    .A2(_14056_),
    .B1(_14058_),
    .B2(_13124_),
    .Y(_14059_));
 INVx1_ASAP7_75t_R _19352_ (.A(_00416_),
    .Y(_14060_));
 INVx1_ASAP7_75t_R _19353_ (.A(_00417_),
    .Y(_14061_));
 NAND2x1_ASAP7_75t_R _19354_ (.A(net329),
    .B(_01705_),
    .Y(_14062_));
 OA21x2_ASAP7_75t_R _19355_ (.A1(net329),
    .A2(_14061_),
    .B(_14062_),
    .Y(_14063_));
 AO221x1_ASAP7_75t_R _19356_ (.A1(_14060_),
    .A2(_13190_),
    .B1(_14063_),
    .B2(net310),
    .C(_13584_),
    .Y(_14064_));
 OA211x2_ASAP7_75t_R _19357_ (.A1(_13598_),
    .A2(_14059_),
    .B(_14064_),
    .C(_00244_),
    .Y(_14065_));
 INVx1_ASAP7_75t_R _19358_ (.A(_00436_),
    .Y(_14066_));
 NAND2x1_ASAP7_75t_R _19359_ (.A(net329),
    .B(_00434_),
    .Y(_14067_));
 OA211x2_ASAP7_75t_R _19360_ (.A1(net329),
    .A2(_14066_),
    .B(_13133_),
    .C(_14067_),
    .Y(_14068_));
 INVx1_ASAP7_75t_R _19361_ (.A(_00437_),
    .Y(_14069_));
 NAND2x1_ASAP7_75t_R _19362_ (.A(net329),
    .B(_00435_),
    .Y(_14070_));
 OA211x2_ASAP7_75t_R _19363_ (.A1(net329),
    .A2(_14069_),
    .B(_13124_),
    .C(_14070_),
    .Y(_14071_));
 INVx1_ASAP7_75t_R _19364_ (.A(_00433_),
    .Y(_14072_));
 NAND2x1_ASAP7_75t_R _19365_ (.A(net328),
    .B(_00431_),
    .Y(_14073_));
 OA21x2_ASAP7_75t_R _19366_ (.A1(net328),
    .A2(_14072_),
    .B(_14073_),
    .Y(_14074_));
 INVx1_ASAP7_75t_R _19367_ (.A(_00432_),
    .Y(_14075_));
 NAND2x1_ASAP7_75t_R _19368_ (.A(net328),
    .B(_00430_),
    .Y(_14076_));
 OA211x2_ASAP7_75t_R _19369_ (.A1(net328),
    .A2(_14075_),
    .B(_13184_),
    .C(_14076_),
    .Y(_14077_));
 AO21x1_ASAP7_75t_R _19370_ (.A1(_13164_),
    .A2(_14074_),
    .B(_14077_),
    .Y(_14078_));
 OR3x1_ASAP7_75t_R _19371_ (.A(_14068_),
    .B(_14071_),
    .C(_14078_),
    .Y(_14079_));
 AO222x2_ASAP7_75t_R _19372_ (.A1(_13215_),
    .A2(_14041_),
    .B1(_14054_),
    .B2(_14065_),
    .C1(_14079_),
    .C2(_13614_),
    .Y(_14080_));
 TIEHIx1_ASAP7_75t_R _34477__489 (.H(net489));
 AND3x2_ASAP7_75t_R _19374_ (.A(_13174_),
    .B(_13299_),
    .C(_13269_),
    .Y(_14082_));
 AOI221x1_ASAP7_75t_R _19375_ (.A1(_14027_),
    .A2(_14028_),
    .B1(_14080_),
    .B2(_13583_),
    .C(_14082_),
    .Y(_14083_));
 CKINVDCx9p33_ASAP7_75t_R _19376_ (.A(_14083_),
    .Y(_14084_));
 TIEHIx1_ASAP7_75t_R _34476__488 (.H(net488));
 TIEHIx1_ASAP7_75t_R _34475__487 (.H(net487));
 INVx1_ASAP7_75t_R _19379_ (.A(_02054_),
    .Y(\cs_registers_i.mhpmcounter[2][44] ));
 INVx1_ASAP7_75t_R _19380_ (.A(_02160_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[44] ));
 INVx1_ASAP7_75t_R _19381_ (.A(_00463_),
    .Y(_14085_));
 NAND2x1_ASAP7_75t_R _19382_ (.A(net341),
    .B(_00461_),
    .Y(_14086_));
 OA211x2_ASAP7_75t_R _19383_ (.A1(net341),
    .A2(_14085_),
    .B(_13164_),
    .C(_14086_),
    .Y(_14087_));
 INVx1_ASAP7_75t_R _19384_ (.A(_00462_),
    .Y(_14088_));
 NAND2x1_ASAP7_75t_R _19385_ (.A(net341),
    .B(_00460_),
    .Y(_14089_));
 OA211x2_ASAP7_75t_R _19386_ (.A1(net341),
    .A2(_14088_),
    .B(_13184_),
    .C(_14089_),
    .Y(_14090_));
 INVx1_ASAP7_75t_R _19387_ (.A(_00466_),
    .Y(_14091_));
 NAND2x1_ASAP7_75t_R _19388_ (.A(net341),
    .B(_00464_),
    .Y(_14092_));
 OA211x2_ASAP7_75t_R _19389_ (.A1(net341),
    .A2(_14091_),
    .B(_13133_),
    .C(_14092_),
    .Y(_14093_));
 INVx1_ASAP7_75t_R _19390_ (.A(_00467_),
    .Y(_14094_));
 NAND2x1_ASAP7_75t_R _19391_ (.A(net341),
    .B(_00465_),
    .Y(_14095_));
 OA211x2_ASAP7_75t_R _19392_ (.A1(net341),
    .A2(_14094_),
    .B(_13124_),
    .C(_14095_),
    .Y(_14096_));
 OR4x1_ASAP7_75t_R _19393_ (.A(_14087_),
    .B(_14090_),
    .C(_14093_),
    .D(_14096_),
    .Y(_14097_));
 INVx1_ASAP7_75t_R _19394_ (.A(_00458_),
    .Y(_14098_));
 NAND2x1_ASAP7_75t_R _19395_ (.A(net347),
    .B(_00456_),
    .Y(_14099_));
 OA21x2_ASAP7_75t_R _19396_ (.A1(net347),
    .A2(_14098_),
    .B(_14099_),
    .Y(_14100_));
 INVx1_ASAP7_75t_R _19397_ (.A(_00454_),
    .Y(_14101_));
 NAND2x1_ASAP7_75t_R _19398_ (.A(net347),
    .B(_00452_),
    .Y(_14102_));
 OA211x2_ASAP7_75t_R _19399_ (.A1(net347),
    .A2(_14101_),
    .B(_13184_),
    .C(_14102_),
    .Y(_14103_));
 AO21x1_ASAP7_75t_R _19400_ (.A1(_13133_),
    .A2(_14100_),
    .B(_14103_),
    .Y(_14104_));
 INVx1_ASAP7_75t_R _19401_ (.A(_00459_),
    .Y(_14105_));
 NAND2x1_ASAP7_75t_R _19402_ (.A(net347),
    .B(_00457_),
    .Y(_14106_));
 OA211x2_ASAP7_75t_R _19403_ (.A1(net347),
    .A2(_14105_),
    .B(_13124_),
    .C(_14106_),
    .Y(_14107_));
 INVx1_ASAP7_75t_R _19404_ (.A(_00455_),
    .Y(_14108_));
 NAND2x1_ASAP7_75t_R _19405_ (.A(net347),
    .B(_00453_),
    .Y(_14109_));
 OA211x2_ASAP7_75t_R _19406_ (.A1(net347),
    .A2(_14108_),
    .B(_13164_),
    .C(_14109_),
    .Y(_14110_));
 OR4x1_ASAP7_75t_R _19407_ (.A(net319),
    .B(_14104_),
    .C(_14107_),
    .D(_14110_),
    .Y(_14111_));
 AND2x2_ASAP7_75t_R _19408_ (.A(net347),
    .B(_00448_),
    .Y(_14112_));
 AO21x1_ASAP7_75t_R _19409_ (.A1(net312),
    .A2(_00450_),
    .B(_14112_),
    .Y(_14113_));
 AND2x2_ASAP7_75t_R _19410_ (.A(net347),
    .B(_00449_),
    .Y(_14114_));
 AO21x1_ASAP7_75t_R _19411_ (.A1(net312),
    .A2(_00451_),
    .B(_14114_),
    .Y(_14115_));
 AOI22x1_ASAP7_75t_R _19412_ (.A1(_13133_),
    .A2(_14113_),
    .B1(_14115_),
    .B2(_13124_),
    .Y(_14116_));
 INVx1_ASAP7_75t_R _19413_ (.A(_00446_),
    .Y(_14117_));
 INVx1_ASAP7_75t_R _19414_ (.A(_00447_),
    .Y(_14118_));
 NAND2x1_ASAP7_75t_R _19415_ (.A(net347),
    .B(_01704_),
    .Y(_14119_));
 OA21x2_ASAP7_75t_R _19416_ (.A1(net347),
    .A2(_14118_),
    .B(_14119_),
    .Y(_14120_));
 AO221x1_ASAP7_75t_R _19417_ (.A1(_14117_),
    .A2(_13190_),
    .B1(_14120_),
    .B2(net310),
    .C(_13584_),
    .Y(_14121_));
 OA211x2_ASAP7_75t_R _19418_ (.A1(_13598_),
    .A2(_14116_),
    .B(_14121_),
    .C(net314),
    .Y(_14122_));
 NAND2x1_ASAP7_75t_R _19419_ (.A(net341),
    .B(_00468_),
    .Y(_14123_));
 NAND2x1_ASAP7_75t_R _19420_ (.A(net313),
    .B(_00470_),
    .Y(_14124_));
 NAND2x1_ASAP7_75t_R _19421_ (.A(net341),
    .B(_00469_),
    .Y(_14125_));
 NAND2x1_ASAP7_75t_R _19422_ (.A(net313),
    .B(_00471_),
    .Y(_14126_));
 AO33x2_ASAP7_75t_R _19423_ (.A1(_13184_),
    .A2(_14123_),
    .A3(_14124_),
    .B1(_14125_),
    .B2(_14126_),
    .B3(_13164_),
    .Y(_14127_));
 INVx1_ASAP7_75t_R _19424_ (.A(_00475_),
    .Y(_14128_));
 NAND2x1_ASAP7_75t_R _19425_ (.A(net341),
    .B(_00473_),
    .Y(_14129_));
 OA211x2_ASAP7_75t_R _19426_ (.A1(net341),
    .A2(_14128_),
    .B(_14129_),
    .C(net309),
    .Y(_14130_));
 INVx1_ASAP7_75t_R _19427_ (.A(_00474_),
    .Y(_14131_));
 NAND2x1_ASAP7_75t_R _19428_ (.A(net341),
    .B(_00472_),
    .Y(_14132_));
 OA211x2_ASAP7_75t_R _19429_ (.A1(net341),
    .A2(_14131_),
    .B(_14132_),
    .C(net359),
    .Y(_14133_));
 AND2x2_ASAP7_75t_R _19430_ (.A(_13132_),
    .B(_13215_),
    .Y(_14134_));
 OA21x2_ASAP7_75t_R _19431_ (.A1(_14130_),
    .A2(_14133_),
    .B(_14134_),
    .Y(_14135_));
 AO21x1_ASAP7_75t_R _19432_ (.A1(_13215_),
    .A2(_14127_),
    .B(_14135_),
    .Y(_14136_));
 AO221x2_ASAP7_75t_R _19433_ (.A1(_13614_),
    .A2(_14097_),
    .B1(_14111_),
    .B2(_14122_),
    .C(_14136_),
    .Y(_14137_));
 OA211x2_ASAP7_75t_R _19434_ (.A1(_13269_),
    .A2(_13653_),
    .B(_13299_),
    .C(_13951_),
    .Y(_14138_));
 AO32x2_ASAP7_75t_R _19435_ (.A1(_13223_),
    .A2(_13248_),
    .A3(_14137_),
    .B1(_14138_),
    .B2(_13306_),
    .Y(_14139_));
 TIEHIx1_ASAP7_75t_R _34474__486 (.H(net486));
 INVx8_ASAP7_75t_R _19437_ (.A(_14139_),
    .Y(_14140_));
 TIEHIx1_ASAP7_75t_R _34473__485 (.H(net485));
 INVx5_ASAP7_75t_R _19439_ (.A(_00283_),
    .Y(_14141_));
 OA211x2_ASAP7_75t_R _19440_ (.A1(_13269_),
    .A2(_13653_),
    .B(_14141_),
    .C(_13951_),
    .Y(_14142_));
 INVx1_ASAP7_75t_R _19441_ (.A(_00497_),
    .Y(_14143_));
 NAND2x1_ASAP7_75t_R _19442_ (.A(net353),
    .B(_00495_),
    .Y(_14144_));
 OA211x2_ASAP7_75t_R _19443_ (.A1(net353),
    .A2(_14143_),
    .B(_14144_),
    .C(net309),
    .Y(_14145_));
 INVx1_ASAP7_75t_R _19444_ (.A(_00496_),
    .Y(_14146_));
 NAND2x1_ASAP7_75t_R _19445_ (.A(net353),
    .B(_00494_),
    .Y(_14147_));
 OA211x2_ASAP7_75t_R _19446_ (.A1(net353),
    .A2(_14146_),
    .B(_14147_),
    .C(_00246_),
    .Y(_14148_));
 OR3x1_ASAP7_75t_R _19447_ (.A(net322),
    .B(_14145_),
    .C(_14148_),
    .Y(_14149_));
 AND2x2_ASAP7_75t_R _19448_ (.A(net352),
    .B(_00490_),
    .Y(_14150_));
 AO21x1_ASAP7_75t_R _19449_ (.A1(net313),
    .A2(_00492_),
    .B(_14150_),
    .Y(_14151_));
 AND2x2_ASAP7_75t_R _19450_ (.A(net352),
    .B(_00491_),
    .Y(_14152_));
 AO21x1_ASAP7_75t_R _19451_ (.A1(net313),
    .A2(_00493_),
    .B(_14152_),
    .Y(_14153_));
 AOI221x1_ASAP7_75t_R _19452_ (.A1(_13184_),
    .A2(_14151_),
    .B1(_14153_),
    .B2(_13164_),
    .C(_13175_),
    .Y(_14154_));
 AND2x4_ASAP7_75t_R _19453_ (.A(net361),
    .B(net352),
    .Y(_14155_));
 OR3x2_ASAP7_75t_R _19454_ (.A(net322),
    .B(_00245_),
    .C(net316),
    .Y(_14156_));
 AOI221x1_ASAP7_75t_R _19455_ (.A1(_00504_),
    .A2(_13190_),
    .B1(_14155_),
    .B2(_00502_),
    .C(_14156_),
    .Y(_14157_));
 AND2x2_ASAP7_75t_R _19456_ (.A(net353),
    .B(_00503_),
    .Y(_14158_));
 AO21x1_ASAP7_75t_R _19457_ (.A1(net313),
    .A2(_00505_),
    .B(_14158_),
    .Y(_14159_));
 NAND2x1_ASAP7_75t_R _19458_ (.A(net309),
    .B(_14159_),
    .Y(_14160_));
 INVx1_ASAP7_75t_R _19459_ (.A(_00501_),
    .Y(_14161_));
 NAND2x1_ASAP7_75t_R _19460_ (.A(net353),
    .B(_00499_),
    .Y(_14162_));
 OA211x2_ASAP7_75t_R _19461_ (.A1(net353),
    .A2(_14161_),
    .B(_14162_),
    .C(net309),
    .Y(_14163_));
 INVx1_ASAP7_75t_R _19462_ (.A(_00500_),
    .Y(_14164_));
 NAND2x1_ASAP7_75t_R _19463_ (.A(net353),
    .B(_00498_),
    .Y(_14165_));
 OA211x2_ASAP7_75t_R _19464_ (.A1(net353),
    .A2(_14164_),
    .B(_14165_),
    .C(net361),
    .Y(_14166_));
 OA211x2_ASAP7_75t_R _19465_ (.A1(_14163_),
    .A2(_14166_),
    .B(net322),
    .C(_13215_),
    .Y(_14167_));
 AO221x2_ASAP7_75t_R _19466_ (.A1(_14149_),
    .A2(_14154_),
    .B1(_14157_),
    .B2(_14160_),
    .C(_14167_),
    .Y(_14168_));
 INVx1_ASAP7_75t_R _19467_ (.A(_00484_),
    .Y(_14169_));
 NAND2x1_ASAP7_75t_R _19468_ (.A(net326),
    .B(_00482_),
    .Y(_14170_));
 OA21x2_ASAP7_75t_R _19469_ (.A1(net353),
    .A2(_14169_),
    .B(_14170_),
    .Y(_14171_));
 INVx1_ASAP7_75t_R _19470_ (.A(_00488_),
    .Y(_14172_));
 NAND2x1_ASAP7_75t_R _19471_ (.A(net326),
    .B(_00486_),
    .Y(_14173_));
 OA21x2_ASAP7_75t_R _19472_ (.A1(net326),
    .A2(_14172_),
    .B(_14173_),
    .Y(_14174_));
 AO221x1_ASAP7_75t_R _19473_ (.A1(_13184_),
    .A2(_14171_),
    .B1(_14174_),
    .B2(_13133_),
    .C(net321),
    .Y(_14175_));
 INVx1_ASAP7_75t_R _19474_ (.A(_00489_),
    .Y(_14176_));
 NAND2x1_ASAP7_75t_R _19475_ (.A(net322),
    .B(_00485_),
    .Y(_14177_));
 OA211x2_ASAP7_75t_R _19476_ (.A1(net322),
    .A2(_14176_),
    .B(_14177_),
    .C(net313),
    .Y(_14178_));
 INVx1_ASAP7_75t_R _19477_ (.A(_00487_),
    .Y(_14179_));
 NAND2x1_ASAP7_75t_R _19478_ (.A(net322),
    .B(_00483_),
    .Y(_14180_));
 OA211x2_ASAP7_75t_R _19479_ (.A1(net322),
    .A2(_14179_),
    .B(_14180_),
    .C(net326),
    .Y(_14181_));
 OA21x2_ASAP7_75t_R _19480_ (.A1(_14178_),
    .A2(_14181_),
    .B(net309),
    .Y(_14182_));
 INVx1_ASAP7_75t_R _19481_ (.A(_00476_),
    .Y(_14183_));
 INVx1_ASAP7_75t_R _19482_ (.A(_00477_),
    .Y(_14184_));
 NAND2x1_ASAP7_75t_R _19483_ (.A(net353),
    .B(_01703_),
    .Y(_14185_));
 OA21x2_ASAP7_75t_R _19484_ (.A1(net353),
    .A2(_14184_),
    .B(_14185_),
    .Y(_14186_));
 AO221x1_ASAP7_75t_R _19485_ (.A1(_14183_),
    .A2(_13190_),
    .B1(_14186_),
    .B2(net309),
    .C(_13584_),
    .Y(_14187_));
 NAND2x2_ASAP7_75t_R _19486_ (.A(_13132_),
    .B(net321),
    .Y(_14188_));
 INVx1_ASAP7_75t_R _19487_ (.A(_00480_),
    .Y(_14189_));
 NAND2x1_ASAP7_75t_R _19488_ (.A(net353),
    .B(_00478_),
    .Y(_14190_));
 OA211x2_ASAP7_75t_R _19489_ (.A1(net353),
    .A2(_14189_),
    .B(_14190_),
    .C(_00246_),
    .Y(_14191_));
 INVx1_ASAP7_75t_R _19490_ (.A(_00481_),
    .Y(_14192_));
 NAND2x1_ASAP7_75t_R _19491_ (.A(net353),
    .B(_00479_),
    .Y(_14193_));
 OA211x2_ASAP7_75t_R _19492_ (.A1(net353),
    .A2(_14192_),
    .B(_14193_),
    .C(net309),
    .Y(_14194_));
 OA31x2_ASAP7_75t_R _19493_ (.A1(_14188_),
    .A2(_14191_),
    .A3(_14194_),
    .B1(_00244_),
    .Y(_14195_));
 OA211x2_ASAP7_75t_R _19494_ (.A1(_14175_),
    .A2(_14182_),
    .B(_14187_),
    .C(_14195_),
    .Y(_14196_));
 OR2x6_ASAP7_75t_R _19495_ (.A(_14168_),
    .B(_14196_),
    .Y(_14197_));
 AND2x2_ASAP7_75t_R _19496_ (.A(_13583_),
    .B(_14197_),
    .Y(_14198_));
 AO21x2_ASAP7_75t_R _19497_ (.A1(_13299_),
    .A2(_14142_),
    .B(_14198_),
    .Y(_18135_));
 INVx1_ASAP7_75t_R _19498_ (.A(_18135_),
    .Y(_18137_));
 INVx2_ASAP7_75t_R _19499_ (.A(_01742_),
    .Y(_14199_));
 TIEHIx1_ASAP7_75t_R _34472__484 (.H(net484));
 INVx1_ASAP7_75t_R _19501_ (.A(_00526_),
    .Y(_14201_));
 NAND2x1_ASAP7_75t_R _19502_ (.A(net340),
    .B(_00524_),
    .Y(_14202_));
 OA211x2_ASAP7_75t_R _19503_ (.A1(net340),
    .A2(_14201_),
    .B(_14202_),
    .C(net359),
    .Y(_14203_));
 INVx1_ASAP7_75t_R _19504_ (.A(_00527_),
    .Y(_14204_));
 NAND2x1_ASAP7_75t_R _19505_ (.A(net340),
    .B(_00525_),
    .Y(_14205_));
 OA211x2_ASAP7_75t_R _19506_ (.A1(net340),
    .A2(_14204_),
    .B(_14205_),
    .C(net309),
    .Y(_14206_));
 OR3x1_ASAP7_75t_R _19507_ (.A(net323),
    .B(_14203_),
    .C(_14206_),
    .Y(_14207_));
 AND2x2_ASAP7_75t_R _19508_ (.A(net340),
    .B(_00520_),
    .Y(_14208_));
 AO21x1_ASAP7_75t_R _19509_ (.A1(net313),
    .A2(_00522_),
    .B(_14208_),
    .Y(_14209_));
 AND2x2_ASAP7_75t_R _19510_ (.A(net340),
    .B(_00521_),
    .Y(_14210_));
 AO21x1_ASAP7_75t_R _19511_ (.A1(net313),
    .A2(_00523_),
    .B(_14210_),
    .Y(_14211_));
 AOI221x1_ASAP7_75t_R _19512_ (.A1(_13184_),
    .A2(_14209_),
    .B1(_14211_),
    .B2(_13164_),
    .C(_13175_),
    .Y(_14212_));
 TIEHIx1_ASAP7_75t_R _34471__483 (.H(net483));
 AND2x2_ASAP7_75t_R _19514_ (.A(net340),
    .B(_00529_),
    .Y(_14214_));
 AO21x1_ASAP7_75t_R _19515_ (.A1(net313),
    .A2(_00531_),
    .B(_14214_),
    .Y(_14215_));
 AND3x1_ASAP7_75t_R _19516_ (.A(net357),
    .B(net340),
    .C(_00528_),
    .Y(_14216_));
 OR3x1_ASAP7_75t_R _19517_ (.A(_13132_),
    .B(_13976_),
    .C(_14216_),
    .Y(_14217_));
 AOI221x1_ASAP7_75t_R _19518_ (.A1(_00530_),
    .A2(_13190_),
    .B1(_14215_),
    .B2(net309),
    .C(_14217_),
    .Y(_14218_));
 INVx1_ASAP7_75t_R _19519_ (.A(_00535_),
    .Y(_14219_));
 NAND2x1_ASAP7_75t_R _19520_ (.A(net340),
    .B(_00533_),
    .Y(_14220_));
 OA211x2_ASAP7_75t_R _19521_ (.A1(net340),
    .A2(_14219_),
    .B(_14220_),
    .C(net309),
    .Y(_14221_));
 INVx1_ASAP7_75t_R _19522_ (.A(_00534_),
    .Y(_14222_));
 NAND2x1_ASAP7_75t_R _19523_ (.A(net340),
    .B(_00532_),
    .Y(_14223_));
 OA211x2_ASAP7_75t_R _19524_ (.A1(net340),
    .A2(_14222_),
    .B(_14223_),
    .C(net359),
    .Y(_14224_));
 OA21x2_ASAP7_75t_R _19525_ (.A1(_14221_),
    .A2(_14224_),
    .B(_14134_),
    .Y(_14225_));
 AO211x2_ASAP7_75t_R _19526_ (.A1(_14207_),
    .A2(_14212_),
    .B(_14218_),
    .C(_14225_),
    .Y(_14226_));
 INVx1_ASAP7_75t_R _19527_ (.A(_00514_),
    .Y(_14227_));
 NAND2x1_ASAP7_75t_R _19528_ (.A(net341),
    .B(_00512_),
    .Y(_14228_));
 OA21x2_ASAP7_75t_R _19529_ (.A1(net341),
    .A2(_14227_),
    .B(_14228_),
    .Y(_14229_));
 INVx1_ASAP7_75t_R _19530_ (.A(_00518_),
    .Y(_14230_));
 NAND2x1_ASAP7_75t_R _19531_ (.A(net341),
    .B(_00516_),
    .Y(_14231_));
 OA21x2_ASAP7_75t_R _19532_ (.A1(net341),
    .A2(_14230_),
    .B(_14231_),
    .Y(_14232_));
 AO221x1_ASAP7_75t_R _19533_ (.A1(_13184_),
    .A2(_14229_),
    .B1(_14232_),
    .B2(_13133_),
    .C(net320),
    .Y(_14233_));
 INVx1_ASAP7_75t_R _19534_ (.A(_00519_),
    .Y(_14234_));
 NAND2x1_ASAP7_75t_R _19535_ (.A(net323),
    .B(_00515_),
    .Y(_14235_));
 OA211x2_ASAP7_75t_R _19536_ (.A1(net323),
    .A2(_14234_),
    .B(_14235_),
    .C(net313),
    .Y(_14236_));
 INVx1_ASAP7_75t_R _19537_ (.A(_00517_),
    .Y(_14237_));
 NAND2x1_ASAP7_75t_R _19538_ (.A(_01744_),
    .B(_00513_),
    .Y(_14238_));
 OA211x2_ASAP7_75t_R _19539_ (.A1(_01744_),
    .A2(_14237_),
    .B(_14238_),
    .C(net351),
    .Y(_14239_));
 OA21x2_ASAP7_75t_R _19540_ (.A1(_14236_),
    .A2(_14239_),
    .B(net309),
    .Y(_14240_));
 INVx1_ASAP7_75t_R _19541_ (.A(_00510_),
    .Y(_14241_));
 NAND2x1_ASAP7_75t_R _19542_ (.A(net351),
    .B(_00508_),
    .Y(_14242_));
 OA211x2_ASAP7_75t_R _19543_ (.A1(net351),
    .A2(_14241_),
    .B(_14242_),
    .C(net360),
    .Y(_14243_));
 INVx1_ASAP7_75t_R _19544_ (.A(_00511_),
    .Y(_14244_));
 NAND2x1_ASAP7_75t_R _19545_ (.A(net351),
    .B(_00509_),
    .Y(_14245_));
 OA211x2_ASAP7_75t_R _19546_ (.A1(net351),
    .A2(_14244_),
    .B(_14245_),
    .C(net309),
    .Y(_14246_));
 OR3x1_ASAP7_75t_R _19547_ (.A(_14188_),
    .B(_14243_),
    .C(_14246_),
    .Y(_14247_));
 INVx1_ASAP7_75t_R _19548_ (.A(_00507_),
    .Y(_14248_));
 NAND2x1_ASAP7_75t_R _19549_ (.A(net339),
    .B(_01702_),
    .Y(_14249_));
 OA211x2_ASAP7_75t_R _19550_ (.A1(net339),
    .A2(_14248_),
    .B(_14249_),
    .C(net309),
    .Y(_14250_));
 INVx1_ASAP7_75t_R _19551_ (.A(_00506_),
    .Y(_14251_));
 AND3x1_ASAP7_75t_R _19552_ (.A(net359),
    .B(net313),
    .C(_14251_),
    .Y(_14252_));
 OA31x2_ASAP7_75t_R _19553_ (.A1(_13584_),
    .A2(_14250_),
    .A3(_14252_),
    .B1(net315),
    .Y(_14253_));
 OA211x2_ASAP7_75t_R _19554_ (.A1(_14233_),
    .A2(_14240_),
    .B(_14247_),
    .C(_14253_),
    .Y(_14254_));
 OA21x2_ASAP7_75t_R _19555_ (.A1(_14226_),
    .A2(_14254_),
    .B(_13583_),
    .Y(_14255_));
 AO21x2_ASAP7_75t_R _19556_ (.A1(_14199_),
    .A2(_14138_),
    .B(_14255_),
    .Y(_14256_));
 TIEHIx1_ASAP7_75t_R _34470__482 (.H(net482));
 INVx1_ASAP7_75t_R _19558_ (.A(_14256_),
    .Y(_18142_));
 TIEHIx1_ASAP7_75t_R _34469__481 (.H(net481));
 TIEHIx1_ASAP7_75t_R _34468__480 (.H(net480));
 INVx1_ASAP7_75t_R _19561_ (.A(_00556_),
    .Y(_14259_));
 TIEHIx1_ASAP7_75t_R _34467__479 (.H(net479));
 NAND2x1_ASAP7_75t_R _19563_ (.A(net352),
    .B(_00554_),
    .Y(_14261_));
 OA211x2_ASAP7_75t_R _19564_ (.A1(net352),
    .A2(_14259_),
    .B(_13133_),
    .C(_14261_),
    .Y(_14262_));
 INVx1_ASAP7_75t_R _19565_ (.A(_00553_),
    .Y(_14263_));
 TIEHIx1_ASAP7_75t_R _34466__478 (.H(net478));
 NAND2x1_ASAP7_75t_R _19567_ (.A(net352),
    .B(_00551_),
    .Y(_14265_));
 OA211x2_ASAP7_75t_R _19568_ (.A1(net352),
    .A2(_14263_),
    .B(_13164_),
    .C(_14265_),
    .Y(_14266_));
 TIEHIx1_ASAP7_75t_R _34465__477 (.H(net477));
 INVx1_ASAP7_75t_R _19570_ (.A(_00552_),
    .Y(_14268_));
 NAND2x1_ASAP7_75t_R _19571_ (.A(net352),
    .B(_00550_),
    .Y(_14269_));
 OA211x2_ASAP7_75t_R _19572_ (.A1(net352),
    .A2(_14268_),
    .B(_13184_),
    .C(_14269_),
    .Y(_14270_));
 INVx1_ASAP7_75t_R _19573_ (.A(_00557_),
    .Y(_14271_));
 NAND2x1_ASAP7_75t_R _19574_ (.A(net352),
    .B(_00555_),
    .Y(_14272_));
 OA211x2_ASAP7_75t_R _19575_ (.A1(net352),
    .A2(_14271_),
    .B(_13124_),
    .C(_14272_),
    .Y(_14273_));
 OR4x1_ASAP7_75t_R _19576_ (.A(_14262_),
    .B(_14266_),
    .C(_14270_),
    .D(_14273_),
    .Y(_14274_));
 INVx1_ASAP7_75t_R _19577_ (.A(_00560_),
    .Y(_14275_));
 NAND2x1_ASAP7_75t_R _19578_ (.A(net350),
    .B(_00558_),
    .Y(_14276_));
 OA211x2_ASAP7_75t_R _19579_ (.A1(net350),
    .A2(_14275_),
    .B(_13184_),
    .C(_14276_),
    .Y(_14277_));
 INVx1_ASAP7_75t_R _19580_ (.A(_00561_),
    .Y(_14278_));
 NAND2x1_ASAP7_75t_R _19581_ (.A(net350),
    .B(_00559_),
    .Y(_14279_));
 OA211x2_ASAP7_75t_R _19582_ (.A1(net350),
    .A2(_14278_),
    .B(_13164_),
    .C(_14279_),
    .Y(_14280_));
 INVx1_ASAP7_75t_R _19583_ (.A(_00565_),
    .Y(_14281_));
 NAND2x1_ASAP7_75t_R _19584_ (.A(net350),
    .B(_00563_),
    .Y(_14282_));
 OA211x2_ASAP7_75t_R _19585_ (.A1(net350),
    .A2(_14281_),
    .B(_13124_),
    .C(_14282_),
    .Y(_14283_));
 INVx1_ASAP7_75t_R _19586_ (.A(_00564_),
    .Y(_14284_));
 NAND2x1_ASAP7_75t_R _19587_ (.A(net350),
    .B(_00562_),
    .Y(_14285_));
 OA211x2_ASAP7_75t_R _19588_ (.A1(net350),
    .A2(_14284_),
    .B(_13133_),
    .C(_14285_),
    .Y(_14286_));
 OR4x1_ASAP7_75t_R _19589_ (.A(_14277_),
    .B(_14280_),
    .C(_14283_),
    .D(_14286_),
    .Y(_14287_));
 INVx1_ASAP7_75t_R _19590_ (.A(_00549_),
    .Y(_14288_));
 NAND2x1_ASAP7_75t_R _19591_ (.A(net352),
    .B(_00547_),
    .Y(_14289_));
 OA211x2_ASAP7_75t_R _19592_ (.A1(net352),
    .A2(_14288_),
    .B(_14289_),
    .C(net310),
    .Y(_14290_));
 INVx1_ASAP7_75t_R _19593_ (.A(_00548_),
    .Y(_14291_));
 NAND2x1_ASAP7_75t_R _19594_ (.A(net352),
    .B(_00546_),
    .Y(_14292_));
 OA211x2_ASAP7_75t_R _19595_ (.A1(net352),
    .A2(_14291_),
    .B(_14292_),
    .C(net361),
    .Y(_14293_));
 OA21x2_ASAP7_75t_R _19596_ (.A1(_14290_),
    .A2(_14293_),
    .B(_13132_),
    .Y(_14294_));
 TIEHIx1_ASAP7_75t_R _34464__476 (.H(net476));
 AND2x2_ASAP7_75t_R _19598_ (.A(net361),
    .B(_00542_),
    .Y(_14296_));
 AOI21x1_ASAP7_75t_R _19599_ (.A1(net310),
    .A2(_00543_),
    .B(_14296_),
    .Y(_14297_));
 INVx1_ASAP7_75t_R _19600_ (.A(_00545_),
    .Y(_14298_));
 NAND2x1_ASAP7_75t_R _19601_ (.A(net361),
    .B(_00544_),
    .Y(_14299_));
 OA21x2_ASAP7_75t_R _19602_ (.A1(net361),
    .A2(_14298_),
    .B(_14299_),
    .Y(_14300_));
 AO221x1_ASAP7_75t_R _19603_ (.A1(_13933_),
    .A2(_14297_),
    .B1(_14300_),
    .B2(_13940_),
    .C(_00245_),
    .Y(_14301_));
 INVx1_ASAP7_75t_R _19604_ (.A(_00541_),
    .Y(_14302_));
 NAND2x1_ASAP7_75t_R _19605_ (.A(net352),
    .B(_00539_),
    .Y(_14303_));
 OA211x2_ASAP7_75t_R _19606_ (.A1(net352),
    .A2(_14302_),
    .B(_14303_),
    .C(net309),
    .Y(_14304_));
 INVx1_ASAP7_75t_R _19607_ (.A(_00540_),
    .Y(_14305_));
 NAND2x1_ASAP7_75t_R _19608_ (.A(net352),
    .B(_00538_),
    .Y(_14306_));
 OA211x2_ASAP7_75t_R _19609_ (.A1(net352),
    .A2(_14305_),
    .B(_14306_),
    .C(net361),
    .Y(_14307_));
 OR3x1_ASAP7_75t_R _19610_ (.A(_14188_),
    .B(_14304_),
    .C(_14307_),
    .Y(_14308_));
 INVx1_ASAP7_75t_R _19611_ (.A(_00537_),
    .Y(_14309_));
 NAND2x1_ASAP7_75t_R _19612_ (.A(net352),
    .B(_01701_),
    .Y(_14310_));
 OA211x2_ASAP7_75t_R _19613_ (.A1(net352),
    .A2(_14309_),
    .B(_14310_),
    .C(net310),
    .Y(_14311_));
 INVx1_ASAP7_75t_R _19614_ (.A(_00536_),
    .Y(_14312_));
 AND3x1_ASAP7_75t_R _19615_ (.A(net361),
    .B(net313),
    .C(_14312_),
    .Y(_14313_));
 OA31x2_ASAP7_75t_R _19616_ (.A1(_13584_),
    .A2(_14311_),
    .A3(_14313_),
    .B1(net314),
    .Y(_14314_));
 OA211x2_ASAP7_75t_R _19617_ (.A1(_14294_),
    .A2(_14301_),
    .B(_14308_),
    .C(_14314_),
    .Y(_14315_));
 AO221x2_ASAP7_75t_R _19618_ (.A1(_13614_),
    .A2(_14274_),
    .B1(_14287_),
    .B2(_13215_),
    .C(_14315_),
    .Y(_14316_));
 TIEHIx1_ASAP7_75t_R _34463__475 (.H(net475));
 INVx2_ASAP7_75t_R _19620_ (.A(_01741_),
    .Y(_14318_));
 AO32x2_ASAP7_75t_R _19621_ (.A1(_13223_),
    .A2(_13248_),
    .A3(_14316_),
    .B1(_14138_),
    .B2(_14318_),
    .Y(_14319_));
 TIEHIx1_ASAP7_75t_R _34462__474 (.H(net474));
 INVx2_ASAP7_75t_R _19623_ (.A(_14319_),
    .Y(_18147_));
 AO221x1_ASAP7_75t_R _19624_ (.A1(_00594_),
    .A2(_13190_),
    .B1(_14155_),
    .B2(_00592_),
    .C(_14156_),
    .Y(_14320_));
 TIEHIx1_ASAP7_75t_R _34461__473 (.H(net473));
 OR2x2_ASAP7_75t_R _19626_ (.A(net353),
    .B(_00595_),
    .Y(_14322_));
 OA211x2_ASAP7_75t_R _19627_ (.A1(net313),
    .A2(_00593_),
    .B(_14322_),
    .C(net309),
    .Y(_14323_));
 NOR2x1_ASAP7_75t_R _19628_ (.A(_14320_),
    .B(_14323_),
    .Y(_14324_));
 INVx1_ASAP7_75t_R _19629_ (.A(_00579_),
    .Y(_14325_));
 NAND2x1_ASAP7_75t_R _19630_ (.A(net322),
    .B(_00575_),
    .Y(_14326_));
 OA211x2_ASAP7_75t_R _19631_ (.A1(net322),
    .A2(_14325_),
    .B(_14326_),
    .C(net313),
    .Y(_14327_));
 INVx1_ASAP7_75t_R _19632_ (.A(_00577_),
    .Y(_14328_));
 NAND2x1_ASAP7_75t_R _19633_ (.A(net322),
    .B(_00573_),
    .Y(_14329_));
 OA211x2_ASAP7_75t_R _19634_ (.A1(net322),
    .A2(_14328_),
    .B(_14329_),
    .C(net330),
    .Y(_14330_));
 OA21x2_ASAP7_75t_R _19635_ (.A1(_14327_),
    .A2(_14330_),
    .B(net310),
    .Y(_14331_));
 INVx1_ASAP7_75t_R _19636_ (.A(_00574_),
    .Y(_14332_));
 NAND2x1_ASAP7_75t_R _19637_ (.A(net326),
    .B(_00572_),
    .Y(_14333_));
 OA21x2_ASAP7_75t_R _19638_ (.A1(net326),
    .A2(_14332_),
    .B(_14333_),
    .Y(_14334_));
 INVx1_ASAP7_75t_R _19639_ (.A(_00578_),
    .Y(_14335_));
 NAND2x1_ASAP7_75t_R _19640_ (.A(net326),
    .B(_00576_),
    .Y(_14336_));
 OA21x2_ASAP7_75t_R _19641_ (.A1(net326),
    .A2(_14335_),
    .B(_14336_),
    .Y(_14337_));
 AO221x1_ASAP7_75t_R _19642_ (.A1(_13184_),
    .A2(_14334_),
    .B1(_14337_),
    .B2(_13133_),
    .C(net321),
    .Y(_14338_));
 INVx1_ASAP7_75t_R _19643_ (.A(_00570_),
    .Y(_14339_));
 NAND2x1_ASAP7_75t_R _19644_ (.A(net326),
    .B(_00568_),
    .Y(_14340_));
 OA211x2_ASAP7_75t_R _19645_ (.A1(net326),
    .A2(_14339_),
    .B(_14340_),
    .C(_00246_),
    .Y(_14341_));
 INVx1_ASAP7_75t_R _19646_ (.A(_00571_),
    .Y(_14342_));
 NAND2x1_ASAP7_75t_R _19647_ (.A(net326),
    .B(_00569_),
    .Y(_14343_));
 OA211x2_ASAP7_75t_R _19648_ (.A1(net326),
    .A2(_14342_),
    .B(_14343_),
    .C(net310),
    .Y(_14344_));
 OR3x1_ASAP7_75t_R _19649_ (.A(_14188_),
    .B(_14341_),
    .C(_14344_),
    .Y(_14345_));
 INVx1_ASAP7_75t_R _19650_ (.A(_00567_),
    .Y(_14346_));
 NAND2x1_ASAP7_75t_R _19651_ (.A(net330),
    .B(_01700_),
    .Y(_14347_));
 OA211x2_ASAP7_75t_R _19652_ (.A1(net330),
    .A2(_14346_),
    .B(_14347_),
    .C(net310),
    .Y(_14348_));
 NOR2x1_ASAP7_75t_R _19653_ (.A(net330),
    .B(_00566_),
    .Y(_14349_));
 AO21x1_ASAP7_75t_R _19654_ (.A1(_00246_),
    .A2(_14349_),
    .B(_13584_),
    .Y(_14350_));
 OA21x2_ASAP7_75t_R _19655_ (.A1(_14348_),
    .A2(_14350_),
    .B(_00244_),
    .Y(_14351_));
 OA211x2_ASAP7_75t_R _19656_ (.A1(_14331_),
    .A2(_14338_),
    .B(_14345_),
    .C(_14351_),
    .Y(_14352_));
 INVx1_ASAP7_75t_R _19657_ (.A(_00590_),
    .Y(_14353_));
 NAND2x1_ASAP7_75t_R _19658_ (.A(net310),
    .B(_00591_),
    .Y(_14354_));
 OA211x2_ASAP7_75t_R _19659_ (.A1(net310),
    .A2(_14353_),
    .B(_13940_),
    .C(_14354_),
    .Y(_14355_));
 INVx1_ASAP7_75t_R _19660_ (.A(_00589_),
    .Y(_14356_));
 NAND2x1_ASAP7_75t_R _19661_ (.A(net361),
    .B(_00588_),
    .Y(_14357_));
 OA211x2_ASAP7_75t_R _19662_ (.A1(net361),
    .A2(_14356_),
    .B(_13933_),
    .C(_14357_),
    .Y(_14358_));
 OA21x2_ASAP7_75t_R _19663_ (.A1(_14355_),
    .A2(_14358_),
    .B(_13215_),
    .Y(_14359_));
 INVx1_ASAP7_75t_R _19664_ (.A(_00587_),
    .Y(_14360_));
 NAND2x1_ASAP7_75t_R _19665_ (.A(net330),
    .B(_00585_),
    .Y(_14361_));
 OA21x2_ASAP7_75t_R _19666_ (.A1(net330),
    .A2(_14360_),
    .B(_14361_),
    .Y(_14362_));
 INVx1_ASAP7_75t_R _19667_ (.A(_00582_),
    .Y(_14363_));
 NAND2x1_ASAP7_75t_R _19668_ (.A(net330),
    .B(_00580_),
    .Y(_14364_));
 OA211x2_ASAP7_75t_R _19669_ (.A1(net330),
    .A2(_14363_),
    .B(_13184_),
    .C(_14364_),
    .Y(_14365_));
 AO21x1_ASAP7_75t_R _19670_ (.A1(_13124_),
    .A2(_14362_),
    .B(_14365_),
    .Y(_14366_));
 NAND2x1_ASAP7_75t_R _19671_ (.A(net330),
    .B(_00584_),
    .Y(_14367_));
 NAND2x1_ASAP7_75t_R _19672_ (.A(net313),
    .B(_00586_),
    .Y(_14368_));
 NAND2x1_ASAP7_75t_R _19673_ (.A(net353),
    .B(_00581_),
    .Y(_14369_));
 NAND2x1_ASAP7_75t_R _19674_ (.A(net313),
    .B(_00583_),
    .Y(_14370_));
 AO33x2_ASAP7_75t_R _19675_ (.A1(_13133_),
    .A2(_14367_),
    .A3(_14368_),
    .B1(_14369_),
    .B2(_14370_),
    .B3(_13164_),
    .Y(_14371_));
 OA21x2_ASAP7_75t_R _19676_ (.A1(_14366_),
    .A2(_14371_),
    .B(_13614_),
    .Y(_14372_));
 OR4x2_ASAP7_75t_R _19677_ (.A(_14324_),
    .B(_14352_),
    .C(_14359_),
    .D(_14372_),
    .Y(_14373_));
 TIEHIx1_ASAP7_75t_R _34460__472 (.H(net472));
 INVx2_ASAP7_75t_R _19679_ (.A(_01740_),
    .Y(_14375_));
 AO32x2_ASAP7_75t_R _19680_ (.A1(_13223_),
    .A2(_13248_),
    .A3(_14373_),
    .B1(_14138_),
    .B2(_14375_),
    .Y(_14376_));
 TIEHIx1_ASAP7_75t_R _34459__471 (.H(net471));
 INVx1_ASAP7_75t_R _19682_ (.A(_14376_),
    .Y(_18152_));
 INVx1_ASAP7_75t_R _19683_ (.A(_00605_),
    .Y(_14377_));
 TIEHIx1_ASAP7_75t_R _34458__470 (.H(net470));
 NAND2x1_ASAP7_75t_R _19685_ (.A(net340),
    .B(_00603_),
    .Y(_14379_));
 OA211x2_ASAP7_75t_R _19686_ (.A1(net340),
    .A2(_14377_),
    .B(_14379_),
    .C(net309),
    .Y(_14380_));
 INVx1_ASAP7_75t_R _19687_ (.A(_00604_),
    .Y(_14381_));
 NAND2x1_ASAP7_75t_R _19688_ (.A(net340),
    .B(_00602_),
    .Y(_14382_));
 TIEHIx1_ASAP7_75t_R _34457__469 (.H(net469));
 OA211x2_ASAP7_75t_R _19690_ (.A1(net340),
    .A2(_14381_),
    .B(_14382_),
    .C(net357),
    .Y(_14384_));
 OAI21x1_ASAP7_75t_R _19691_ (.A1(_14380_),
    .A2(_14384_),
    .B(net324),
    .Y(_14385_));
 INVx1_ASAP7_75t_R _19692_ (.A(_00606_),
    .Y(_14386_));
 TIEHIx1_ASAP7_75t_R _34456__468 (.H(net468));
 NOR2x1_ASAP7_75t_R _19694_ (.A(net340),
    .B(_00608_),
    .Y(_14388_));
 AO21x1_ASAP7_75t_R _19695_ (.A1(net340),
    .A2(_14386_),
    .B(_14388_),
    .Y(_14389_));
 INVx1_ASAP7_75t_R _19696_ (.A(_00609_),
    .Y(_14390_));
 NAND2x1_ASAP7_75t_R _19697_ (.A(net340),
    .B(_00607_),
    .Y(_14391_));
 OA211x2_ASAP7_75t_R _19698_ (.A1(net340),
    .A2(_14390_),
    .B(_13124_),
    .C(_14391_),
    .Y(_14392_));
 AOI21x1_ASAP7_75t_R _19699_ (.A1(_13133_),
    .A2(_14389_),
    .B(_14392_),
    .Y(_14393_));
 AND3x1_ASAP7_75t_R _19700_ (.A(_13598_),
    .B(_14385_),
    .C(_14393_),
    .Y(_14394_));
 INVx1_ASAP7_75t_R _19701_ (.A(_00601_),
    .Y(_14395_));
 NAND2x1_ASAP7_75t_R _19702_ (.A(net340),
    .B(_00599_),
    .Y(_14396_));
 OA211x2_ASAP7_75t_R _19703_ (.A1(net340),
    .A2(_14395_),
    .B(_14396_),
    .C(net309),
    .Y(_14397_));
 INVx1_ASAP7_75t_R _19704_ (.A(_00600_),
    .Y(_14398_));
 NAND2x1_ASAP7_75t_R _19705_ (.A(net340),
    .B(_00598_),
    .Y(_14399_));
 OA211x2_ASAP7_75t_R _19706_ (.A1(net340),
    .A2(_14398_),
    .B(_14399_),
    .C(net357),
    .Y(_14400_));
 OR3x1_ASAP7_75t_R _19707_ (.A(_14188_),
    .B(_14397_),
    .C(_14400_),
    .Y(_14401_));
 INVx1_ASAP7_75t_R _19708_ (.A(_00596_),
    .Y(_14402_));
 INVx1_ASAP7_75t_R _19709_ (.A(_00597_),
    .Y(_14403_));
 NAND2x1_ASAP7_75t_R _19710_ (.A(net346),
    .B(_01699_),
    .Y(_14404_));
 OA21x2_ASAP7_75t_R _19711_ (.A1(net346),
    .A2(_14403_),
    .B(_14404_),
    .Y(_14405_));
 AO221x1_ASAP7_75t_R _19712_ (.A1(_14402_),
    .A2(_13190_),
    .B1(_14405_),
    .B2(net310),
    .C(_13584_),
    .Y(_14406_));
 NAND3x1_ASAP7_75t_R _19713_ (.A(net314),
    .B(_14401_),
    .C(_14406_),
    .Y(_14407_));
 TIEHIx1_ASAP7_75t_R _34455__467 (.H(net467));
 INVx1_ASAP7_75t_R _19715_ (.A(_00621_),
    .Y(_14409_));
 NAND2x1_ASAP7_75t_R _19716_ (.A(net347),
    .B(_00619_),
    .Y(_14410_));
 OA21x2_ASAP7_75t_R _19717_ (.A1(net347),
    .A2(_14409_),
    .B(_14410_),
    .Y(_14411_));
 INVx1_ASAP7_75t_R _19718_ (.A(_00620_),
    .Y(_14412_));
 NAND2x1_ASAP7_75t_R _19719_ (.A(net347),
    .B(_00618_),
    .Y(_14413_));
 OA211x2_ASAP7_75t_R _19720_ (.A1(net347),
    .A2(_14412_),
    .B(_14413_),
    .C(net357),
    .Y(_14414_));
 AOI211x1_ASAP7_75t_R _19721_ (.A1(net310),
    .A2(_14411_),
    .B(_14414_),
    .C(_13132_),
    .Y(_14415_));
 AND2x2_ASAP7_75t_R _19722_ (.A(net347),
    .B(_00623_),
    .Y(_14416_));
 AO21x1_ASAP7_75t_R _19723_ (.A1(net312),
    .A2(_00625_),
    .B(_14416_),
    .Y(_14417_));
 AND2x2_ASAP7_75t_R _19724_ (.A(net347),
    .B(_00622_),
    .Y(_14418_));
 AO21x1_ASAP7_75t_R _19725_ (.A1(net312),
    .A2(_00624_),
    .B(_14418_),
    .Y(_14419_));
 AO22x1_ASAP7_75t_R _19726_ (.A1(_13124_),
    .A2(_14417_),
    .B1(_14419_),
    .B2(_13133_),
    .Y(_14420_));
 INVx1_ASAP7_75t_R _19727_ (.A(_00617_),
    .Y(_14421_));
 NAND2x1_ASAP7_75t_R _19728_ (.A(net346),
    .B(_00615_),
    .Y(_14422_));
 OA21x2_ASAP7_75t_R _19729_ (.A1(net346),
    .A2(_14421_),
    .B(_14422_),
    .Y(_14423_));
 INVx1_ASAP7_75t_R _19730_ (.A(_00616_),
    .Y(_14424_));
 NAND2x1_ASAP7_75t_R _19731_ (.A(net346),
    .B(_00614_),
    .Y(_14425_));
 OA211x2_ASAP7_75t_R _19732_ (.A1(net346),
    .A2(_14424_),
    .B(_14425_),
    .C(net357),
    .Y(_14426_));
 AOI211x1_ASAP7_75t_R _19733_ (.A1(net310),
    .A2(_14423_),
    .B(_14426_),
    .C(net324),
    .Y(_14427_));
 AND2x2_ASAP7_75t_R _19734_ (.A(net347),
    .B(_00610_),
    .Y(_14428_));
 AO21x1_ASAP7_75t_R _19735_ (.A1(net312),
    .A2(_00612_),
    .B(_14428_),
    .Y(_14429_));
 AND2x2_ASAP7_75t_R _19736_ (.A(net347),
    .B(_00611_),
    .Y(_14430_));
 AO21x1_ASAP7_75t_R _19737_ (.A1(net312),
    .A2(_00613_),
    .B(_14430_),
    .Y(_14431_));
 AO22x1_ASAP7_75t_R _19738_ (.A1(_13184_),
    .A2(_14429_),
    .B1(_14431_),
    .B2(_13164_),
    .Y(_14432_));
 OA33x2_ASAP7_75t_R _19739_ (.A1(_13976_),
    .A2(_14415_),
    .A3(_14420_),
    .B1(_14427_),
    .B2(_14432_),
    .B3(_13175_),
    .Y(_14433_));
 OAI21x1_ASAP7_75t_R _19740_ (.A1(_14394_),
    .A2(_14407_),
    .B(_14433_),
    .Y(_14434_));
 NAND2x2_ASAP7_75t_R _19741_ (.A(_13583_),
    .B(_14434_),
    .Y(_14435_));
 NAND2x2_ASAP7_75t_R _19742_ (.A(_13223_),
    .B(_13291_),
    .Y(_14436_));
 AO21x1_ASAP7_75t_R _19743_ (.A1(_13298_),
    .A2(_14436_),
    .B(_13275_),
    .Y(_14437_));
 OR3x1_ASAP7_75t_R _19744_ (.A(_01739_),
    .B(_13583_),
    .C(_14437_),
    .Y(_14438_));
 NAND2x2_ASAP7_75t_R _19745_ (.A(_14435_),
    .B(_14438_),
    .Y(_18155_));
 INVx1_ASAP7_75t_R _19746_ (.A(_18155_),
    .Y(_18157_));
 INVx1_ASAP7_75t_R _19747_ (.A(_00638_),
    .Y(_14439_));
 NAND2x1_ASAP7_75t_R _19748_ (.A(net330),
    .B(_00636_),
    .Y(_14440_));
 OA21x2_ASAP7_75t_R _19749_ (.A1(net330),
    .A2(_14439_),
    .B(_14440_),
    .Y(_14441_));
 INVx1_ASAP7_75t_R _19750_ (.A(_00634_),
    .Y(_14442_));
 NAND2x1_ASAP7_75t_R _19751_ (.A(net330),
    .B(_00632_),
    .Y(_14443_));
 OA211x2_ASAP7_75t_R _19752_ (.A1(net330),
    .A2(_14442_),
    .B(_13184_),
    .C(_14443_),
    .Y(_14444_));
 AO21x1_ASAP7_75t_R _19753_ (.A1(_13133_),
    .A2(_14441_),
    .B(_14444_),
    .Y(_14445_));
 INVx1_ASAP7_75t_R _19754_ (.A(_00639_),
    .Y(_14446_));
 NAND2x1_ASAP7_75t_R _19755_ (.A(net330),
    .B(_00637_),
    .Y(_14447_));
 OA211x2_ASAP7_75t_R _19756_ (.A1(net330),
    .A2(_14446_),
    .B(_13124_),
    .C(_14447_),
    .Y(_14448_));
 INVx1_ASAP7_75t_R _19757_ (.A(_00635_),
    .Y(_14449_));
 NAND2x1_ASAP7_75t_R _19758_ (.A(net349),
    .B(_00633_),
    .Y(_14450_));
 OA211x2_ASAP7_75t_R _19759_ (.A1(net349),
    .A2(_14449_),
    .B(_13164_),
    .C(_14450_),
    .Y(_14451_));
 OR4x1_ASAP7_75t_R _19760_ (.A(net321),
    .B(_14445_),
    .C(_14448_),
    .D(_14451_),
    .Y(_14452_));
 AND2x2_ASAP7_75t_R _19761_ (.A(net348),
    .B(_00628_),
    .Y(_14453_));
 AO21x1_ASAP7_75t_R _19762_ (.A1(net312),
    .A2(_00630_),
    .B(_14453_),
    .Y(_14454_));
 AND2x2_ASAP7_75t_R _19763_ (.A(net350),
    .B(_00629_),
    .Y(_14455_));
 AO21x1_ASAP7_75t_R _19764_ (.A1(net312),
    .A2(_00631_),
    .B(_14455_),
    .Y(_14456_));
 AOI22x1_ASAP7_75t_R _19765_ (.A1(_13133_),
    .A2(_14454_),
    .B1(_14456_),
    .B2(_13124_),
    .Y(_14457_));
 INVx1_ASAP7_75t_R _19766_ (.A(_00626_),
    .Y(_14458_));
 INVx1_ASAP7_75t_R _19767_ (.A(_00627_),
    .Y(_14459_));
 NAND2x1_ASAP7_75t_R _19768_ (.A(net348),
    .B(_01698_),
    .Y(_14460_));
 OA21x2_ASAP7_75t_R _19769_ (.A1(net348),
    .A2(_14459_),
    .B(_14460_),
    .Y(_14461_));
 AO221x1_ASAP7_75t_R _19770_ (.A1(_14458_),
    .A2(_13190_),
    .B1(_14461_),
    .B2(net310),
    .C(_13584_),
    .Y(_14462_));
 OA211x2_ASAP7_75t_R _19771_ (.A1(_13598_),
    .A2(_14457_),
    .B(_14462_),
    .C(net314),
    .Y(_14463_));
 INVx1_ASAP7_75t_R _19772_ (.A(_00643_),
    .Y(_14464_));
 NAND2x1_ASAP7_75t_R _19773_ (.A(net350),
    .B(_00641_),
    .Y(_14465_));
 OA211x2_ASAP7_75t_R _19774_ (.A1(net350),
    .A2(_14464_),
    .B(_13164_),
    .C(_14465_),
    .Y(_14466_));
 INVx1_ASAP7_75t_R _19775_ (.A(_00642_),
    .Y(_14467_));
 NAND2x1_ASAP7_75t_R _19776_ (.A(net350),
    .B(_00640_),
    .Y(_14468_));
 OA211x2_ASAP7_75t_R _19777_ (.A1(net350),
    .A2(_14467_),
    .B(_13184_),
    .C(_14468_),
    .Y(_14469_));
 INVx1_ASAP7_75t_R _19778_ (.A(_00646_),
    .Y(_14470_));
 NAND2x1_ASAP7_75t_R _19779_ (.A(net350),
    .B(_00644_),
    .Y(_14471_));
 OA211x2_ASAP7_75t_R _19780_ (.A1(net350),
    .A2(_14470_),
    .B(_13133_),
    .C(_14471_),
    .Y(_14472_));
 INVx1_ASAP7_75t_R _19781_ (.A(_00647_),
    .Y(_14473_));
 NAND2x1_ASAP7_75t_R _19782_ (.A(net350),
    .B(_00645_),
    .Y(_14474_));
 OA211x2_ASAP7_75t_R _19783_ (.A1(net350),
    .A2(_14473_),
    .B(_13124_),
    .C(_14474_),
    .Y(_14475_));
 OR4x1_ASAP7_75t_R _19784_ (.A(_14466_),
    .B(_14469_),
    .C(_14472_),
    .D(_14475_),
    .Y(_14476_));
 INVx1_ASAP7_75t_R _19785_ (.A(_00650_),
    .Y(_14477_));
 NOR2x1_ASAP7_75t_R _19786_ (.A(net360),
    .B(_00651_),
    .Y(_14478_));
 AO21x1_ASAP7_75t_R _19787_ (.A1(net360),
    .A2(_14477_),
    .B(_14478_),
    .Y(_14479_));
 INVx1_ASAP7_75t_R _19788_ (.A(_00649_),
    .Y(_14480_));
 NAND2x1_ASAP7_75t_R _19789_ (.A(net359),
    .B(_00648_),
    .Y(_14481_));
 OA211x2_ASAP7_75t_R _19790_ (.A1(net359),
    .A2(_14480_),
    .B(_13933_),
    .C(_14481_),
    .Y(_14482_));
 AO21x1_ASAP7_75t_R _19791_ (.A1(_13940_),
    .A2(_14479_),
    .B(_14482_),
    .Y(_14483_));
 AND2x2_ASAP7_75t_R _19792_ (.A(net352),
    .B(_00653_),
    .Y(_14484_));
 AO21x1_ASAP7_75t_R _19793_ (.A1(net313),
    .A2(_00655_),
    .B(_14484_),
    .Y(_14485_));
 AO21x1_ASAP7_75t_R _19794_ (.A1(_00652_),
    .A2(_14155_),
    .B(_14156_),
    .Y(_14486_));
 AOI221x1_ASAP7_75t_R _19795_ (.A1(_00654_),
    .A2(_13190_),
    .B1(_14485_),
    .B2(net309),
    .C(_14486_),
    .Y(_14487_));
 AO21x1_ASAP7_75t_R _19796_ (.A1(_13215_),
    .A2(_14483_),
    .B(_14487_),
    .Y(_14488_));
 AO221x2_ASAP7_75t_R _19797_ (.A1(_14452_),
    .A2(_14463_),
    .B1(_14476_),
    .B2(_13614_),
    .C(_14488_),
    .Y(_14489_));
 TIEHIx1_ASAP7_75t_R _34454__466 (.H(net466));
 AND2x2_ASAP7_75t_R _19799_ (.A(net309),
    .B(_14436_),
    .Y(_14491_));
 OR4x2_ASAP7_75t_R _19800_ (.A(_13273_),
    .B(_01746_),
    .C(_13543_),
    .D(_13245_),
    .Y(_14492_));
 OR3x1_ASAP7_75t_R _19801_ (.A(_00323_),
    .B(_13328_),
    .C(_14492_),
    .Y(_14493_));
 OA31x2_ASAP7_75t_R _19802_ (.A1(_00280_),
    .A2(_13288_),
    .A3(_13287_),
    .B1(_14493_),
    .Y(_14494_));
 OR3x2_ASAP7_75t_R _19803_ (.A(_13270_),
    .B(_13248_),
    .C(_13281_),
    .Y(_14495_));
 NOR2x2_ASAP7_75t_R _19804_ (.A(_14494_),
    .B(_14495_),
    .Y(_14496_));
 AOI221x1_ASAP7_75t_R _19805_ (.A1(_13583_),
    .A2(_14489_),
    .B1(_14491_),
    .B2(_13269_),
    .C(_14496_),
    .Y(_14497_));
 TIEHIx1_ASAP7_75t_R _34453__465 (.H(net465));
 INVx4_ASAP7_75t_R _19807_ (.A(_14497_),
    .Y(_18162_));
 INVx1_ASAP7_75t_R _19808_ (.A(_01476_),
    .Y(\cs_registers_i.mhpmcounter[2][12] ));
 INVx1_ASAP7_75t_R _19809_ (.A(_01507_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[12] ));
 TIEHIx1_ASAP7_75t_R _34452__464 (.H(net464));
 AND5x2_ASAP7_75t_R _19811_ (.A(_00290_),
    .B(_00289_),
    .C(net374),
    .D(_00287_),
    .E(_00286_),
    .Y(_14499_));
 AND2x2_ASAP7_75t_R _19812_ (.A(_13323_),
    .B(_14499_),
    .Y(_14500_));
 OR3x4_ASAP7_75t_R _19813_ (.A(_00281_),
    .B(_13547_),
    .C(_14500_),
    .Y(_17594_));
 INVx1_ASAP7_75t_R _19814_ (.A(_17594_),
    .Y(_17598_));
 NOR3x2_ASAP7_75t_R _19815_ (.B(_13547_),
    .C(_14499_),
    .Y(_14501_),
    .A(_00282_));
 CKINVDCx11_ASAP7_75t_R _19816_ (.A(_14501_),
    .Y(_14502_));
 TIEHIx1_ASAP7_75t_R _34451__463 (.H(net463));
 INVx3_ASAP7_75t_R _19818_ (.A(_00196_),
    .Y(\cs_registers_i.pc_id_i[11] ));
 NOR2x2_ASAP7_75t_R _19819_ (.A(_13879_),
    .B(_13561_),
    .Y(_14503_));
 TIEHIx1_ASAP7_75t_R _34450__462 (.H(net462));
 TIEHIx1_ASAP7_75t_R _34449__461 (.H(net461));
 TIEHIx1_ASAP7_75t_R _34448__460 (.H(net460));
 TIEHIx1_ASAP7_75t_R _34447__459 (.H(net459));
 NAND2x1_ASAP7_75t_R _19824_ (.A(net383),
    .B(_00640_),
    .Y(_14508_));
 OA211x2_ASAP7_75t_R _19825_ (.A1(net383),
    .A2(_14467_),
    .B(_14508_),
    .C(net374),
    .Y(_14509_));
 NAND2x1_ASAP7_75t_R _19826_ (.A(net383),
    .B(_00644_),
    .Y(_14510_));
 OA211x2_ASAP7_75t_R _19827_ (.A1(net383),
    .A2(_14470_),
    .B(_14510_),
    .C(_13397_),
    .Y(_14511_));
 OR3x1_ASAP7_75t_R _19828_ (.A(net304),
    .B(_14509_),
    .C(_14511_),
    .Y(_14512_));
 NAND2x1_ASAP7_75t_R _19829_ (.A(net383),
    .B(_00641_),
    .Y(_14513_));
 OA211x2_ASAP7_75t_R _19830_ (.A1(net383),
    .A2(_14464_),
    .B(_14513_),
    .C(net374),
    .Y(_14514_));
 NAND2x1_ASAP7_75t_R _19831_ (.A(net383),
    .B(_00645_),
    .Y(_14515_));
 OA211x2_ASAP7_75t_R _19832_ (.A1(net383),
    .A2(_14473_),
    .B(_14515_),
    .C(_13397_),
    .Y(_14516_));
 OR3x1_ASAP7_75t_R _19833_ (.A(net412),
    .B(_14514_),
    .C(_14516_),
    .Y(_14517_));
 TIEHIx1_ASAP7_75t_R _34446__458 (.H(net458));
 INVx1_ASAP7_75t_R _19835_ (.A(_00631_),
    .Y(_14519_));
 NAND2x1_ASAP7_75t_R _19836_ (.A(net383),
    .B(_00629_),
    .Y(_14520_));
 OA211x2_ASAP7_75t_R _19837_ (.A1(net383),
    .A2(_14519_),
    .B(_14520_),
    .C(net305),
    .Y(_14521_));
 INVx1_ASAP7_75t_R _19838_ (.A(_00630_),
    .Y(_14522_));
 NAND2x1_ASAP7_75t_R _19839_ (.A(net383),
    .B(_00628_),
    .Y(_14523_));
 OA211x2_ASAP7_75t_R _19840_ (.A1(net383),
    .A2(_14522_),
    .B(_14523_),
    .C(net405),
    .Y(_14524_));
 OR3x1_ASAP7_75t_R _19841_ (.A(net298),
    .B(_14521_),
    .C(_14524_),
    .Y(_14525_));
 TIEHIx1_ASAP7_75t_R _34445__457 (.H(net457));
 TIELOx1_ASAP7_75t_R _36363__455 (.L(net455));
 NAND2x1_ASAP7_75t_R _19844_ (.A(net383),
    .B(_01698_),
    .Y(_14528_));
 TIELOx1_ASAP7_75t_R _36362__454 (.L(net454));
 OA211x2_ASAP7_75t_R _19846_ (.A1(net383),
    .A2(_14459_),
    .B(_14528_),
    .C(net304),
    .Y(_14530_));
 AND3x1_ASAP7_75t_R _19847_ (.A(net405),
    .B(net303),
    .C(_14458_),
    .Y(_14531_));
 OA31x2_ASAP7_75t_R _19848_ (.A1(net301),
    .A2(_14530_),
    .A3(_14531_),
    .B1(net363),
    .Y(_14532_));
 AO32x1_ASAP7_75t_R _19849_ (.A1(_13392_),
    .A2(_14512_),
    .A3(_14517_),
    .B1(_14525_),
    .B2(_14532_),
    .Y(_14533_));
 TIELOx1_ASAP7_75t_R _36331__453 (.L(net453));
 TIELOx1_ASAP7_75t_R _36330__452 (.L(net452));
 TIELOx1_ASAP7_75t_R _36329__451 (.L(net451));
 NAND2x1_ASAP7_75t_R _19853_ (.A(net383),
    .B(_00633_),
    .Y(_14537_));
 OA211x2_ASAP7_75t_R _19854_ (.A1(net381),
    .A2(_14449_),
    .B(_14537_),
    .C(net304),
    .Y(_14538_));
 TIELOx1_ASAP7_75t_R ibex_core_450 (.L(net450));
 BUFx16f_ASAP7_75t_R load_slew449 (.A(net148),
    .Y(net449));
 NAND2x1_ASAP7_75t_R _19857_ (.A(net381),
    .B(_00632_),
    .Y(_14541_));
 OA211x2_ASAP7_75t_R _19858_ (.A1(net381),
    .A2(_14442_),
    .B(_14541_),
    .C(net404),
    .Y(_14542_));
 OR3x1_ASAP7_75t_R _19859_ (.A(_13397_),
    .B(_14538_),
    .C(_14542_),
    .Y(_14543_));
 BUFx16f_ASAP7_75t_R load_slew448 (.A(net148),
    .Y(net448));
 NAND2x1_ASAP7_75t_R _19861_ (.A(net381),
    .B(_00637_),
    .Y(_14545_));
 BUFx16f_ASAP7_75t_R load_slew447 (.A(net448),
    .Y(net447));
 OA211x2_ASAP7_75t_R _19863_ (.A1(net381),
    .A2(_14446_),
    .B(_14545_),
    .C(net304),
    .Y(_14547_));
 BUFx16f_ASAP7_75t_R load_slew446 (.A(net447),
    .Y(net446));
 NAND2x1_ASAP7_75t_R _19865_ (.A(net381),
    .B(_00636_),
    .Y(_14549_));
 BUFx16f_ASAP7_75t_R load_slew445 (.A(net447),
    .Y(net445));
 OA211x2_ASAP7_75t_R _19867_ (.A1(net381),
    .A2(_14439_),
    .B(_14549_),
    .C(net404),
    .Y(_14551_));
 OR3x1_ASAP7_75t_R _19868_ (.A(net374),
    .B(_14547_),
    .C(_14551_),
    .Y(_14552_));
 AND2x2_ASAP7_75t_R _19869_ (.A(_14543_),
    .B(_14552_),
    .Y(_14553_));
 AND2x2_ASAP7_75t_R _19870_ (.A(_14525_),
    .B(_14532_),
    .Y(_14554_));
 BUFx16f_ASAP7_75t_R load_slew444 (.A(net445),
    .Y(net444));
 BUFx16f_ASAP7_75t_R load_slew443 (.A(net447),
    .Y(net443));
 BUFx16f_ASAP7_75t_R load_slew442 (.A(net443),
    .Y(net442));
 NOR2x1_ASAP7_75t_R _19874_ (.A(net374),
    .B(_00654_),
    .Y(_14558_));
 AO21x1_ASAP7_75t_R _19875_ (.A1(net374),
    .A2(_14477_),
    .B(_14558_),
    .Y(_14559_));
 INVx1_ASAP7_75t_R _19876_ (.A(_00655_),
    .Y(_14560_));
 NAND2x1_ASAP7_75t_R _19877_ (.A(net373),
    .B(_00651_),
    .Y(_14561_));
 OA211x2_ASAP7_75t_R _19878_ (.A1(net373),
    .A2(_14560_),
    .B(_14561_),
    .C(net305),
    .Y(_14562_));
 AO21x1_ASAP7_75t_R _19879_ (.A1(net411),
    .A2(_14559_),
    .B(_14562_),
    .Y(_14563_));
 BUFx16f_ASAP7_75t_R load_slew441 (.A(net442),
    .Y(net441));
 NAND2x1_ASAP7_75t_R _19881_ (.A(net411),
    .B(_00648_),
    .Y(_14565_));
 OA211x2_ASAP7_75t_R _19882_ (.A1(net411),
    .A2(_14480_),
    .B(_14565_),
    .C(net373),
    .Y(_14566_));
 INVx1_ASAP7_75t_R _19883_ (.A(_00653_),
    .Y(_14567_));
 NAND2x1_ASAP7_75t_R _19884_ (.A(net411),
    .B(_00652_),
    .Y(_14568_));
 OA211x2_ASAP7_75t_R _19885_ (.A1(net411),
    .A2(_14567_),
    .B(_14568_),
    .C(_13397_),
    .Y(_14569_));
 OR3x1_ASAP7_75t_R _19886_ (.A(_13433_),
    .B(_14566_),
    .C(_14569_),
    .Y(_14570_));
 NOR2x2_ASAP7_75t_R _19887_ (.A(net366),
    .B(net363),
    .Y(_14571_));
 BUFx16f_ASAP7_75t_R load_slew440 (.A(net443),
    .Y(net440));
 OA211x2_ASAP7_75t_R _19889_ (.A1(net384),
    .A2(_14563_),
    .B(_14570_),
    .C(_14571_),
    .Y(_14573_));
 AO221x2_ASAP7_75t_R _19890_ (.A1(net367),
    .A2(_14533_),
    .B1(_14553_),
    .B2(_14554_),
    .C(_14573_),
    .Y(_14574_));
 NOR2x1_ASAP7_75t_R _19891_ (.A(_01630_),
    .B(_13223_),
    .Y(_14575_));
 AOI221x1_ASAP7_75t_R _19892_ (.A1(\cs_registers_i.pc_id_i[11] ),
    .A2(_14503_),
    .B1(_14574_),
    .B2(_13563_),
    .C(_14575_),
    .Y(_14576_));
 BUFx16f_ASAP7_75t_R load_slew439 (.A(net440),
    .Y(net439));
 INVx1_ASAP7_75t_R _19894_ (.A(_01487_),
    .Y(\cs_registers_i.mhpmcounter[2][1] ));
 INVx1_ASAP7_75t_R _19895_ (.A(_01518_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[1] ));
 INVx1_ASAP7_75t_R _19896_ (.A(_02066_),
    .Y(\cs_registers_i.mhpmcounter[2][32] ));
 INVx1_ASAP7_75t_R _19897_ (.A(_02172_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[32] ));
 INVx2_ASAP7_75t_R _19898_ (.A(_01732_),
    .Y(_14577_));
 BUFx16f_ASAP7_75t_R load_slew438 (.A(net440),
    .Y(net438));
 BUFx16f_ASAP7_75t_R max_length437 (.A(net449),
    .Y(net437));
 INVx4_ASAP7_75t_R _19901_ (.A(_01717_),
    .Y(_14580_));
 INVx2_ASAP7_75t_R _19902_ (.A(_01715_),
    .Y(_14581_));
 BUFx16f_ASAP7_75t_R load_slew436 (.A(net449),
    .Y(net436));
 AND3x4_ASAP7_75t_R _19904_ (.A(_01714_),
    .B(_14581_),
    .C(_01716_),
    .Y(_14583_));
 AND2x2_ASAP7_75t_R _19905_ (.A(_14580_),
    .B(_14583_),
    .Y(_14584_));
 AND3x4_ASAP7_75t_R _19906_ (.A(_13227_),
    .B(_01721_),
    .C(_14584_),
    .Y(_14585_));
 BUFx16f_ASAP7_75t_R load_slew435 (.A(net449),
    .Y(net435));
 OR2x2_ASAP7_75t_R _19908_ (.A(_13358_),
    .B(_13379_),
    .Y(_14587_));
 AO22x1_ASAP7_75t_R _19909_ (.A1(_00279_),
    .A2(_13369_),
    .B1(_01743_),
    .B2(_13323_),
    .Y(_14588_));
 AND2x2_ASAP7_75t_R _19910_ (.A(_13261_),
    .B(_14588_),
    .Y(_14589_));
 AND3x1_ASAP7_75t_R _19911_ (.A(_01739_),
    .B(_13372_),
    .C(_13335_),
    .Y(_14590_));
 INVx1_ASAP7_75t_R _19912_ (.A(_14590_),
    .Y(_14591_));
 OA211x2_ASAP7_75t_R _19913_ (.A1(_14587_),
    .A2(_14589_),
    .B(_14591_),
    .C(_13317_),
    .Y(_14592_));
 NAND2x1_ASAP7_75t_R _19914_ (.A(_00281_),
    .B(_00282_),
    .Y(_14593_));
 NOR2x1_ASAP7_75t_R _19915_ (.A(_13547_),
    .B(_14593_),
    .Y(_14594_));
 AND4x2_ASAP7_75t_R _19916_ (.A(net316),
    .B(_01739_),
    .C(_01742_),
    .D(_01743_),
    .Y(_14595_));
 NAND3x2_ASAP7_75t_R _19917_ (.B(_00283_),
    .C(_14595_),
    .Y(_14596_),
    .A(_00280_));
 INVx1_ASAP7_75t_R _19918_ (.A(_00280_),
    .Y(_14597_));
 OR3x1_ASAP7_75t_R _19919_ (.A(net316),
    .B(_01739_),
    .C(_01743_),
    .Y(_14598_));
 OR4x2_ASAP7_75t_R _19920_ (.A(_14597_),
    .B(_14141_),
    .C(_01742_),
    .D(_14598_),
    .Y(_14599_));
 OR5x2_ASAP7_75t_R _19921_ (.A(net309),
    .B(_01745_),
    .C(_01740_),
    .D(_01741_),
    .E(_13584_),
    .Y(_14600_));
 AO21x2_ASAP7_75t_R _19922_ (.A1(_14596_),
    .A2(_14599_),
    .B(_14600_),
    .Y(_14601_));
 OR3x1_ASAP7_75t_R _19923_ (.A(net360),
    .B(_01744_),
    .C(_01741_),
    .Y(_14602_));
 OA21x2_ASAP7_75t_R _19924_ (.A1(_13132_),
    .A2(_14318_),
    .B(_14602_),
    .Y(_14603_));
 OR5x1_ASAP7_75t_R _19925_ (.A(_13127_),
    .B(_13598_),
    .C(_14375_),
    .D(_14596_),
    .E(_14603_),
    .Y(_14604_));
 OR4x1_ASAP7_75t_R _19926_ (.A(_00172_),
    .B(_13245_),
    .C(_13546_),
    .D(_14593_),
    .Y(_14605_));
 AND4x1_ASAP7_75t_R _19927_ (.A(_00323_),
    .B(_00184_),
    .C(_00187_),
    .D(_00191_),
    .Y(_14606_));
 AND4x1_ASAP7_75t_R _19928_ (.A(_00279_),
    .B(_00194_),
    .C(_14499_),
    .D(_14606_),
    .Y(_14607_));
 OAI21x1_ASAP7_75t_R _19929_ (.A1(_14605_),
    .A2(_14607_),
    .B(_01847_),
    .Y(_14608_));
 AO31x2_ASAP7_75t_R _19930_ (.A1(_14594_),
    .A2(_14601_),
    .A3(_14604_),
    .B(_14608_),
    .Y(_14609_));
 AND2x2_ASAP7_75t_R _19931_ (.A(_00165_),
    .B(_13238_),
    .Y(_14610_));
 OA21x2_ASAP7_75t_R _19932_ (.A1(_00165_),
    .A2(_13273_),
    .B(_00278_),
    .Y(_14611_));
 OA21x2_ASAP7_75t_R _19933_ (.A1(_14610_),
    .A2(_14611_),
    .B(_00168_),
    .Y(_14612_));
 AND3x1_ASAP7_75t_R _19934_ (.A(_13271_),
    .B(_00172_),
    .C(_13347_),
    .Y(_14613_));
 OA21x2_ASAP7_75t_R _19935_ (.A1(_13323_),
    .A2(_13238_),
    .B(_13325_),
    .Y(_14614_));
 AND5x2_ASAP7_75t_R _19936_ (.A(_00278_),
    .B(_13272_),
    .C(_00172_),
    .D(_13230_),
    .E(_13252_),
    .Y(_14615_));
 OAI21x1_ASAP7_75t_R _19937_ (.A1(_13335_),
    .A2(_14614_),
    .B(_14615_),
    .Y(_14616_));
 OAI21x1_ASAP7_75t_R _19938_ (.A1(_14612_),
    .A2(_14613_),
    .B(_14616_),
    .Y(_14617_));
 AND2x2_ASAP7_75t_R _19939_ (.A(_13271_),
    .B(_13352_),
    .Y(_14618_));
 OAI21x1_ASAP7_75t_R _19940_ (.A1(_13381_),
    .A2(_14618_),
    .B(_13280_),
    .Y(_14619_));
 NAND3x1_ASAP7_75t_R _19941_ (.A(_13259_),
    .B(_13345_),
    .C(_14619_),
    .Y(_14620_));
 OR4x1_ASAP7_75t_R _19942_ (.A(_13255_),
    .B(_00163_),
    .C(_00172_),
    .D(_01746_),
    .Y(_14621_));
 OR4x1_ASAP7_75t_R _19943_ (.A(_13245_),
    .B(_13350_),
    .C(_14621_),
    .D(_13338_),
    .Y(_14622_));
 NOR2x1_ASAP7_75t_R _19944_ (.A(_13238_),
    .B(_14622_),
    .Y(_14623_));
 OR4x2_ASAP7_75t_R _19945_ (.A(_14609_),
    .B(_14617_),
    .C(_14620_),
    .D(_14623_),
    .Y(_14624_));
 NOR2x2_ASAP7_75t_R _19946_ (.A(_14592_),
    .B(_14624_),
    .Y(_14625_));
 AND3x4_ASAP7_75t_R _19947_ (.A(_13576_),
    .B(_14585_),
    .C(_14625_),
    .Y(_14626_));
 BUFx16f_ASAP7_75t_R load_slew434 (.A(net435),
    .Y(net434));
 NAND2x2_ASAP7_75t_R _19949_ (.A(_00279_),
    .B(_14626_),
    .Y(_14628_));
 BUFx16f_ASAP7_75t_R wire433 (.A(net435),
    .Y(net433));
 BUFx16f_ASAP7_75t_R wire432 (.A(net433),
    .Y(net432));
 AO21x1_ASAP7_75t_R _19952_ (.A1(_13313_),
    .A2(_13550_),
    .B(_01874_),
    .Y(_14631_));
 AOI211x1_ASAP7_75t_R _19953_ (.A1(_01314_),
    .A2(_14631_),
    .B(_14628_),
    .C(_14141_),
    .Y(_14632_));
 AO21x1_ASAP7_75t_R _19954_ (.A1(_14577_),
    .A2(_14628_),
    .B(_14632_),
    .Y(_00000_));
 INVx2_ASAP7_75t_R _19955_ (.A(_00162_),
    .Y(\cs_registers_i.pc_id_i[2] ));
 NAND2x1_ASAP7_75t_R _19956_ (.A(net401),
    .B(_00374_),
    .Y(_14633_));
 OA211x2_ASAP7_75t_R _19957_ (.A1(net401),
    .A2(_13887_),
    .B(_14633_),
    .C(net307),
    .Y(_14634_));
 BUFx16f_ASAP7_75t_R load_slew431 (.A(net432),
    .Y(net431));
 NAND2x1_ASAP7_75t_R _19959_ (.A(net401),
    .B(_00373_),
    .Y(_14636_));
 OA211x2_ASAP7_75t_R _19960_ (.A1(net401),
    .A2(_13883_),
    .B(_14636_),
    .C(net411),
    .Y(_14637_));
 OR3x1_ASAP7_75t_R _19961_ (.A(net373),
    .B(_14634_),
    .C(_14637_),
    .Y(_14638_));
 NAND2x1_ASAP7_75t_R _19962_ (.A(net401),
    .B(_00370_),
    .Y(_14639_));
 OA211x2_ASAP7_75t_R _19963_ (.A1(net401),
    .A2(_13890_),
    .B(_14639_),
    .C(net307),
    .Y(_14640_));
 NAND2x1_ASAP7_75t_R _19964_ (.A(net401),
    .B(_00369_),
    .Y(_14641_));
 OA211x2_ASAP7_75t_R _19965_ (.A1(net401),
    .A2(_13893_),
    .B(_14641_),
    .C(net411),
    .Y(_14642_));
 OR3x1_ASAP7_75t_R _19966_ (.A(_13397_),
    .B(_14640_),
    .C(_14642_),
    .Y(_14643_));
 INVx1_ASAP7_75t_R _19967_ (.A(_00360_),
    .Y(_14644_));
 NAND2x1_ASAP7_75t_R _19968_ (.A(net401),
    .B(_00358_),
    .Y(_14645_));
 OA211x2_ASAP7_75t_R _19969_ (.A1(net401),
    .A2(_14644_),
    .B(_14645_),
    .C(net307),
    .Y(_14646_));
 INVx1_ASAP7_75t_R _19970_ (.A(_00359_),
    .Y(_14647_));
 NAND2x1_ASAP7_75t_R _19971_ (.A(net400),
    .B(_00357_),
    .Y(_14648_));
 OA211x2_ASAP7_75t_R _19972_ (.A1(net400),
    .A2(_14647_),
    .B(_14648_),
    .C(net411),
    .Y(_14649_));
 OR3x1_ASAP7_75t_R _19973_ (.A(net298),
    .B(_14646_),
    .C(_14649_),
    .Y(_14650_));
 INVx1_ASAP7_75t_R _19974_ (.A(_00356_),
    .Y(_14651_));
 NAND2x1_ASAP7_75t_R _19975_ (.A(net411),
    .B(_00355_),
    .Y(_14652_));
 OA211x2_ASAP7_75t_R _19976_ (.A1(net411),
    .A2(_14651_),
    .B(_14652_),
    .C(net302),
    .Y(_14653_));
 AND3x1_ASAP7_75t_R _19977_ (.A(net307),
    .B(net401),
    .C(_13918_),
    .Y(_14654_));
 OA31x2_ASAP7_75t_R _19978_ (.A1(net300),
    .A2(_14653_),
    .A3(_14654_),
    .B1(net362),
    .Y(_14655_));
 AO32x1_ASAP7_75t_R _19979_ (.A1(_13392_),
    .A2(_14638_),
    .A3(_14643_),
    .B1(_14650_),
    .B2(_14655_),
    .Y(_14656_));
 NAND2x1_ASAP7_75t_R _19980_ (.A(net383),
    .B(_00366_),
    .Y(_14657_));
 OA211x2_ASAP7_75t_R _19981_ (.A1(net383),
    .A2(_13903_),
    .B(_14657_),
    .C(net305),
    .Y(_14658_));
 NAND2x1_ASAP7_75t_R _19982_ (.A(net383),
    .B(_00365_),
    .Y(_14659_));
 OA211x2_ASAP7_75t_R _19983_ (.A1(net383),
    .A2(_13900_),
    .B(_14659_),
    .C(net411),
    .Y(_14660_));
 OR3x1_ASAP7_75t_R _19984_ (.A(net373),
    .B(_14658_),
    .C(_14660_),
    .Y(_14661_));
 NAND2x1_ASAP7_75t_R _19985_ (.A(net383),
    .B(_00362_),
    .Y(_14662_));
 OA211x2_ASAP7_75t_R _19986_ (.A1(net383),
    .A2(_13908_),
    .B(_14662_),
    .C(net305),
    .Y(_14663_));
 NAND2x1_ASAP7_75t_R _19987_ (.A(net401),
    .B(_00361_),
    .Y(_14664_));
 OA211x2_ASAP7_75t_R _19988_ (.A1(net401),
    .A2(_13897_),
    .B(_14664_),
    .C(net411),
    .Y(_14665_));
 OR3x1_ASAP7_75t_R _19989_ (.A(_13397_),
    .B(_14663_),
    .C(_14665_),
    .Y(_14666_));
 AND2x2_ASAP7_75t_R _19990_ (.A(_14661_),
    .B(_14666_),
    .Y(_14667_));
 AND2x2_ASAP7_75t_R _19991_ (.A(_14650_),
    .B(_14655_),
    .Y(_14668_));
 BUFx16f_ASAP7_75t_R load_slew430 (.A(net433),
    .Y(net430));
 BUFx16f_ASAP7_75t_R load_slew429 (.A(net430),
    .Y(net429));
 BUFx16f_ASAP7_75t_R load_slew428 (.A(net429),
    .Y(net428));
 NOR2x1_ASAP7_75t_R _19995_ (.A(net383),
    .B(_00383_),
    .Y(_14672_));
 AO21x1_ASAP7_75t_R _19996_ (.A1(net383),
    .A2(_13925_),
    .B(_14672_),
    .Y(_14673_));
 NAND2x1_ASAP7_75t_R _19997_ (.A(net383),
    .B(_00382_),
    .Y(_14674_));
 OA211x2_ASAP7_75t_R _19998_ (.A1(net383),
    .A2(_13929_),
    .B(_14674_),
    .C(net305),
    .Y(_14675_));
 AO21x1_ASAP7_75t_R _19999_ (.A1(net411),
    .A2(_14673_),
    .B(_14675_),
    .Y(_14676_));
 INVx1_ASAP7_75t_R _20000_ (.A(_00380_),
    .Y(_14677_));
 NAND2x1_ASAP7_75t_R _20001_ (.A(net384),
    .B(_00378_),
    .Y(_14678_));
 OA211x2_ASAP7_75t_R _20002_ (.A1(net384),
    .A2(_14677_),
    .B(_14678_),
    .C(net305),
    .Y(_14679_));
 NAND2x1_ASAP7_75t_R _20003_ (.A(net384),
    .B(_00377_),
    .Y(_14680_));
 OA211x2_ASAP7_75t_R _20004_ (.A1(net384),
    .A2(_13937_),
    .B(_14680_),
    .C(net411),
    .Y(_14681_));
 OR3x1_ASAP7_75t_R _20005_ (.A(_13397_),
    .B(_14679_),
    .C(_14681_),
    .Y(_14682_));
 OA211x2_ASAP7_75t_R _20006_ (.A1(net373),
    .A2(_14676_),
    .B(_14682_),
    .C(_14571_),
    .Y(_14683_));
 AO221x2_ASAP7_75t_R _20007_ (.A1(net367),
    .A2(_14656_),
    .B1(_14667_),
    .B2(_14668_),
    .C(_14683_),
    .Y(_14684_));
 BUFx16f_ASAP7_75t_R load_slew427 (.A(net428),
    .Y(net427));
 NAND2x2_ASAP7_75t_R _20009_ (.A(_13223_),
    .B(_13551_),
    .Y(_14686_));
 OAI22x1_ASAP7_75t_R _20010_ (.A1(_01639_),
    .A2(_13223_),
    .B1(_14686_),
    .B2(net374),
    .Y(_14687_));
 AOI221x1_ASAP7_75t_R _20011_ (.A1(\cs_registers_i.pc_id_i[2] ),
    .A2(_14503_),
    .B1(_14684_),
    .B2(_13563_),
    .C(_14687_),
    .Y(_14688_));
 BUFx16f_ASAP7_75t_R load_slew426 (.A(net428),
    .Y(net426));
 XNOR2x1_ASAP7_75t_R _20013_ (.B(_14026_),
    .Y(_14689_),
    .A(_13387_));
 BUFx16f_ASAP7_75t_R load_slew425 (.A(net429),
    .Y(net425));
 NAND2x1_ASAP7_75t_R _20015_ (.A(net382),
    .B(_00409_),
    .Y(_14691_));
 OA211x2_ASAP7_75t_R _20016_ (.A1(net382),
    .A2(_13972_),
    .B(_14691_),
    .C(net305),
    .Y(_14692_));
 BUFx16f_ASAP7_75t_R load_slew424 (.A(net429),
    .Y(net424));
 INVx1_ASAP7_75t_R _20018_ (.A(_00410_),
    .Y(_14694_));
 NAND2x1_ASAP7_75t_R _20019_ (.A(net386),
    .B(_00408_),
    .Y(_14695_));
 BUFx16f_ASAP7_75t_R load_slew423 (.A(net424),
    .Y(net423));
 OA211x2_ASAP7_75t_R _20021_ (.A1(net386),
    .A2(_14694_),
    .B(_14695_),
    .C(net404),
    .Y(_14697_));
 OR3x1_ASAP7_75t_R _20022_ (.A(_13397_),
    .B(_14692_),
    .C(_14697_),
    .Y(_14698_));
 NAND2x1_ASAP7_75t_R _20023_ (.A(net382),
    .B(_00413_),
    .Y(_14699_));
 OA211x2_ASAP7_75t_R _20024_ (.A1(net382),
    .A2(_13968_),
    .B(_14699_),
    .C(net305),
    .Y(_14700_));
 BUFx16f_ASAP7_75t_R load_slew422 (.A(net425),
    .Y(net422));
 INVx1_ASAP7_75t_R _20026_ (.A(_00414_),
    .Y(_14702_));
 BUFx16f_ASAP7_75t_R max_cap421 (.A(_01722_),
    .Y(net421));
 NAND2x1_ASAP7_75t_R _20028_ (.A(net382),
    .B(_00412_),
    .Y(_14704_));
 OA211x2_ASAP7_75t_R _20029_ (.A1(net382),
    .A2(_14702_),
    .B(_14704_),
    .C(net404),
    .Y(_14705_));
 OR3x1_ASAP7_75t_R _20030_ (.A(net369),
    .B(_14700_),
    .C(_14705_),
    .Y(_14706_));
 AO21x1_ASAP7_75t_R _20031_ (.A1(_14698_),
    .A2(_14706_),
    .B(net368),
    .Y(_14707_));
 BUFx16f_ASAP7_75t_R load_slew420 (.A(_01643_),
    .Y(net420));
 BUFx16f_ASAP7_75t_R max_cap419 (.A(net420),
    .Y(net419));
 NAND2x1_ASAP7_75t_R _20034_ (.A(net386),
    .B(_00401_),
    .Y(_14710_));
 OA211x2_ASAP7_75t_R _20035_ (.A1(net386),
    .A2(_13993_),
    .B(_14710_),
    .C(net305),
    .Y(_14711_));
 NAND2x1_ASAP7_75t_R _20036_ (.A(net386),
    .B(_00400_),
    .Y(_14712_));
 OA21x2_ASAP7_75t_R _20037_ (.A1(net386),
    .A2(_13996_),
    .B(_14712_),
    .Y(_14713_));
 AO21x1_ASAP7_75t_R _20038_ (.A1(net405),
    .A2(_14713_),
    .B(net301),
    .Y(_14714_));
 INVx1_ASAP7_75t_R _20039_ (.A(_00407_),
    .Y(_14715_));
 BUFx16f_ASAP7_75t_R max_cap418 (.A(_01642_),
    .Y(net418));
 NAND2x1_ASAP7_75t_R _20041_ (.A(net385),
    .B(_00405_),
    .Y(_14717_));
 BUFx16f_ASAP7_75t_R load_slew417 (.A(_00662_),
    .Y(net417));
 OA211x2_ASAP7_75t_R _20043_ (.A1(net385),
    .A2(_14715_),
    .B(_14717_),
    .C(net305),
    .Y(_14719_));
 INVx1_ASAP7_75t_R _20044_ (.A(_00406_),
    .Y(_14720_));
 BUFx16f_ASAP7_75t_R max_cap416 (.A(net417),
    .Y(net416));
 NAND2x1_ASAP7_75t_R _20046_ (.A(net385),
    .B(_00404_),
    .Y(_14722_));
 OA211x2_ASAP7_75t_R _20047_ (.A1(net385),
    .A2(_14720_),
    .B(_14722_),
    .C(net405),
    .Y(_14723_));
 OR3x1_ASAP7_75t_R _20048_ (.A(net298),
    .B(_14719_),
    .C(_14723_),
    .Y(_14724_));
 OA21x2_ASAP7_75t_R _20049_ (.A1(_14711_),
    .A2(_14714_),
    .B(_14724_),
    .Y(_14725_));
 INVx1_ASAP7_75t_R _20050_ (.A(_00391_),
    .Y(_14726_));
 NAND2x1_ASAP7_75t_R _20051_ (.A(net386),
    .B(_00389_),
    .Y(_14727_));
 OA211x2_ASAP7_75t_R _20052_ (.A1(net386),
    .A2(_14726_),
    .B(_14727_),
    .C(net305),
    .Y(_14728_));
 INVx1_ASAP7_75t_R _20053_ (.A(_00390_),
    .Y(_14729_));
 NAND2x1_ASAP7_75t_R _20054_ (.A(net386),
    .B(_00388_),
    .Y(_14730_));
 OA211x2_ASAP7_75t_R _20055_ (.A1(net386),
    .A2(_14729_),
    .B(_14730_),
    .C(net405),
    .Y(_14731_));
 OR3x1_ASAP7_75t_R _20056_ (.A(_13484_),
    .B(_14728_),
    .C(_14731_),
    .Y(_14732_));
 NAND2x1_ASAP7_75t_R _20057_ (.A(net382),
    .B(_00397_),
    .Y(_14733_));
 OA211x2_ASAP7_75t_R _20058_ (.A1(net382),
    .A2(_14006_),
    .B(_14733_),
    .C(net305),
    .Y(_14734_));
 NAND2x1_ASAP7_75t_R _20059_ (.A(net382),
    .B(_00396_),
    .Y(_14735_));
 OA211x2_ASAP7_75t_R _20060_ (.A1(net382),
    .A2(_14015_),
    .B(_14735_),
    .C(net404),
    .Y(_14736_));
 OR3x1_ASAP7_75t_R _20061_ (.A(net368),
    .B(_14734_),
    .C(_14736_),
    .Y(_14737_));
 BUFx16f_ASAP7_75t_R load_slew415 (.A(_00237_),
    .Y(net415));
 AO21x1_ASAP7_75t_R _20063_ (.A1(_14732_),
    .A2(_14737_),
    .B(net369),
    .Y(_14739_));
 AND2x2_ASAP7_75t_R _20064_ (.A(net386),
    .B(_01706_),
    .Y(_14740_));
 AO21x1_ASAP7_75t_R _20065_ (.A1(net303),
    .A2(_00387_),
    .B(_14740_),
    .Y(_14741_));
 OAI22x1_ASAP7_75t_R _20066_ (.A1(_00386_),
    .A2(_13471_),
    .B1(_14741_),
    .B2(net405),
    .Y(_14742_));
 NAND2x2_ASAP7_75t_R _20067_ (.A(net373),
    .B(_13484_),
    .Y(_14743_));
 INVx1_ASAP7_75t_R _20068_ (.A(_00395_),
    .Y(_14744_));
 NAND2x1_ASAP7_75t_R _20069_ (.A(net386),
    .B(_00393_),
    .Y(_14745_));
 OA211x2_ASAP7_75t_R _20070_ (.A1(net386),
    .A2(_14744_),
    .B(_14745_),
    .C(net305),
    .Y(_14746_));
 INVx1_ASAP7_75t_R _20071_ (.A(_00394_),
    .Y(_14747_));
 NAND2x1_ASAP7_75t_R _20072_ (.A(net386),
    .B(_00392_),
    .Y(_14748_));
 OA211x2_ASAP7_75t_R _20073_ (.A1(net386),
    .A2(_14747_),
    .B(_14748_),
    .C(net405),
    .Y(_14749_));
 OR3x1_ASAP7_75t_R _20074_ (.A(_14743_),
    .B(_14746_),
    .C(_14749_),
    .Y(_14750_));
 OA211x2_ASAP7_75t_R _20075_ (.A1(net301),
    .A2(_14742_),
    .B(_14750_),
    .C(net363),
    .Y(_14751_));
 AO32x2_ASAP7_75t_R _20076_ (.A1(_13392_),
    .A2(_14707_),
    .A3(_14725_),
    .B1(_14739_),
    .B2(_14751_),
    .Y(_14752_));
 BUFx16f_ASAP7_75t_R load_slew414 (.A(_00240_),
    .Y(net414));
 AOI22x1_ASAP7_75t_R _20078_ (.A1(_13530_),
    .A2(_00665_),
    .B1(_01449_),
    .B2(_13533_),
    .Y(_14754_));
 OA211x2_ASAP7_75t_R _20079_ (.A1(_00284_),
    .A2(_14752_),
    .B(_14754_),
    .C(_13763_),
    .Y(_14755_));
 AOI211x1_ASAP7_75t_R _20080_ (.A1(_13528_),
    .A2(_14019_),
    .B(_14755_),
    .C(net295),
    .Y(_14756_));
 AO21x1_ASAP7_75t_R _20081_ (.A1(net294),
    .A2(_14689_),
    .B(_14756_),
    .Y(_17542_));
 INVx1_ASAP7_75t_R _20082_ (.A(_17542_),
    .Y(_16505_));
 INVx2_ASAP7_75t_R _20083_ (.A(_00170_),
    .Y(\cs_registers_i.pc_id_i[3] ));
 INVx1_ASAP7_75t_R _20084_ (.A(_13561_),
    .Y(_14757_));
 AND2x2_ASAP7_75t_R _20085_ (.A(\cs_registers_i.pc_id_i[3] ),
    .B(_13553_),
    .Y(_14758_));
 AO21x1_ASAP7_75t_R _20086_ (.A1(_13879_),
    .A2(_14752_),
    .B(_14758_),
    .Y(_14759_));
 OAI22x1_ASAP7_75t_R _20087_ (.A1(_01638_),
    .A2(_13223_),
    .B1(_14686_),
    .B2(_00287_),
    .Y(_14760_));
 AO21x2_ASAP7_75t_R _20088_ (.A1(_14757_),
    .A2(_14759_),
    .B(_14760_),
    .Y(_14761_));
 BUFx16f_ASAP7_75t_R max_cap413 (.A(_01815_),
    .Y(net413));
 INVx1_ASAP7_75t_R _20090_ (.A(_14761_),
    .Y(_18121_));
 OAI21x1_ASAP7_75t_R _20091_ (.A1(_00665_),
    .A2(_13574_),
    .B(_13576_),
    .Y(_14762_));
 OA21x2_ASAP7_75t_R _20092_ (.A1(_13576_),
    .A2(_14761_),
    .B(_14762_),
    .Y(_17543_));
 INVx1_ASAP7_75t_R _20093_ (.A(_17543_),
    .Y(_16506_));
 INVx1_ASAP7_75t_R _20094_ (.A(_17539_),
    .Y(_16496_));
 OA21x2_ASAP7_75t_R _20095_ (.A1(_00292_),
    .A2(_16496_),
    .B(_00664_),
    .Y(_14763_));
 OA21x2_ASAP7_75t_R _20096_ (.A1(_02262_),
    .A2(_14763_),
    .B(_00667_),
    .Y(_16504_));
 INVx1_ASAP7_75t_R _20097_ (.A(_00174_),
    .Y(_14764_));
 BUFx16f_ASAP7_75t_R max_cap412 (.A(_00290_),
    .Y(net412));
 NAND2x1_ASAP7_75t_R _20099_ (.A(net376),
    .B(_00435_),
    .Y(_14766_));
 BUFx16f_ASAP7_75t_R load_slew411 (.A(_00290_),
    .Y(net411));
 OA211x2_ASAP7_75t_R _20101_ (.A1(net376),
    .A2(_14069_),
    .B(_14766_),
    .C(net304),
    .Y(_14768_));
 NAND2x1_ASAP7_75t_R _20102_ (.A(net376),
    .B(_00434_),
    .Y(_14769_));
 OA211x2_ASAP7_75t_R _20103_ (.A1(net376),
    .A2(_14066_),
    .B(_14769_),
    .C(net406),
    .Y(_14770_));
 OR3x1_ASAP7_75t_R _20104_ (.A(net375),
    .B(_14768_),
    .C(_14770_),
    .Y(_14771_));
 BUFx16f_ASAP7_75t_R load_slew410 (.A(_00290_),
    .Y(net410));
 NAND2x1_ASAP7_75t_R _20106_ (.A(net376),
    .B(_00431_),
    .Y(_14773_));
 OA211x2_ASAP7_75t_R _20107_ (.A1(net376),
    .A2(_14072_),
    .B(_14773_),
    .C(net304),
    .Y(_14774_));
 NAND2x1_ASAP7_75t_R _20108_ (.A(net376),
    .B(_00430_),
    .Y(_14775_));
 OA211x2_ASAP7_75t_R _20109_ (.A1(net376),
    .A2(_14075_),
    .B(_14775_),
    .C(net406),
    .Y(_14776_));
 OR3x1_ASAP7_75t_R _20110_ (.A(_13397_),
    .B(_14774_),
    .C(_14776_),
    .Y(_14777_));
 BUFx16f_ASAP7_75t_R max_cap409 (.A(net410),
    .Y(net409));
 INVx1_ASAP7_75t_R _20112_ (.A(_00420_),
    .Y(_14779_));
 NAND2x1_ASAP7_75t_R _20113_ (.A(net377),
    .B(_00418_),
    .Y(_14780_));
 OA211x2_ASAP7_75t_R _20114_ (.A1(net377),
    .A2(_14779_),
    .B(_14780_),
    .C(net412),
    .Y(_14781_));
 INVx1_ASAP7_75t_R _20115_ (.A(_00421_),
    .Y(_14782_));
 NAND2x1_ASAP7_75t_R _20116_ (.A(net377),
    .B(_00419_),
    .Y(_14783_));
 OA211x2_ASAP7_75t_R _20117_ (.A1(net377),
    .A2(_14782_),
    .B(_14783_),
    .C(net304),
    .Y(_14784_));
 OR3x1_ASAP7_75t_R _20118_ (.A(net298),
    .B(_14781_),
    .C(_14784_),
    .Y(_14785_));
 NAND2x1_ASAP7_75t_R _20119_ (.A(net376),
    .B(_01705_),
    .Y(_14786_));
 OA211x2_ASAP7_75t_R _20120_ (.A1(net376),
    .A2(_14061_),
    .B(_14786_),
    .C(net304),
    .Y(_14787_));
 AND3x1_ASAP7_75t_R _20121_ (.A(net406),
    .B(_13433_),
    .C(_14060_),
    .Y(_14788_));
 OA31x2_ASAP7_75t_R _20122_ (.A1(net301),
    .A2(_14787_),
    .A3(_14788_),
    .B1(_00286_),
    .Y(_14789_));
 AO32x1_ASAP7_75t_R _20123_ (.A1(_13392_),
    .A2(_14771_),
    .A3(_14777_),
    .B1(_14785_),
    .B2(_14789_),
    .Y(_14790_));
 OR2x2_ASAP7_75t_R _20124_ (.A(net377),
    .B(_00424_),
    .Y(_14791_));
 OAI21x1_ASAP7_75t_R _20125_ (.A1(_13433_),
    .A2(_00422_),
    .B(_14791_),
    .Y(_14792_));
 BUFx12f_ASAP7_75t_R load_slew408 (.A(net410),
    .Y(net408));
 INVx1_ASAP7_75t_R _20127_ (.A(_00425_),
    .Y(_14794_));
 BUFx16f_ASAP7_75t_R load_slew407 (.A(net409),
    .Y(net407));
 NAND2x1_ASAP7_75t_R _20129_ (.A(net377),
    .B(_00423_),
    .Y(_14796_));
 BUFx16f_ASAP7_75t_R load_slew406 (.A(net412),
    .Y(net406));
 OA211x2_ASAP7_75t_R _20131_ (.A1(net377),
    .A2(_14794_),
    .B(_14796_),
    .C(net304),
    .Y(_14798_));
 AO21x1_ASAP7_75t_R _20132_ (.A1(net412),
    .A2(_14792_),
    .B(_14798_),
    .Y(_14799_));
 NAND2x1_ASAP7_75t_R _20133_ (.A(net377),
    .B(_00427_),
    .Y(_14800_));
 OA211x2_ASAP7_75t_R _20134_ (.A1(net377),
    .A2(_14051_),
    .B(_14800_),
    .C(net304),
    .Y(_14801_));
 NAND2x1_ASAP7_75t_R _20135_ (.A(net377),
    .B(_00426_),
    .Y(_14802_));
 BUFx16f_ASAP7_75t_R max_cap405 (.A(net412),
    .Y(net405));
 OA211x2_ASAP7_75t_R _20137_ (.A1(net377),
    .A2(_14042_),
    .B(_14802_),
    .C(net412),
    .Y(_14804_));
 OA21x2_ASAP7_75t_R _20138_ (.A1(_14801_),
    .A2(_14804_),
    .B(_13397_),
    .Y(_14805_));
 AO21x1_ASAP7_75t_R _20139_ (.A1(net375),
    .A2(_14799_),
    .B(_14805_),
    .Y(_14806_));
 AND2x2_ASAP7_75t_R _20140_ (.A(_14785_),
    .B(_14789_),
    .Y(_14807_));
 INVx1_ASAP7_75t_R _20141_ (.A(_00441_),
    .Y(_14808_));
 NAND2x1_ASAP7_75t_R _20142_ (.A(net376),
    .B(_00439_),
    .Y(_14809_));
 OA211x2_ASAP7_75t_R _20143_ (.A1(net376),
    .A2(_14808_),
    .B(_14809_),
    .C(net304),
    .Y(_14810_));
 NAND2x1_ASAP7_75t_R _20144_ (.A(net376),
    .B(_00438_),
    .Y(_14811_));
 OA211x2_ASAP7_75t_R _20145_ (.A1(net376),
    .A2(_14029_),
    .B(_14811_),
    .C(net406),
    .Y(_14812_));
 OR3x1_ASAP7_75t_R _20146_ (.A(_13397_),
    .B(_14810_),
    .C(_14812_),
    .Y(_14813_));
 NAND2x1_ASAP7_75t_R _20147_ (.A(net376),
    .B(_00443_),
    .Y(_14814_));
 OA211x2_ASAP7_75t_R _20148_ (.A1(net376),
    .A2(_14038_),
    .B(_14814_),
    .C(net304),
    .Y(_14815_));
 NAND2x1_ASAP7_75t_R _20149_ (.A(net376),
    .B(_00442_),
    .Y(_14816_));
 OA211x2_ASAP7_75t_R _20150_ (.A1(net376),
    .A2(_14035_),
    .B(_14816_),
    .C(net406),
    .Y(_14817_));
 OR3x1_ASAP7_75t_R _20151_ (.A(net375),
    .B(_14815_),
    .C(_14817_),
    .Y(_14818_));
 AND3x1_ASAP7_75t_R _20152_ (.A(_14571_),
    .B(_14813_),
    .C(_14818_),
    .Y(_14819_));
 AO221x2_ASAP7_75t_R _20153_ (.A1(net368),
    .A2(_14790_),
    .B1(_14806_),
    .B2(_14807_),
    .C(_14819_),
    .Y(_14820_));
 OAI22x1_ASAP7_75t_R _20154_ (.A1(_01637_),
    .A2(_13223_),
    .B1(_14686_),
    .B2(_00286_),
    .Y(_14821_));
 AOI221x1_ASAP7_75t_R _20155_ (.A1(_14764_),
    .A2(_14503_),
    .B1(_14820_),
    .B2(_13563_),
    .C(_14821_),
    .Y(_14822_));
 BUFx16f_ASAP7_75t_R max_cap404 (.A(net412),
    .Y(net404));
 XNOR2x1_ASAP7_75t_R _20157_ (.B(_14140_),
    .Y(_14823_),
    .A(_13387_));
 NAND2x1_ASAP7_75t_R _20158_ (.A(net401),
    .B(_00465_),
    .Y(_14824_));
 OA211x2_ASAP7_75t_R _20159_ (.A1(net401),
    .A2(_14094_),
    .B(_14824_),
    .C(net307),
    .Y(_14825_));
 NAND2x1_ASAP7_75t_R _20160_ (.A(net401),
    .B(_00464_),
    .Y(_14826_));
 OA211x2_ASAP7_75t_R _20161_ (.A1(net401),
    .A2(_14091_),
    .B(_14826_),
    .C(net411),
    .Y(_14827_));
 OR3x1_ASAP7_75t_R _20162_ (.A(net373),
    .B(_14825_),
    .C(_14827_),
    .Y(_14828_));
 BUFx12f_ASAP7_75t_R load_slew403 (.A(_00289_),
    .Y(net403));
 NAND2x1_ASAP7_75t_R _20164_ (.A(net401),
    .B(_00461_),
    .Y(_14830_));
 OA211x2_ASAP7_75t_R _20165_ (.A1(net401),
    .A2(_14085_),
    .B(_14830_),
    .C(net307),
    .Y(_14831_));
 NAND2x1_ASAP7_75t_R _20166_ (.A(net401),
    .B(_00460_),
    .Y(_14832_));
 OA211x2_ASAP7_75t_R _20167_ (.A1(net401),
    .A2(_14088_),
    .B(_14832_),
    .C(net411),
    .Y(_14833_));
 OR3x1_ASAP7_75t_R _20168_ (.A(_13397_),
    .B(_14831_),
    .C(_14833_),
    .Y(_14834_));
 BUFx16f_ASAP7_75t_R load_slew402 (.A(_00289_),
    .Y(net402));
 INVx1_ASAP7_75t_R _20170_ (.A(_00451_),
    .Y(_14836_));
 NAND2x1_ASAP7_75t_R _20171_ (.A(net386),
    .B(_00449_),
    .Y(_14837_));
 OA211x2_ASAP7_75t_R _20172_ (.A1(net386),
    .A2(_14836_),
    .B(_14837_),
    .C(net305),
    .Y(_14838_));
 INVx1_ASAP7_75t_R _20173_ (.A(_00450_),
    .Y(_14839_));
 NAND2x1_ASAP7_75t_R _20174_ (.A(net386),
    .B(_00448_),
    .Y(_14840_));
 OA211x2_ASAP7_75t_R _20175_ (.A1(net386),
    .A2(_14839_),
    .B(_14840_),
    .C(net405),
    .Y(_14841_));
 OR3x1_ASAP7_75t_R _20176_ (.A(net298),
    .B(_14838_),
    .C(_14841_),
    .Y(_14842_));
 NAND2x1_ASAP7_75t_R _20177_ (.A(net386),
    .B(_01704_),
    .Y(_14843_));
 OA211x2_ASAP7_75t_R _20178_ (.A1(net386),
    .A2(_14118_),
    .B(_14843_),
    .C(net305),
    .Y(_14844_));
 AND3x1_ASAP7_75t_R _20179_ (.A(net405),
    .B(net302),
    .C(_14117_),
    .Y(_14845_));
 OA31x2_ASAP7_75t_R _20180_ (.A1(net300),
    .A2(_14844_),
    .A3(_14845_),
    .B1(net362),
    .Y(_14846_));
 AO32x1_ASAP7_75t_R _20181_ (.A1(_13392_),
    .A2(_14828_),
    .A3(_14834_),
    .B1(_14842_),
    .B2(_14846_),
    .Y(_14847_));
 NAND2x1_ASAP7_75t_R _20182_ (.A(net386),
    .B(_00457_),
    .Y(_14848_));
 OA211x2_ASAP7_75t_R _20183_ (.A1(net386),
    .A2(_14105_),
    .B(_14848_),
    .C(net305),
    .Y(_14849_));
 NAND2x1_ASAP7_75t_R _20184_ (.A(net386),
    .B(_00456_),
    .Y(_14850_));
 OA211x2_ASAP7_75t_R _20185_ (.A1(net386),
    .A2(_14098_),
    .B(_14850_),
    .C(net405),
    .Y(_14851_));
 OR3x1_ASAP7_75t_R _20186_ (.A(net373),
    .B(_14849_),
    .C(_14851_),
    .Y(_14852_));
 NAND2x1_ASAP7_75t_R _20187_ (.A(net401),
    .B(_00453_),
    .Y(_14853_));
 OA211x2_ASAP7_75t_R _20188_ (.A1(net401),
    .A2(_14108_),
    .B(_14853_),
    .C(net305),
    .Y(_14854_));
 NAND2x1_ASAP7_75t_R _20189_ (.A(net401),
    .B(_00452_),
    .Y(_14855_));
 OA211x2_ASAP7_75t_R _20190_ (.A1(net401),
    .A2(_14101_),
    .B(_14855_),
    .C(net405),
    .Y(_14856_));
 OR3x1_ASAP7_75t_R _20191_ (.A(_13397_),
    .B(_14854_),
    .C(_14856_),
    .Y(_14857_));
 AND2x2_ASAP7_75t_R _20192_ (.A(_14852_),
    .B(_14857_),
    .Y(_14858_));
 AND2x2_ASAP7_75t_R _20193_ (.A(_14842_),
    .B(_14846_),
    .Y(_14859_));
 NAND2x1_ASAP7_75t_R _20194_ (.A(net400),
    .B(_00473_),
    .Y(_14860_));
 OA211x2_ASAP7_75t_R _20195_ (.A1(net400),
    .A2(_14128_),
    .B(_14860_),
    .C(net307),
    .Y(_14861_));
 NAND2x1_ASAP7_75t_R _20196_ (.A(net400),
    .B(_00472_),
    .Y(_14862_));
 OA211x2_ASAP7_75t_R _20197_ (.A1(net400),
    .A2(_14131_),
    .B(_14862_),
    .C(net411),
    .Y(_14863_));
 OR3x1_ASAP7_75t_R _20198_ (.A(net373),
    .B(_14861_),
    .C(_14863_),
    .Y(_14864_));
 INVx1_ASAP7_75t_R _20199_ (.A(_00471_),
    .Y(_14865_));
 NAND2x1_ASAP7_75t_R _20200_ (.A(net400),
    .B(_00469_),
    .Y(_14866_));
 OA211x2_ASAP7_75t_R _20201_ (.A1(net400),
    .A2(_14865_),
    .B(_14866_),
    .C(net307),
    .Y(_14867_));
 INVx1_ASAP7_75t_R _20202_ (.A(_00470_),
    .Y(_14868_));
 NAND2x1_ASAP7_75t_R _20203_ (.A(net400),
    .B(_00468_),
    .Y(_14869_));
 OA211x2_ASAP7_75t_R _20204_ (.A1(net400),
    .A2(_14868_),
    .B(_14869_),
    .C(net411),
    .Y(_14870_));
 OR3x1_ASAP7_75t_R _20205_ (.A(_13397_),
    .B(_14867_),
    .C(_14870_),
    .Y(_14871_));
 AND3x1_ASAP7_75t_R _20206_ (.A(_14571_),
    .B(_14864_),
    .C(_14871_),
    .Y(_14872_));
 AO221x2_ASAP7_75t_R _20207_ (.A1(net366),
    .A2(_14847_),
    .B1(_14858_),
    .B2(_14859_),
    .C(_14872_),
    .Y(_14873_));
 BUFx16f_ASAP7_75t_R load_slew401 (.A(_00289_),
    .Y(net401));
 AO22x1_ASAP7_75t_R _20209_ (.A1(_13530_),
    .A2(_00670_),
    .B1(_01447_),
    .B2(_13533_),
    .Y(_14875_));
 INVx1_ASAP7_75t_R _20210_ (.A(_14875_),
    .Y(_14876_));
 OA211x2_ASAP7_75t_R _20211_ (.A1(_13763_),
    .A2(_14137_),
    .B(_14876_),
    .C(_13576_),
    .Y(_14877_));
 OA21x2_ASAP7_75t_R _20212_ (.A1(_00284_),
    .A2(_14873_),
    .B(_14877_),
    .Y(_14878_));
 AOI21x1_ASAP7_75t_R _20213_ (.A1(net294),
    .A2(_14823_),
    .B(_14878_),
    .Y(_17546_));
 INVx1_ASAP7_75t_R _20214_ (.A(_17546_),
    .Y(_16507_));
 INVx1_ASAP7_75t_R _20215_ (.A(_00177_),
    .Y(\cs_registers_i.pc_id_i[5] ));
 NOR2x1_ASAP7_75t_R _20216_ (.A(_01636_),
    .B(_13223_),
    .Y(_14879_));
 AOI21x1_ASAP7_75t_R _20217_ (.A1(_00177_),
    .A2(_13553_),
    .B(_13561_),
    .Y(_14880_));
 OAI22x1_ASAP7_75t_R _20218_ (.A1(_13782_),
    .A2(_14873_),
    .B1(_14879_),
    .B2(_14880_),
    .Y(_18133_));
 OR3x2_ASAP7_75t_R _20219_ (.A(_00670_),
    .B(net295),
    .C(_13574_),
    .Y(_14881_));
 OAI21x1_ASAP7_75t_R _20220_ (.A1(_13576_),
    .A2(_18133_),
    .B(_14881_),
    .Y(_17547_));
 INVx1_ASAP7_75t_R _20221_ (.A(_17547_),
    .Y(_16508_));
 OR3x1_ASAP7_75t_R _20222_ (.A(_00666_),
    .B(_02264_),
    .C(_02262_),
    .Y(_14882_));
 OA21x2_ASAP7_75t_R _20223_ (.A1(_00667_),
    .A2(_00666_),
    .B(_00669_),
    .Y(_14883_));
 OA21x2_ASAP7_75t_R _20224_ (.A1(_02264_),
    .A2(_14883_),
    .B(_02263_),
    .Y(_14884_));
 OA21x2_ASAP7_75t_R _20225_ (.A1(_14763_),
    .A2(_14882_),
    .B(_14884_),
    .Y(_16509_));
 INVx2_ASAP7_75t_R _20226_ (.A(_01635_),
    .Y(_14885_));
 NAND2x1_ASAP7_75t_R _20227_ (.A(net379),
    .B(_00494_),
    .Y(_14886_));
 OA211x2_ASAP7_75t_R _20228_ (.A1(net379),
    .A2(_14146_),
    .B(_14886_),
    .C(net406),
    .Y(_14887_));
 NAND2x1_ASAP7_75t_R _20229_ (.A(net379),
    .B(_00495_),
    .Y(_14888_));
 OA211x2_ASAP7_75t_R _20230_ (.A1(net379),
    .A2(_14143_),
    .B(_14888_),
    .C(net304),
    .Y(_14889_));
 OR3x1_ASAP7_75t_R _20231_ (.A(net298),
    .B(_14887_),
    .C(_14889_),
    .Y(_14890_));
 INVx1_ASAP7_75t_R _20232_ (.A(_00492_),
    .Y(_14891_));
 NAND2x1_ASAP7_75t_R _20233_ (.A(net384),
    .B(_00490_),
    .Y(_14892_));
 OA211x2_ASAP7_75t_R _20234_ (.A1(net384),
    .A2(_14891_),
    .B(_14892_),
    .C(net411),
    .Y(_14893_));
 INVx1_ASAP7_75t_R _20235_ (.A(_00493_),
    .Y(_14894_));
 NAND2x1_ASAP7_75t_R _20236_ (.A(net384),
    .B(_00491_),
    .Y(_14895_));
 OA211x2_ASAP7_75t_R _20237_ (.A1(net384),
    .A2(_14894_),
    .B(_14895_),
    .C(net305),
    .Y(_14896_));
 OR3x2_ASAP7_75t_R _20238_ (.A(net300),
    .B(_14893_),
    .C(_14896_),
    .Y(_14897_));
 AND3x1_ASAP7_75t_R _20239_ (.A(_13392_),
    .B(_14890_),
    .C(_14897_),
    .Y(_14898_));
 BUFx16f_ASAP7_75t_R max_cap400 (.A(net401),
    .Y(net400));
 OR2x2_ASAP7_75t_R _20241_ (.A(net378),
    .B(_00504_),
    .Y(_14900_));
 OAI21x1_ASAP7_75t_R _20242_ (.A1(_13433_),
    .A2(_00502_),
    .B(_14900_),
    .Y(_14901_));
 INVx1_ASAP7_75t_R _20243_ (.A(_00505_),
    .Y(_14902_));
 NAND2x1_ASAP7_75t_R _20244_ (.A(net379),
    .B(_00503_),
    .Y(_14903_));
 OA211x2_ASAP7_75t_R _20245_ (.A1(net379),
    .A2(_14902_),
    .B(_14903_),
    .C(net304),
    .Y(_14904_));
 AO21x1_ASAP7_75t_R _20246_ (.A1(net412),
    .A2(_14901_),
    .B(_14904_),
    .Y(_14905_));
 BUFx16f_ASAP7_75t_R load_slew399 (.A(net400),
    .Y(net399));
 NAND2x1_ASAP7_75t_R _20248_ (.A(net379),
    .B(_00499_),
    .Y(_14907_));
 OA211x2_ASAP7_75t_R _20249_ (.A1(net379),
    .A2(_14161_),
    .B(_14907_),
    .C(net304),
    .Y(_14908_));
 NAND2x1_ASAP7_75t_R _20250_ (.A(net378),
    .B(_00498_),
    .Y(_14909_));
 OA211x2_ASAP7_75t_R _20251_ (.A1(net378),
    .A2(_14164_),
    .B(_14909_),
    .C(net412),
    .Y(_14910_));
 OR3x1_ASAP7_75t_R _20252_ (.A(_13397_),
    .B(_14908_),
    .C(_14910_),
    .Y(_14911_));
 OA21x2_ASAP7_75t_R _20253_ (.A1(net374),
    .A2(_14905_),
    .B(_14911_),
    .Y(_14912_));
 NAND2x1_ASAP7_75t_R _20254_ (.A(net403),
    .B(_00478_),
    .Y(_14913_));
 OA211x2_ASAP7_75t_R _20255_ (.A1(net403),
    .A2(_14189_),
    .B(_14913_),
    .C(net412),
    .Y(_14914_));
 NAND2x1_ASAP7_75t_R _20256_ (.A(net403),
    .B(_00479_),
    .Y(_14915_));
 OA211x2_ASAP7_75t_R _20257_ (.A1(net403),
    .A2(_14192_),
    .B(_14915_),
    .C(net304),
    .Y(_14916_));
 OR3x1_ASAP7_75t_R _20258_ (.A(net298),
    .B(_14914_),
    .C(_14916_),
    .Y(_14917_));
 NAND2x1_ASAP7_75t_R _20259_ (.A(net379),
    .B(_01703_),
    .Y(_14918_));
 OA211x2_ASAP7_75t_R _20260_ (.A1(net379),
    .A2(_14184_),
    .B(_14918_),
    .C(net304),
    .Y(_14919_));
 BUFx16f_ASAP7_75t_R max_cap398 (.A(net399),
    .Y(net398));
 AND3x1_ASAP7_75t_R _20262_ (.A(net412),
    .B(_13433_),
    .C(_14183_),
    .Y(_14921_));
 OA31x2_ASAP7_75t_R _20263_ (.A1(net300),
    .A2(_14919_),
    .A3(_14921_),
    .B1(_00286_),
    .Y(_14922_));
 AO32x1_ASAP7_75t_R _20264_ (.A1(_13392_),
    .A2(_14890_),
    .A3(_14897_),
    .B1(_14917_),
    .B2(_14922_),
    .Y(_14923_));
 NAND2x1_ASAP7_75t_R _20265_ (.A(net379),
    .B(_00487_),
    .Y(_14924_));
 OA211x2_ASAP7_75t_R _20266_ (.A1(net379),
    .A2(_14176_),
    .B(_14924_),
    .C(net304),
    .Y(_14925_));
 NAND2x1_ASAP7_75t_R _20267_ (.A(net403),
    .B(_00486_),
    .Y(_14926_));
 OA211x2_ASAP7_75t_R _20268_ (.A1(net403),
    .A2(_14172_),
    .B(_14926_),
    .C(net412),
    .Y(_14927_));
 OR3x1_ASAP7_75t_R _20269_ (.A(net375),
    .B(_14925_),
    .C(_14927_),
    .Y(_14928_));
 INVx1_ASAP7_75t_R _20270_ (.A(_00485_),
    .Y(_14929_));
 NAND2x1_ASAP7_75t_R _20271_ (.A(net379),
    .B(_00483_),
    .Y(_14930_));
 OA211x2_ASAP7_75t_R _20272_ (.A1(net379),
    .A2(_14929_),
    .B(_14930_),
    .C(net304),
    .Y(_14931_));
 NAND2x1_ASAP7_75t_R _20273_ (.A(net403),
    .B(_00482_),
    .Y(_14932_));
 OA211x2_ASAP7_75t_R _20274_ (.A1(net403),
    .A2(_14169_),
    .B(_14932_),
    .C(net412),
    .Y(_14933_));
 OR3x1_ASAP7_75t_R _20275_ (.A(_13397_),
    .B(_14931_),
    .C(_14933_),
    .Y(_14934_));
 AND4x1_ASAP7_75t_R _20276_ (.A(_14917_),
    .B(_14922_),
    .C(_14928_),
    .D(_14934_),
    .Y(_14935_));
 AO221x2_ASAP7_75t_R _20277_ (.A1(_14898_),
    .A2(_14912_),
    .B1(_14923_),
    .B2(net368),
    .C(_14935_),
    .Y(_14936_));
 INVx2_ASAP7_75t_R _20278_ (.A(_00180_),
    .Y(_14937_));
 AO222x2_ASAP7_75t_R _20279_ (.A1(_14885_),
    .A2(_13270_),
    .B1(_13563_),
    .B2(_14936_),
    .C1(_14503_),
    .C2(_14937_),
    .Y(_14938_));
 BUFx16f_ASAP7_75t_R load_slew397 (.A(net399),
    .Y(net397));
 INVx2_ASAP7_75t_R _20281_ (.A(_14938_),
    .Y(_18138_));
 INVx2_ASAP7_75t_R _20282_ (.A(_00182_),
    .Y(\cs_registers_i.pc_id_i[7] ));
 INVx1_ASAP7_75t_R _20283_ (.A(_00515_),
    .Y(_14939_));
 NAND2x1_ASAP7_75t_R _20284_ (.A(_00289_),
    .B(_00513_),
    .Y(_14940_));
 OA211x2_ASAP7_75t_R _20285_ (.A1(_00289_),
    .A2(_14939_),
    .B(_14940_),
    .C(net307),
    .Y(_14941_));
 NAND2x1_ASAP7_75t_R _20286_ (.A(net401),
    .B(_00512_),
    .Y(_14942_));
 OA211x2_ASAP7_75t_R _20287_ (.A1(_00289_),
    .A2(_14227_),
    .B(_14942_),
    .C(net411),
    .Y(_14943_));
 NAND2x1_ASAP7_75t_R _20288_ (.A(net398),
    .B(_01702_),
    .Y(_14944_));
 OA211x2_ASAP7_75t_R _20289_ (.A1(net398),
    .A2(_14248_),
    .B(_14944_),
    .C(net306),
    .Y(_14945_));
 AND3x1_ASAP7_75t_R _20290_ (.A(_00290_),
    .B(net302),
    .C(_14251_),
    .Y(_14946_));
 OA33x2_ASAP7_75t_R _20291_ (.A1(_14743_),
    .A2(_14941_),
    .A3(_14943_),
    .B1(_14945_),
    .B2(_14946_),
    .B3(_13828_),
    .Y(_14947_));
 NAND2x1_ASAP7_75t_R _20292_ (.A(_00289_),
    .B(_00509_),
    .Y(_14948_));
 BUFx16f_ASAP7_75t_R load_slew396 (.A(net397),
    .Y(net396));
 OA211x2_ASAP7_75t_R _20294_ (.A1(_00289_),
    .A2(_14244_),
    .B(_14948_),
    .C(net307),
    .Y(_14950_));
 NAND2x1_ASAP7_75t_R _20295_ (.A(_00289_),
    .B(_00508_),
    .Y(_14951_));
 BUFx16f_ASAP7_75t_R load_slew395 (.A(net400),
    .Y(net395));
 OA211x2_ASAP7_75t_R _20297_ (.A1(_00289_),
    .A2(_14241_),
    .B(_14951_),
    .C(_00290_),
    .Y(_14953_));
 OR3x1_ASAP7_75t_R _20298_ (.A(_13484_),
    .B(_14950_),
    .C(_14953_),
    .Y(_14954_));
 NAND2x1_ASAP7_75t_R _20299_ (.A(_00289_),
    .B(_00517_),
    .Y(_14955_));
 OA211x2_ASAP7_75t_R _20300_ (.A1(_00289_),
    .A2(_14234_),
    .B(_14955_),
    .C(net307),
    .Y(_14956_));
 NAND2x1_ASAP7_75t_R _20301_ (.A(_00289_),
    .B(_00516_),
    .Y(_14957_));
 OA211x2_ASAP7_75t_R _20302_ (.A1(_00289_),
    .A2(_14230_),
    .B(_14957_),
    .C(net411),
    .Y(_14958_));
 OR3x1_ASAP7_75t_R _20303_ (.A(net367),
    .B(_14956_),
    .C(_14958_),
    .Y(_14959_));
 AO21x1_ASAP7_75t_R _20304_ (.A1(_14954_),
    .A2(_14959_),
    .B(net373),
    .Y(_14960_));
 AO21x2_ASAP7_75t_R _20305_ (.A1(_14947_),
    .A2(_14960_),
    .B(_13392_),
    .Y(_14961_));
 INVx1_ASAP7_75t_R _20306_ (.A(_00531_),
    .Y(_14962_));
 NAND2x1_ASAP7_75t_R _20307_ (.A(net411),
    .B(_00530_),
    .Y(_14963_));
 OA211x2_ASAP7_75t_R _20308_ (.A1(net411),
    .A2(_14962_),
    .B(_14963_),
    .C(net302),
    .Y(_14964_));
 INVx1_ASAP7_75t_R _20309_ (.A(_00529_),
    .Y(_14965_));
 NAND2x1_ASAP7_75t_R _20310_ (.A(net411),
    .B(_00528_),
    .Y(_14966_));
 OA211x2_ASAP7_75t_R _20311_ (.A1(net411),
    .A2(_14965_),
    .B(_14966_),
    .C(net400),
    .Y(_14967_));
 OR3x1_ASAP7_75t_R _20312_ (.A(_13397_),
    .B(_14964_),
    .C(_14967_),
    .Y(_14968_));
 NAND2x1_ASAP7_75t_R _20313_ (.A(net400),
    .B(_00533_),
    .Y(_14969_));
 OA211x2_ASAP7_75t_R _20314_ (.A1(net400),
    .A2(_14219_),
    .B(_14969_),
    .C(net307),
    .Y(_14970_));
 BUFx16f_ASAP7_75t_R wire394 (.A(net400),
    .Y(net394));
 NAND2x1_ASAP7_75t_R _20316_ (.A(net400),
    .B(_00532_),
    .Y(_14972_));
 OA211x2_ASAP7_75t_R _20317_ (.A1(net400),
    .A2(_14222_),
    .B(_14972_),
    .C(net411),
    .Y(_14973_));
 OR3x1_ASAP7_75t_R _20318_ (.A(net372),
    .B(_14970_),
    .C(_14973_),
    .Y(_14974_));
 AND3x1_ASAP7_75t_R _20319_ (.A(_13484_),
    .B(_14968_),
    .C(_14974_),
    .Y(_14975_));
 NAND2x1_ASAP7_75t_R _20320_ (.A(net400),
    .B(_00524_),
    .Y(_14976_));
 OA211x2_ASAP7_75t_R _20321_ (.A1(net400),
    .A2(_14201_),
    .B(_14976_),
    .C(_13397_),
    .Y(_14977_));
 INVx1_ASAP7_75t_R _20322_ (.A(_00522_),
    .Y(_14978_));
 NAND2x1_ASAP7_75t_R _20323_ (.A(net400),
    .B(_00520_),
    .Y(_14979_));
 OA211x2_ASAP7_75t_R _20324_ (.A1(net400),
    .A2(_14978_),
    .B(_14979_),
    .C(net372),
    .Y(_14980_));
 OR3x1_ASAP7_75t_R _20325_ (.A(net307),
    .B(_14977_),
    .C(_14980_),
    .Y(_14981_));
 INVx1_ASAP7_75t_R _20326_ (.A(_00523_),
    .Y(_14982_));
 NAND2x1_ASAP7_75t_R _20327_ (.A(net400),
    .B(_00521_),
    .Y(_14983_));
 OA211x2_ASAP7_75t_R _20328_ (.A1(net400),
    .A2(_14982_),
    .B(_14983_),
    .C(net372),
    .Y(_14984_));
 NAND2x1_ASAP7_75t_R _20329_ (.A(net399),
    .B(_00525_),
    .Y(_14985_));
 OA211x2_ASAP7_75t_R _20330_ (.A1(net399),
    .A2(_14204_),
    .B(_14985_),
    .C(_13397_),
    .Y(_14986_));
 OR3x1_ASAP7_75t_R _20331_ (.A(net411),
    .B(_14984_),
    .C(_14986_),
    .Y(_14987_));
 AND3x1_ASAP7_75t_R _20332_ (.A(net367),
    .B(_14981_),
    .C(_14987_),
    .Y(_14988_));
 OR3x4_ASAP7_75t_R _20333_ (.A(net362),
    .B(_14975_),
    .C(_14988_),
    .Y(_14989_));
 AND3x4_ASAP7_75t_R _20334_ (.A(_13563_),
    .B(_14961_),
    .C(_14989_),
    .Y(_14990_));
 INVx1_ASAP7_75t_R _20335_ (.A(_01634_),
    .Y(_14991_));
 AO32x2_ASAP7_75t_R _20336_ (.A1(\cs_registers_i.pc_id_i[7] ),
    .A2(_13553_),
    .A3(_14757_),
    .B1(_14991_),
    .B2(_13270_),
    .Y(_14992_));
 NOR2x2_ASAP7_75t_R _20337_ (.A(_14990_),
    .B(_14992_),
    .Y(_18143_));
 OA21x2_ASAP7_75t_R _20338_ (.A1(_00673_),
    .A2(_02266_),
    .B(_02265_),
    .Y(_14993_));
 OR3x1_ASAP7_75t_R _20339_ (.A(_00671_),
    .B(_02266_),
    .C(_16509_),
    .Y(_14994_));
 NAND2x1_ASAP7_75t_R _20340_ (.A(_14993_),
    .B(_14994_),
    .Y(_16512_));
 INVx1_ASAP7_75t_R _20341_ (.A(_01633_),
    .Y(_14995_));
 AND2x2_ASAP7_75t_R _20342_ (.A(_14995_),
    .B(_13270_),
    .Y(_14996_));
 BUFx12f_ASAP7_75t_R load_slew393 (.A(net394),
    .Y(net393));
 AOI21x1_ASAP7_75t_R _20344_ (.A1(_00186_),
    .A2(_13553_),
    .B(_13561_),
    .Y(_14998_));
 NAND2x1_ASAP7_75t_R _20345_ (.A(net402),
    .B(_00551_),
    .Y(_14999_));
 OA211x2_ASAP7_75t_R _20346_ (.A1(net402),
    .A2(_14263_),
    .B(_14999_),
    .C(net305),
    .Y(_15000_));
 NAND2x1_ASAP7_75t_R _20347_ (.A(net402),
    .B(_00550_),
    .Y(_15001_));
 OA211x2_ASAP7_75t_R _20348_ (.A1(net402),
    .A2(_14268_),
    .B(_15001_),
    .C(net411),
    .Y(_15002_));
 OR3x1_ASAP7_75t_R _20349_ (.A(_13397_),
    .B(_15000_),
    .C(_15002_),
    .Y(_15003_));
 NAND2x1_ASAP7_75t_R _20350_ (.A(net402),
    .B(_00555_),
    .Y(_15004_));
 OA211x2_ASAP7_75t_R _20351_ (.A1(net402),
    .A2(_14271_),
    .B(_15004_),
    .C(net305),
    .Y(_15005_));
 NAND2x1_ASAP7_75t_R _20352_ (.A(net402),
    .B(_00554_),
    .Y(_15006_));
 OA211x2_ASAP7_75t_R _20353_ (.A1(net402),
    .A2(_14259_),
    .B(_15006_),
    .C(net411),
    .Y(_15007_));
 OR3x1_ASAP7_75t_R _20354_ (.A(net374),
    .B(_15005_),
    .C(_15007_),
    .Y(_15008_));
 NAND2x1_ASAP7_75t_R _20355_ (.A(net402),
    .B(_00539_),
    .Y(_15009_));
 OA211x2_ASAP7_75t_R _20356_ (.A1(net402),
    .A2(_14302_),
    .B(_15009_),
    .C(net305),
    .Y(_15010_));
 NAND2x1_ASAP7_75t_R _20357_ (.A(net402),
    .B(_00538_),
    .Y(_15011_));
 OA211x2_ASAP7_75t_R _20358_ (.A1(net402),
    .A2(_14305_),
    .B(_15011_),
    .C(net411),
    .Y(_15012_));
 OR3x1_ASAP7_75t_R _20359_ (.A(net298),
    .B(_15010_),
    .C(_15012_),
    .Y(_15013_));
 NAND2x1_ASAP7_75t_R _20360_ (.A(net402),
    .B(_01701_),
    .Y(_15014_));
 OA211x2_ASAP7_75t_R _20361_ (.A1(net402),
    .A2(_14309_),
    .B(_15014_),
    .C(net305),
    .Y(_15015_));
 AND3x1_ASAP7_75t_R _20362_ (.A(net411),
    .B(_13433_),
    .C(_14312_),
    .Y(_15016_));
 OA31x2_ASAP7_75t_R _20363_ (.A1(net300),
    .A2(_15015_),
    .A3(_15016_),
    .B1(net363),
    .Y(_15017_));
 AO32x1_ASAP7_75t_R _20364_ (.A1(_13392_),
    .A2(_15003_),
    .A3(_15008_),
    .B1(_15013_),
    .B2(_15017_),
    .Y(_15018_));
 OR2x2_ASAP7_75t_R _20365_ (.A(net384),
    .B(_00544_),
    .Y(_15019_));
 OAI21x1_ASAP7_75t_R _20366_ (.A1(net303),
    .A2(_00542_),
    .B(_15019_),
    .Y(_15020_));
 NAND2x1_ASAP7_75t_R _20367_ (.A(net384),
    .B(_00543_),
    .Y(_15021_));
 OA211x2_ASAP7_75t_R _20368_ (.A1(net384),
    .A2(_14298_),
    .B(_15021_),
    .C(net304),
    .Y(_15022_));
 AO21x1_ASAP7_75t_R _20369_ (.A1(net412),
    .A2(_15020_),
    .B(_15022_),
    .Y(_15023_));
 NAND2x1_ASAP7_75t_R _20370_ (.A(net384),
    .B(_00547_),
    .Y(_15024_));
 OA211x2_ASAP7_75t_R _20371_ (.A1(net384),
    .A2(_14288_),
    .B(_15024_),
    .C(net304),
    .Y(_15025_));
 NAND2x1_ASAP7_75t_R _20372_ (.A(net384),
    .B(_00546_),
    .Y(_15026_));
 OA211x2_ASAP7_75t_R _20373_ (.A1(net384),
    .A2(_14291_),
    .B(_15026_),
    .C(net412),
    .Y(_15027_));
 OA21x2_ASAP7_75t_R _20374_ (.A1(_15025_),
    .A2(_15027_),
    .B(_13397_),
    .Y(_15028_));
 AO21x1_ASAP7_75t_R _20375_ (.A1(net374),
    .A2(_15023_),
    .B(_15028_),
    .Y(_15029_));
 AND2x2_ASAP7_75t_R _20376_ (.A(_15013_),
    .B(_15017_),
    .Y(_15030_));
 NAND2x1_ASAP7_75t_R _20377_ (.A(net384),
    .B(_00563_),
    .Y(_15031_));
 OA211x2_ASAP7_75t_R _20378_ (.A1(net384),
    .A2(_14281_),
    .B(_15031_),
    .C(net305),
    .Y(_15032_));
 NAND2x1_ASAP7_75t_R _20379_ (.A(net384),
    .B(_00562_),
    .Y(_15033_));
 OA211x2_ASAP7_75t_R _20380_ (.A1(net384),
    .A2(_14284_),
    .B(_15033_),
    .C(net412),
    .Y(_15034_));
 OR3x1_ASAP7_75t_R _20381_ (.A(net374),
    .B(_15032_),
    .C(_15034_),
    .Y(_15035_));
 NAND2x1_ASAP7_75t_R _20382_ (.A(net384),
    .B(_00559_),
    .Y(_15036_));
 OA211x2_ASAP7_75t_R _20383_ (.A1(net384),
    .A2(_14278_),
    .B(_15036_),
    .C(net305),
    .Y(_15037_));
 NAND2x1_ASAP7_75t_R _20384_ (.A(net384),
    .B(_00558_),
    .Y(_15038_));
 OA211x2_ASAP7_75t_R _20385_ (.A1(net384),
    .A2(_14275_),
    .B(_15038_),
    .C(net411),
    .Y(_15039_));
 OR3x1_ASAP7_75t_R _20386_ (.A(_13397_),
    .B(_15037_),
    .C(_15039_),
    .Y(_15040_));
 AND3x1_ASAP7_75t_R _20387_ (.A(_14571_),
    .B(_15035_),
    .C(_15040_),
    .Y(_15041_));
 AO221x2_ASAP7_75t_R _20388_ (.A1(net367),
    .A2(_15018_),
    .B1(_15029_),
    .B2(_15030_),
    .C(_15041_),
    .Y(_15042_));
 OAI22x1_ASAP7_75t_R _20389_ (.A1(_14996_),
    .A2(_14998_),
    .B1(_15042_),
    .B2(_13782_),
    .Y(_18148_));
 XOR2x1_ASAP7_75t_R _20390_ (.A(_13387_),
    .Y(_15043_),
    .B(_14376_));
 INVx1_ASAP7_75t_R _20391_ (.A(_15043_),
    .Y(_15044_));
 NAND2x1_ASAP7_75t_R _20392_ (.A(net378),
    .B(_00585_),
    .Y(_15045_));
 OA211x2_ASAP7_75t_R _20393_ (.A1(net378),
    .A2(_14360_),
    .B(_15045_),
    .C(net304),
    .Y(_15046_));
 INVx1_ASAP7_75t_R _20394_ (.A(_00586_),
    .Y(_15047_));
 NAND2x1_ASAP7_75t_R _20395_ (.A(net378),
    .B(_00584_),
    .Y(_15048_));
 OA211x2_ASAP7_75t_R _20396_ (.A1(net378),
    .A2(_15047_),
    .B(_15048_),
    .C(net406),
    .Y(_15049_));
 OR3x1_ASAP7_75t_R _20397_ (.A(net298),
    .B(_15046_),
    .C(_15049_),
    .Y(_15050_));
 NAND2x1_ASAP7_75t_R _20398_ (.A(net378),
    .B(_00580_),
    .Y(_15051_));
 OA211x2_ASAP7_75t_R _20399_ (.A1(net378),
    .A2(_14363_),
    .B(_15051_),
    .C(net406),
    .Y(_15052_));
 INVx1_ASAP7_75t_R _20400_ (.A(_00583_),
    .Y(_15053_));
 NAND2x1_ASAP7_75t_R _20401_ (.A(net378),
    .B(_00581_),
    .Y(_15054_));
 OA211x2_ASAP7_75t_R _20402_ (.A1(net378),
    .A2(_15053_),
    .B(_15054_),
    .C(net304),
    .Y(_15055_));
 OR3x1_ASAP7_75t_R _20403_ (.A(net300),
    .B(_15052_),
    .C(_15055_),
    .Y(_15056_));
 AND3x1_ASAP7_75t_R _20404_ (.A(_13392_),
    .B(_15050_),
    .C(_15056_),
    .Y(_15057_));
 OR2x2_ASAP7_75t_R _20405_ (.A(net378),
    .B(_00594_),
    .Y(_15058_));
 OAI21x1_ASAP7_75t_R _20406_ (.A1(_13433_),
    .A2(_00592_),
    .B(_15058_),
    .Y(_15059_));
 INVx1_ASAP7_75t_R _20407_ (.A(_00595_),
    .Y(_15060_));
 NAND2x1_ASAP7_75t_R _20408_ (.A(net378),
    .B(_00593_),
    .Y(_15061_));
 OA211x2_ASAP7_75t_R _20409_ (.A1(net378),
    .A2(_15060_),
    .B(_15061_),
    .C(net304),
    .Y(_15062_));
 AO21x1_ASAP7_75t_R _20410_ (.A1(net412),
    .A2(_15059_),
    .B(_15062_),
    .Y(_15063_));
 BUFx16f_ASAP7_75t_R load_slew392 (.A(net400),
    .Y(net392));
 INVx1_ASAP7_75t_R _20412_ (.A(_00591_),
    .Y(_15065_));
 NAND2x1_ASAP7_75t_R _20413_ (.A(net378),
    .B(_00589_),
    .Y(_15066_));
 OA211x2_ASAP7_75t_R _20414_ (.A1(net378),
    .A2(_15065_),
    .B(_15066_),
    .C(net304),
    .Y(_15067_));
 BUFx16f_ASAP7_75t_R load_slew391 (.A(net392),
    .Y(net391));
 NAND2x1_ASAP7_75t_R _20416_ (.A(net378),
    .B(_00588_),
    .Y(_15069_));
 OA211x2_ASAP7_75t_R _20417_ (.A1(net378),
    .A2(_14353_),
    .B(_15069_),
    .C(net412),
    .Y(_15070_));
 OR3x1_ASAP7_75t_R _20418_ (.A(_13397_),
    .B(_15067_),
    .C(_15070_),
    .Y(_15071_));
 OA21x2_ASAP7_75t_R _20419_ (.A1(net374),
    .A2(_15063_),
    .B(_15071_),
    .Y(_15072_));
 NAND2x1_ASAP7_75t_R _20420_ (.A(net379),
    .B(_00568_),
    .Y(_15073_));
 OA211x2_ASAP7_75t_R _20421_ (.A1(net379),
    .A2(_14339_),
    .B(_15073_),
    .C(net412),
    .Y(_15074_));
 NAND2x1_ASAP7_75t_R _20422_ (.A(net379),
    .B(_00569_),
    .Y(_15075_));
 OA211x2_ASAP7_75t_R _20423_ (.A1(net379),
    .A2(_14342_),
    .B(_15075_),
    .C(net304),
    .Y(_15076_));
 OR3x1_ASAP7_75t_R _20424_ (.A(net298),
    .B(_15074_),
    .C(_15076_),
    .Y(_15077_));
 NAND2x1_ASAP7_75t_R _20425_ (.A(net378),
    .B(_01700_),
    .Y(_15078_));
 OA211x2_ASAP7_75t_R _20426_ (.A1(net378),
    .A2(_14346_),
    .B(_15078_),
    .C(net304),
    .Y(_15079_));
 INVx1_ASAP7_75t_R _20427_ (.A(_00566_),
    .Y(_15080_));
 AND3x1_ASAP7_75t_R _20428_ (.A(net406),
    .B(_13433_),
    .C(_15080_),
    .Y(_15081_));
 OA31x2_ASAP7_75t_R _20429_ (.A1(net300),
    .A2(_15079_),
    .A3(_15081_),
    .B1(_00286_),
    .Y(_15082_));
 AO32x1_ASAP7_75t_R _20430_ (.A1(_13392_),
    .A2(_15050_),
    .A3(_15056_),
    .B1(_15077_),
    .B2(_15082_),
    .Y(_15083_));
 NAND2x1_ASAP7_75t_R _20431_ (.A(net379),
    .B(_00577_),
    .Y(_15084_));
 OA211x2_ASAP7_75t_R _20432_ (.A1(net379),
    .A2(_14325_),
    .B(_15084_),
    .C(net304),
    .Y(_15085_));
 NAND2x1_ASAP7_75t_R _20433_ (.A(net379),
    .B(_00576_),
    .Y(_15086_));
 OA211x2_ASAP7_75t_R _20434_ (.A1(net379),
    .A2(_14335_),
    .B(_15086_),
    .C(net412),
    .Y(_15087_));
 OR3x1_ASAP7_75t_R _20435_ (.A(net375),
    .B(_15085_),
    .C(_15087_),
    .Y(_15088_));
 INVx1_ASAP7_75t_R _20436_ (.A(_00575_),
    .Y(_15089_));
 NAND2x1_ASAP7_75t_R _20437_ (.A(net379),
    .B(_00573_),
    .Y(_15090_));
 OA211x2_ASAP7_75t_R _20438_ (.A1(net379),
    .A2(_15089_),
    .B(_15090_),
    .C(net304),
    .Y(_15091_));
 NAND2x1_ASAP7_75t_R _20439_ (.A(net379),
    .B(_00572_),
    .Y(_15092_));
 OA211x2_ASAP7_75t_R _20440_ (.A1(net379),
    .A2(_14332_),
    .B(_15092_),
    .C(net412),
    .Y(_15093_));
 OR3x1_ASAP7_75t_R _20441_ (.A(_13397_),
    .B(_15091_),
    .C(_15093_),
    .Y(_15094_));
 AND4x1_ASAP7_75t_R _20442_ (.A(_15077_),
    .B(_15082_),
    .C(_15088_),
    .D(_15094_),
    .Y(_15095_));
 AO221x2_ASAP7_75t_R _20443_ (.A1(_15057_),
    .A2(_15072_),
    .B1(_15083_),
    .B2(net368),
    .C(_15095_),
    .Y(_15096_));
 NOR2x1_ASAP7_75t_R _20444_ (.A(_00284_),
    .B(_15096_),
    .Y(_15097_));
 BUFx16f_ASAP7_75t_R load_slew390 (.A(net391),
    .Y(net390));
 AO221x1_ASAP7_75t_R _20446_ (.A1(_13530_),
    .A2(_00680_),
    .B1(_01443_),
    .B2(_13533_),
    .C(_13528_),
    .Y(_15099_));
 NAND2x1_ASAP7_75t_R _20447_ (.A(_13528_),
    .B(_14373_),
    .Y(_15100_));
 OA211x2_ASAP7_75t_R _20448_ (.A1(_15097_),
    .A2(_15099_),
    .B(_13576_),
    .C(_15100_),
    .Y(_15101_));
 AO21x1_ASAP7_75t_R _20449_ (.A1(net294),
    .A2(_15044_),
    .B(_15101_),
    .Y(_17552_));
 INVx1_ASAP7_75t_R _20450_ (.A(_17552_),
    .Y(_16513_));
 INVx1_ASAP7_75t_R _20451_ (.A(_00189_),
    .Y(\cs_registers_i.pc_id_i[9] ));
 OA211x2_ASAP7_75t_R _20452_ (.A1(_13549_),
    .A2(_13552_),
    .B(_00189_),
    .C(_13223_),
    .Y(_15102_));
 OAI22x1_ASAP7_75t_R _20453_ (.A1(_01632_),
    .A2(_13223_),
    .B1(_13561_),
    .B2(_15102_),
    .Y(_15103_));
 OA21x2_ASAP7_75t_R _20454_ (.A1(_13782_),
    .A2(_15096_),
    .B(_15103_),
    .Y(_15104_));
 BUFx16f_ASAP7_75t_R load_slew389 (.A(net392),
    .Y(net389));
 INVx2_ASAP7_75t_R _20456_ (.A(_15104_),
    .Y(_18153_));
 OR3x1_ASAP7_75t_R _20457_ (.A(_00680_),
    .B(net295),
    .C(_13574_),
    .Y(_15105_));
 OAI21x1_ASAP7_75t_R _20458_ (.A1(_13576_),
    .A2(_18153_),
    .B(_15105_),
    .Y(_17553_));
 INVx1_ASAP7_75t_R _20459_ (.A(_17553_),
    .Y(_16514_));
 OR2x2_ASAP7_75t_R _20460_ (.A(_00675_),
    .B(_02268_),
    .Y(_15106_));
 AO21x1_ASAP7_75t_R _20461_ (.A1(_14993_),
    .A2(_14994_),
    .B(_15106_),
    .Y(_15107_));
 OA21x2_ASAP7_75t_R _20462_ (.A1(_00678_),
    .A2(_02268_),
    .B(_02267_),
    .Y(_15108_));
 AND2x2_ASAP7_75t_R _20463_ (.A(_15107_),
    .B(_15108_),
    .Y(_16515_));
 INVx2_ASAP7_75t_R _20464_ (.A(_01631_),
    .Y(_15109_));
 NAND2x1_ASAP7_75t_R _20465_ (.A(net395),
    .B(_00615_),
    .Y(_15110_));
 OA211x2_ASAP7_75t_R _20466_ (.A1(net395),
    .A2(_14421_),
    .B(_15110_),
    .C(net307),
    .Y(_15111_));
 NAND2x1_ASAP7_75t_R _20467_ (.A(net395),
    .B(_00614_),
    .Y(_15112_));
 OA211x2_ASAP7_75t_R _20468_ (.A1(net395),
    .A2(_14424_),
    .B(_15112_),
    .C(net405),
    .Y(_15113_));
 OR3x1_ASAP7_75t_R _20469_ (.A(net373),
    .B(_15111_),
    .C(_15113_),
    .Y(_15114_));
 INVx1_ASAP7_75t_R _20470_ (.A(_00613_),
    .Y(_15115_));
 NAND2x1_ASAP7_75t_R _20471_ (.A(net385),
    .B(_00611_),
    .Y(_15116_));
 OA211x2_ASAP7_75t_R _20472_ (.A1(net385),
    .A2(_15115_),
    .B(_15116_),
    .C(net305),
    .Y(_15117_));
 INVx1_ASAP7_75t_R _20473_ (.A(_00612_),
    .Y(_15118_));
 NAND2x1_ASAP7_75t_R _20474_ (.A(net385),
    .B(_00610_),
    .Y(_15119_));
 OA211x2_ASAP7_75t_R _20475_ (.A1(net385),
    .A2(_15118_),
    .B(_15119_),
    .C(net405),
    .Y(_15120_));
 OR3x1_ASAP7_75t_R _20476_ (.A(_13397_),
    .B(_15117_),
    .C(_15120_),
    .Y(_15121_));
 NAND2x1_ASAP7_75t_R _20477_ (.A(net395),
    .B(_00598_),
    .Y(_15122_));
 OA211x2_ASAP7_75t_R _20478_ (.A1(net395),
    .A2(_14398_),
    .B(_15122_),
    .C(net405),
    .Y(_15123_));
 NAND2x1_ASAP7_75t_R _20479_ (.A(net395),
    .B(_00599_),
    .Y(_15124_));
 OA211x2_ASAP7_75t_R _20480_ (.A1(net395),
    .A2(_14395_),
    .B(_15124_),
    .C(net307),
    .Y(_15125_));
 OR3x1_ASAP7_75t_R _20481_ (.A(net298),
    .B(_15123_),
    .C(_15125_),
    .Y(_15126_));
 NAND2x1_ASAP7_75t_R _20482_ (.A(net385),
    .B(_01699_),
    .Y(_15127_));
 OA211x2_ASAP7_75t_R _20483_ (.A1(net385),
    .A2(_14403_),
    .B(_15127_),
    .C(net307),
    .Y(_15128_));
 AND3x1_ASAP7_75t_R _20484_ (.A(net405),
    .B(net302),
    .C(_14402_),
    .Y(_15129_));
 OA31x2_ASAP7_75t_R _20485_ (.A1(net300),
    .A2(_15128_),
    .A3(_15129_),
    .B1(net362),
    .Y(_15130_));
 AO32x1_ASAP7_75t_R _20486_ (.A1(_13392_),
    .A2(_15114_),
    .A3(_15121_),
    .B1(_15126_),
    .B2(_15130_),
    .Y(_15131_));
 NOR2x1_ASAP7_75t_R _20487_ (.A(net401),
    .B(_00608_),
    .Y(_15132_));
 AO21x1_ASAP7_75t_R _20488_ (.A1(net401),
    .A2(_14386_),
    .B(_15132_),
    .Y(_15133_));
 NAND2x1_ASAP7_75t_R _20489_ (.A(net401),
    .B(_00607_),
    .Y(_15134_));
 OA211x2_ASAP7_75t_R _20490_ (.A1(net401),
    .A2(_14390_),
    .B(_15134_),
    .C(net307),
    .Y(_15135_));
 AO21x1_ASAP7_75t_R _20491_ (.A1(net405),
    .A2(_15133_),
    .B(_15135_),
    .Y(_15136_));
 NAND2x1_ASAP7_75t_R _20492_ (.A(net395),
    .B(_00603_),
    .Y(_15137_));
 OA211x2_ASAP7_75t_R _20493_ (.A1(net395),
    .A2(_14377_),
    .B(_15137_),
    .C(net307),
    .Y(_15138_));
 NAND2x1_ASAP7_75t_R _20494_ (.A(net395),
    .B(_00602_),
    .Y(_15139_));
 OA211x2_ASAP7_75t_R _20495_ (.A1(net395),
    .A2(_14381_),
    .B(_15139_),
    .C(net405),
    .Y(_15140_));
 OA21x2_ASAP7_75t_R _20496_ (.A1(_15138_),
    .A2(_15140_),
    .B(net373),
    .Y(_15141_));
 AO21x1_ASAP7_75t_R _20497_ (.A1(_13397_),
    .A2(_15136_),
    .B(_15141_),
    .Y(_15142_));
 AND2x2_ASAP7_75t_R _20498_ (.A(_15126_),
    .B(_15130_),
    .Y(_15143_));
 INVx1_ASAP7_75t_R _20499_ (.A(_00625_),
    .Y(_15144_));
 NAND2x1_ASAP7_75t_R _20500_ (.A(net385),
    .B(_00623_),
    .Y(_15145_));
 OA211x2_ASAP7_75t_R _20501_ (.A1(net385),
    .A2(_15144_),
    .B(_15145_),
    .C(net305),
    .Y(_15146_));
 INVx1_ASAP7_75t_R _20502_ (.A(_00624_),
    .Y(_15147_));
 NAND2x1_ASAP7_75t_R _20503_ (.A(net385),
    .B(_00622_),
    .Y(_15148_));
 OA211x2_ASAP7_75t_R _20504_ (.A1(net385),
    .A2(_15147_),
    .B(_15148_),
    .C(net405),
    .Y(_15149_));
 OR3x1_ASAP7_75t_R _20505_ (.A(net373),
    .B(_15146_),
    .C(_15149_),
    .Y(_15150_));
 NAND2x1_ASAP7_75t_R _20506_ (.A(net385),
    .B(_00619_),
    .Y(_15151_));
 OA211x2_ASAP7_75t_R _20507_ (.A1(net385),
    .A2(_14409_),
    .B(_15151_),
    .C(net305),
    .Y(_15152_));
 NAND2x1_ASAP7_75t_R _20508_ (.A(net385),
    .B(_00618_),
    .Y(_15153_));
 OA211x2_ASAP7_75t_R _20509_ (.A1(net385),
    .A2(_14412_),
    .B(_15153_),
    .C(net405),
    .Y(_15154_));
 OR3x1_ASAP7_75t_R _20510_ (.A(_13397_),
    .B(_15152_),
    .C(_15154_),
    .Y(_15155_));
 AND3x1_ASAP7_75t_R _20511_ (.A(_14571_),
    .B(_15150_),
    .C(_15155_),
    .Y(_15156_));
 AO221x2_ASAP7_75t_R _20512_ (.A1(net366),
    .A2(_15131_),
    .B1(_15142_),
    .B2(_15143_),
    .C(_15156_),
    .Y(_15157_));
 INVx2_ASAP7_75t_R _20513_ (.A(_00193_),
    .Y(_15158_));
 AO222x2_ASAP7_75t_R _20514_ (.A1(_15109_),
    .A2(_13270_),
    .B1(_13563_),
    .B2(_15157_),
    .C1(_14503_),
    .C2(_15158_),
    .Y(_15159_));
 BUFx16f_ASAP7_75t_R max_cap388 (.A(net389),
    .Y(net388));
 INVx2_ASAP7_75t_R _20516_ (.A(_15159_),
    .Y(_18158_));
 INVx2_ASAP7_75t_R _20517_ (.A(_14489_),
    .Y(_15160_));
 NOR2x1_ASAP7_75t_R _20518_ (.A(_00284_),
    .B(_14574_),
    .Y(_15161_));
 BUFx16f_ASAP7_75t_R load_slew387 (.A(net395),
    .Y(net387));
 AO221x1_ASAP7_75t_R _20520_ (.A1(_13530_),
    .A2(_00684_),
    .B1(_01441_),
    .B2(_13533_),
    .C(_13528_),
    .Y(_15163_));
 OA22x2_ASAP7_75t_R _20521_ (.A1(_13763_),
    .A2(_15160_),
    .B1(_15161_),
    .B2(_15163_),
    .Y(_15164_));
 XNOR2x1_ASAP7_75t_R _20522_ (.B(_18162_),
    .Y(_15165_),
    .A(_13387_));
 AND2x2_ASAP7_75t_R _20523_ (.A(net294),
    .B(_15165_),
    .Y(_15166_));
 AO21x1_ASAP7_75t_R _20524_ (.A1(_13576_),
    .A2(_15164_),
    .B(_15166_),
    .Y(_17557_));
 INVx1_ASAP7_75t_R _20525_ (.A(_17557_),
    .Y(_16518_));
 OA21x2_ASAP7_75t_R _20526_ (.A1(_00684_),
    .A2(_13574_),
    .B(_13576_),
    .Y(_15167_));
 AOI21x1_ASAP7_75t_R _20527_ (.A1(net294),
    .A2(_14576_),
    .B(_15167_),
    .Y(_17556_));
 INVx1_ASAP7_75t_R _20528_ (.A(_17556_),
    .Y(_16516_));
 OA21x2_ASAP7_75t_R _20529_ (.A1(_00681_),
    .A2(_16515_),
    .B(_00683_),
    .Y(_15168_));
 OA21x2_ASAP7_75t_R _20530_ (.A1(_02270_),
    .A2(_15168_),
    .B(_02269_),
    .Y(_16517_));
 BUFx16f_ASAP7_75t_R load_slew386 (.A(net401),
    .Y(net386));
 BUFx16f_ASAP7_75t_R load_slew385 (.A(net386),
    .Y(net385));
 BUFx16f_ASAP7_75t_R max_cap384 (.A(net402),
    .Y(net384));
 BUFx16f_ASAP7_75t_R wire383 (.A(net384),
    .Y(net383));
 BUFx16f_ASAP7_75t_R load_slew382 (.A(net383),
    .Y(net382));
 BUFx16f_ASAP7_75t_R load_slew381 (.A(net383),
    .Y(net381));
 BUFx16f_ASAP7_75t_R load_slew380 (.A(net381),
    .Y(net380));
 BUFx16f_ASAP7_75t_R load_slew379 (.A(net403),
    .Y(net379));
 BUFx16f_ASAP7_75t_R max_cap378 (.A(net379),
    .Y(net378));
 BUFx16f_ASAP7_75t_R load_slew377 (.A(net379),
    .Y(net377));
 BUFx16f_ASAP7_75t_R load_slew376 (.A(net378),
    .Y(net376));
 BUFx16f_ASAP7_75t_R max_cap375 (.A(_00288_),
    .Y(net375));
 AND2x2_ASAP7_75t_R _20543_ (.A(net327),
    .B(_01697_),
    .Y(_15181_));
 AO21x1_ASAP7_75t_R _20544_ (.A1(net312),
    .A2(_00326_),
    .B(_15181_),
    .Y(_15182_));
 BUFx16f_ASAP7_75t_R max_cap374 (.A(_00288_),
    .Y(net374));
 BUFx16f_ASAP7_75t_R load_slew373 (.A(net374),
    .Y(net373));
 BUFx12f_ASAP7_75t_R load_slew372 (.A(net373),
    .Y(net372));
 BUFx16f_ASAP7_75t_R load_slew371 (.A(net372),
    .Y(net371));
 OAI22x1_ASAP7_75t_R _20549_ (.A1(_00325_),
    .A2(_13586_),
    .B1(_15182_),
    .B2(net354),
    .Y(_15187_));
 BUFx16f_ASAP7_75t_R wire370 (.A(net372),
    .Y(net370));
 BUFx16f_ASAP7_75t_R load_slew369 (.A(net373),
    .Y(net369));
 BUFx12f_ASAP7_75t_R load_slew368 (.A(_00287_),
    .Y(net368));
 BUFx16f_ASAP7_75t_R load_slew367 (.A(_00287_),
    .Y(net367));
 BUFx12f_ASAP7_75t_R load_slew366 (.A(net367),
    .Y(net366));
 BUFx16f_ASAP7_75t_R load_slew365 (.A(net367),
    .Y(net365));
 BUFx16f_ASAP7_75t_R load_slew364 (.A(_00286_),
    .Y(net364));
 NAND2x1_ASAP7_75t_R _20557_ (.A(net327),
    .B(_00332_),
    .Y(_15195_));
 BUFx16f_ASAP7_75t_R load_slew363 (.A(_00286_),
    .Y(net363));
 BUFx12f_ASAP7_75t_R load_slew362 (.A(net363),
    .Y(net362));
 OA211x2_ASAP7_75t_R _20560_ (.A1(net327),
    .A2(_13802_),
    .B(_15195_),
    .C(net311),
    .Y(_15198_));
 NAND2x1_ASAP7_75t_R _20561_ (.A(net327),
    .B(_00331_),
    .Y(_15199_));
 BUFx16f_ASAP7_75t_R load_slew361 (.A(_00246_),
    .Y(net361));
 OA211x2_ASAP7_75t_R _20563_ (.A1(net327),
    .A2(_13808_),
    .B(_15199_),
    .C(net354),
    .Y(_15201_));
 OR3x1_ASAP7_75t_R _20564_ (.A(net321),
    .B(_15198_),
    .C(_15201_),
    .Y(_15202_));
 BUFx12f_ASAP7_75t_R load_slew360 (.A(net361),
    .Y(net360));
 BUFx16f_ASAP7_75t_R load_slew359 (.A(net360),
    .Y(net359));
 BUFx16f_ASAP7_75t_R load_slew358 (.A(net359),
    .Y(net358));
 OA211x2_ASAP7_75t_R _20568_ (.A1(_13598_),
    .A2(_15187_),
    .B(_15202_),
    .C(net323),
    .Y(_15206_));
 BUFx16f_ASAP7_75t_R wire357 (.A(net359),
    .Y(net357));
 BUFx16f_ASAP7_75t_R load_slew356 (.A(net357),
    .Y(net356));
 BUFx16f_ASAP7_75t_R load_slew355 (.A(net356),
    .Y(net355));
 BUFx16f_ASAP7_75t_R load_slew354 (.A(_00246_),
    .Y(net354));
 BUFx16f_ASAP7_75t_R load_slew353 (.A(_01745_),
    .Y(net353));
 BUFx16f_ASAP7_75t_R max_cap352 (.A(net353),
    .Y(net352));
 NOR2x1_ASAP7_75t_R _20575_ (.A(net327),
    .B(_00337_),
    .Y(_15213_));
 AO21x1_ASAP7_75t_R _20576_ (.A1(net327),
    .A2(_13789_),
    .B(_15213_),
    .Y(_15214_));
 BUFx16f_ASAP7_75t_R max_cap351 (.A(net352),
    .Y(net351));
 BUFx16f_ASAP7_75t_R load_slew350 (.A(net352),
    .Y(net350));
 BUFx16f_ASAP7_75t_R load_slew349 (.A(net350),
    .Y(net349));
 NAND2x1_ASAP7_75t_R _20580_ (.A(net327),
    .B(_00336_),
    .Y(_15218_));
 BUFx16f_ASAP7_75t_R load_slew348 (.A(net350),
    .Y(net348));
 BUFx16f_ASAP7_75t_R max_cap347 (.A(net348),
    .Y(net347));
 OA211x2_ASAP7_75t_R _20583_ (.A1(net327),
    .A2(_13794_),
    .B(_15218_),
    .C(net311),
    .Y(_15221_));
 AO21x1_ASAP7_75t_R _20584_ (.A1(net354),
    .A2(_15214_),
    .B(_15221_),
    .Y(_15222_));
 NAND2x1_ASAP7_75t_R _20585_ (.A(net327),
    .B(_00328_),
    .Y(_15223_));
 OA211x2_ASAP7_75t_R _20586_ (.A1(net327),
    .A2(_13821_),
    .B(_15223_),
    .C(net311),
    .Y(_15224_));
 BUFx16f_ASAP7_75t_R load_slew346 (.A(net347),
    .Y(net346));
 BUFx16f_ASAP7_75t_R load_slew345 (.A(net346),
    .Y(net345));
 NAND2x1_ASAP7_75t_R _20589_ (.A(net327),
    .B(_00327_),
    .Y(_15227_));
 OA211x2_ASAP7_75t_R _20590_ (.A1(net327),
    .A2(_13818_),
    .B(_15227_),
    .C(net354),
    .Y(_15228_));
 OR3x1_ASAP7_75t_R _20591_ (.A(_13598_),
    .B(_15224_),
    .C(_15228_),
    .Y(_15229_));
 BUFx16f_ASAP7_75t_R load_slew344 (.A(net345),
    .Y(net344));
 BUFx16f_ASAP7_75t_R load_slew343 (.A(net348),
    .Y(net343));
 OA211x2_ASAP7_75t_R _20594_ (.A1(net321),
    .A2(_15222_),
    .B(_15229_),
    .C(_13132_),
    .Y(_15232_));
 OR3x1_ASAP7_75t_R _20595_ (.A(_13174_),
    .B(_15206_),
    .C(_15232_),
    .Y(_15233_));
 BUFx16f_ASAP7_75t_R load_slew342 (.A(net343),
    .Y(net342));
 BUFx16f_ASAP7_75t_R load_slew341 (.A(net351),
    .Y(net341));
 NAND2x1_ASAP7_75t_R _20598_ (.A(net327),
    .B(_00340_),
    .Y(_15236_));
 OA211x2_ASAP7_75t_R _20599_ (.A1(net327),
    .A2(_13847_),
    .B(_15236_),
    .C(net311),
    .Y(_15237_));
 BUFx16f_ASAP7_75t_R load_slew340 (.A(net341),
    .Y(net340));
 BUFx16f_ASAP7_75t_R load_slew339 (.A(net340),
    .Y(net339));
 BUFx16f_ASAP7_75t_R load_slew338 (.A(net339),
    .Y(net338));
 NAND2x1_ASAP7_75t_R _20603_ (.A(net327),
    .B(_00339_),
    .Y(_15241_));
 BUFx16f_ASAP7_75t_R load_slew337 (.A(net338),
    .Y(net337));
 OA211x2_ASAP7_75t_R _20605_ (.A1(net327),
    .A2(_13835_),
    .B(_15241_),
    .C(net354),
    .Y(_15243_));
 OR3x1_ASAP7_75t_R _20606_ (.A(_13132_),
    .B(_15237_),
    .C(_15243_),
    .Y(_15244_));
 NAND2x1_ASAP7_75t_R _20607_ (.A(net327),
    .B(_00344_),
    .Y(_15245_));
 BUFx12f_ASAP7_75t_R load_slew336 (.A(net337),
    .Y(net336));
 OA211x2_ASAP7_75t_R _20609_ (.A1(net327),
    .A2(_13852_),
    .B(_15245_),
    .C(net311),
    .Y(_15247_));
 NAND2x1_ASAP7_75t_R _20610_ (.A(net327),
    .B(_00343_),
    .Y(_15248_));
 OA211x2_ASAP7_75t_R _20611_ (.A1(net327),
    .A2(_13839_),
    .B(_15248_),
    .C(net354),
    .Y(_15249_));
 OR3x1_ASAP7_75t_R _20612_ (.A(net323),
    .B(_15247_),
    .C(_15249_),
    .Y(_15250_));
 AND3x1_ASAP7_75t_R _20613_ (.A(net321),
    .B(_15244_),
    .C(_15250_),
    .Y(_15251_));
 NAND2x1_ASAP7_75t_R _20614_ (.A(net327),
    .B(_00352_),
    .Y(_15252_));
 OA211x2_ASAP7_75t_R _20615_ (.A1(net327),
    .A2(_13872_),
    .B(_15252_),
    .C(net311),
    .Y(_15253_));
 NAND2x1_ASAP7_75t_R _20616_ (.A(net327),
    .B(_00351_),
    .Y(_15254_));
 OA211x2_ASAP7_75t_R _20617_ (.A1(net327),
    .A2(_13864_),
    .B(_15254_),
    .C(net354),
    .Y(_15255_));
 OR3x1_ASAP7_75t_R _20618_ (.A(net322),
    .B(_15253_),
    .C(_15255_),
    .Y(_15256_));
 NAND2x1_ASAP7_75t_R _20619_ (.A(net327),
    .B(_00348_),
    .Y(_15257_));
 OA211x2_ASAP7_75t_R _20620_ (.A1(net327),
    .A2(_13868_),
    .B(_15257_),
    .C(net311),
    .Y(_15258_));
 BUFx16f_ASAP7_75t_R load_slew335 (.A(net340),
    .Y(net335));
 BUFx16f_ASAP7_75t_R load_slew334 (.A(net335),
    .Y(net334));
 NAND2x1_ASAP7_75t_R _20623_ (.A(net327),
    .B(_00347_),
    .Y(_15261_));
 OA211x2_ASAP7_75t_R _20624_ (.A1(net327),
    .A2(_13860_),
    .B(_15261_),
    .C(net354),
    .Y(_15262_));
 OR3x1_ASAP7_75t_R _20625_ (.A(_13132_),
    .B(_15258_),
    .C(_15262_),
    .Y(_15263_));
 AND3x1_ASAP7_75t_R _20626_ (.A(_13598_),
    .B(_15256_),
    .C(_15263_),
    .Y(_15264_));
 OR3x2_ASAP7_75t_R _20627_ (.A(net314),
    .B(_15251_),
    .C(_15264_),
    .Y(_15265_));
 NAND2x2_ASAP7_75t_R _20628_ (.A(_15233_),
    .B(_15265_),
    .Y(_15266_));
 NAND2x2_ASAP7_75t_R _20629_ (.A(_13223_),
    .B(_13275_),
    .Y(_15267_));
 OA21x2_ASAP7_75t_R _20630_ (.A1(_13298_),
    .A2(_13653_),
    .B(_15267_),
    .Y(_15268_));
 OA21x2_ASAP7_75t_R _20631_ (.A1(_00280_),
    .A2(_13282_),
    .B(_13299_),
    .Y(_15269_));
 OA21x2_ASAP7_75t_R _20632_ (.A1(_00281_),
    .A2(_15268_),
    .B(_15269_),
    .Y(_15270_));
 AOI21x1_ASAP7_75t_R _20633_ (.A1(_13583_),
    .A2(_15266_),
    .B(_15270_),
    .Y(_18166_));
 BUFx16f_ASAP7_75t_R max_cap333 (.A(net334),
    .Y(net333));
 BUFx16f_ASAP7_75t_R load_slew332 (.A(net335),
    .Y(net332));
 BUFx16f_ASAP7_75t_R load_slew331 (.A(net332),
    .Y(net331));
 BUFx16f_ASAP7_75t_R load_slew330 (.A(net353),
    .Y(net330));
 BUFx16f_ASAP7_75t_R load_slew329 (.A(net330),
    .Y(net329));
 INVx1_ASAP7_75t_R _20639_ (.A(_00698_),
    .Y(_15276_));
 BUFx16f_ASAP7_75t_R load_slew328 (.A(net329),
    .Y(net328));
 NOR2x1_ASAP7_75t_R _20641_ (.A(net332),
    .B(_00700_),
    .Y(_15278_));
 AO21x1_ASAP7_75t_R _20642_ (.A1(net332),
    .A2(_15276_),
    .B(_15278_),
    .Y(_15279_));
 BUFx16f_ASAP7_75t_R load_slew327 (.A(net329),
    .Y(net327));
 INVx1_ASAP7_75t_R _20644_ (.A(_00701_),
    .Y(_15281_));
 BUFx16f_ASAP7_75t_R load_slew326 (.A(net353),
    .Y(net326));
 BUFx16f_ASAP7_75t_R load_slew325 (.A(_01744_),
    .Y(net325));
 NAND2x1_ASAP7_75t_R _20647_ (.A(net332),
    .B(_00699_),
    .Y(_15284_));
 BUFx16f_ASAP7_75t_R load_slew324 (.A(_01744_),
    .Y(net324));
 BUFx16f_ASAP7_75t_R load_slew323 (.A(_01744_),
    .Y(net323));
 OA211x2_ASAP7_75t_R _20650_ (.A1(net332),
    .A2(_15281_),
    .B(_15284_),
    .C(net310),
    .Y(_15287_));
 AO21x1_ASAP7_75t_R _20651_ (.A1(net356),
    .A2(_15279_),
    .B(_15287_),
    .Y(_15288_));
 BUFx16f_ASAP7_75t_R wire322 (.A(_01744_),
    .Y(net322));
 BUFx16f_ASAP7_75t_R load_slew321 (.A(_00245_),
    .Y(net321));
 BUFx16f_ASAP7_75t_R load_slew320 (.A(_00245_),
    .Y(net320));
 INVx1_ASAP7_75t_R _20655_ (.A(_00693_),
    .Y(_15292_));
 NAND2x1_ASAP7_75t_R _20656_ (.A(net332),
    .B(_00691_),
    .Y(_15293_));
 BUFx16f_ASAP7_75t_R load_slew319 (.A(net320),
    .Y(net319));
 OA211x2_ASAP7_75t_R _20658_ (.A1(net332),
    .A2(_15292_),
    .B(_15293_),
    .C(net308),
    .Y(_15295_));
 INVx1_ASAP7_75t_R _20659_ (.A(_00692_),
    .Y(_15296_));
 NAND2x1_ASAP7_75t_R _20660_ (.A(net332),
    .B(_00690_),
    .Y(_15297_));
 OA211x2_ASAP7_75t_R _20661_ (.A1(net332),
    .A2(_15296_),
    .B(_15297_),
    .C(net356),
    .Y(_15298_));
 OR3x1_ASAP7_75t_R _20662_ (.A(_13598_),
    .B(_15295_),
    .C(_15298_),
    .Y(_15299_));
 OA21x2_ASAP7_75t_R _20663_ (.A1(net318),
    .A2(_15288_),
    .B(_15299_),
    .Y(_15300_));
 INVx1_ASAP7_75t_R _20664_ (.A(_00688_),
    .Y(_15301_));
 INVx1_ASAP7_75t_R _20665_ (.A(_00689_),
    .Y(_15302_));
 NAND2x1_ASAP7_75t_R _20666_ (.A(net332),
    .B(_01696_),
    .Y(_15303_));
 BUFx16f_ASAP7_75t_R load_slew318 (.A(net319),
    .Y(net318));
 OA211x2_ASAP7_75t_R _20668_ (.A1(net332),
    .A2(_15302_),
    .B(_15303_),
    .C(net310),
    .Y(_15305_));
 AO21x1_ASAP7_75t_R _20669_ (.A1(_15301_),
    .A2(_13190_),
    .B(_15305_),
    .Y(_15306_));
 INVx1_ASAP7_75t_R _20670_ (.A(_00697_),
    .Y(_15307_));
 NAND2x1_ASAP7_75t_R _20671_ (.A(net332),
    .B(_00695_),
    .Y(_15308_));
 OA211x2_ASAP7_75t_R _20672_ (.A1(net332),
    .A2(_15307_),
    .B(_15308_),
    .C(net308),
    .Y(_15309_));
 INVx1_ASAP7_75t_R _20673_ (.A(_00696_),
    .Y(_15310_));
 NAND2x1_ASAP7_75t_R _20674_ (.A(net332),
    .B(_00694_),
    .Y(_15311_));
 OA211x2_ASAP7_75t_R _20675_ (.A1(net332),
    .A2(_15310_),
    .B(_15311_),
    .C(net356),
    .Y(_15312_));
 OR3x1_ASAP7_75t_R _20676_ (.A(net318),
    .B(_15309_),
    .C(_15312_),
    .Y(_15313_));
 OA211x2_ASAP7_75t_R _20677_ (.A1(_13598_),
    .A2(_15306_),
    .B(_15313_),
    .C(net325),
    .Y(_15314_));
 AO21x1_ASAP7_75t_R _20678_ (.A1(_13132_),
    .A2(_15300_),
    .B(_15314_),
    .Y(_15315_));
 BUFx12f_ASAP7_75t_R load_slew317 (.A(net320),
    .Y(net317));
 INVx1_ASAP7_75t_R _20680_ (.A(_00705_),
    .Y(_15317_));
 BUFx12f_ASAP7_75t_R load_slew316 (.A(_00244_),
    .Y(net316));
 NAND2x1_ASAP7_75t_R _20682_ (.A(net344),
    .B(_00703_),
    .Y(_15319_));
 OA211x2_ASAP7_75t_R _20683_ (.A1(net344),
    .A2(_15317_),
    .B(_15319_),
    .C(net308),
    .Y(_15320_));
 BUFx12f_ASAP7_75t_R load_slew315 (.A(net316),
    .Y(net315));
 INVx1_ASAP7_75t_R _20685_ (.A(_00704_),
    .Y(_15322_));
 NAND2x1_ASAP7_75t_R _20686_ (.A(net344),
    .B(_00702_),
    .Y(_15323_));
 OA211x2_ASAP7_75t_R _20687_ (.A1(net344),
    .A2(_15322_),
    .B(_15323_),
    .C(net356),
    .Y(_15324_));
 OR3x1_ASAP7_75t_R _20688_ (.A(_13132_),
    .B(_15320_),
    .C(_15324_),
    .Y(_15325_));
 BUFx16f_ASAP7_75t_R load_slew314 (.A(net316),
    .Y(net314));
 INVx1_ASAP7_75t_R _20690_ (.A(_00709_),
    .Y(_15327_));
 NAND2x1_ASAP7_75t_R _20691_ (.A(net344),
    .B(_00707_),
    .Y(_15328_));
 OA211x2_ASAP7_75t_R _20692_ (.A1(net344),
    .A2(_15327_),
    .B(_15328_),
    .C(net308),
    .Y(_15329_));
 BUFx16f_ASAP7_75t_R max_length313 (.A(_13127_),
    .Y(net313));
 INVx1_ASAP7_75t_R _20694_ (.A(_00708_),
    .Y(_15331_));
 NAND2x1_ASAP7_75t_R _20695_ (.A(net344),
    .B(_00706_),
    .Y(_15332_));
 OA211x2_ASAP7_75t_R _20696_ (.A1(net344),
    .A2(_15331_),
    .B(_15332_),
    .C(net356),
    .Y(_15333_));
 OR3x1_ASAP7_75t_R _20697_ (.A(net325),
    .B(_15329_),
    .C(_15333_),
    .Y(_15334_));
 AND3x1_ASAP7_75t_R _20698_ (.A(net318),
    .B(_15325_),
    .C(_15334_),
    .Y(_15335_));
 INVx1_ASAP7_75t_R _20699_ (.A(_00712_),
    .Y(_15336_));
 NAND2x1_ASAP7_75t_R _20700_ (.A(net344),
    .B(_00710_),
    .Y(_15337_));
 OA211x2_ASAP7_75t_R _20701_ (.A1(net344),
    .A2(_15336_),
    .B(_15337_),
    .C(net356),
    .Y(_15338_));
 INVx1_ASAP7_75t_R _20702_ (.A(_00713_),
    .Y(_15339_));
 NAND2x1_ASAP7_75t_R _20703_ (.A(net344),
    .B(_00711_),
    .Y(_15340_));
 OA211x2_ASAP7_75t_R _20704_ (.A1(net344),
    .A2(_15339_),
    .B(_15340_),
    .C(net308),
    .Y(_15341_));
 OR3x1_ASAP7_75t_R _20705_ (.A(_13132_),
    .B(_15338_),
    .C(_15341_),
    .Y(_15342_));
 INVx1_ASAP7_75t_R _20706_ (.A(_00717_),
    .Y(_15343_));
 NAND2x1_ASAP7_75t_R _20707_ (.A(net344),
    .B(_00715_),
    .Y(_15344_));
 OA211x2_ASAP7_75t_R _20708_ (.A1(net344),
    .A2(_15343_),
    .B(_15344_),
    .C(_13145_),
    .Y(_15345_));
 INVx1_ASAP7_75t_R _20709_ (.A(_00716_),
    .Y(_15346_));
 NAND2x1_ASAP7_75t_R _20710_ (.A(net344),
    .B(_00714_),
    .Y(_15347_));
 OA211x2_ASAP7_75t_R _20711_ (.A1(net344),
    .A2(_15346_),
    .B(_15347_),
    .C(net356),
    .Y(_15348_));
 OR3x1_ASAP7_75t_R _20712_ (.A(net325),
    .B(_15345_),
    .C(_15348_),
    .Y(_15349_));
 AND3x1_ASAP7_75t_R _20713_ (.A(_13598_),
    .B(_15342_),
    .C(_15349_),
    .Y(_15350_));
 OR3x1_ASAP7_75t_R _20714_ (.A(net315),
    .B(_15335_),
    .C(_15350_),
    .Y(_15351_));
 OAI21x1_ASAP7_75t_R _20715_ (.A1(_13174_),
    .A2(_15315_),
    .B(_15351_),
    .Y(_15352_));
 BUFx16f_ASAP7_75t_R max_length312 (.A(net313),
    .Y(net312));
 OA21x2_ASAP7_75t_R _20717_ (.A1(_00282_),
    .A2(_15268_),
    .B(_15269_),
    .Y(_15354_));
 AO21x2_ASAP7_75t_R _20718_ (.A1(_13583_),
    .A2(_15352_),
    .B(_15354_),
    .Y(_18173_));
 INVx1_ASAP7_75t_R _20719_ (.A(_18173_),
    .Y(_18171_));
 XNOR2x1_ASAP7_75t_R _20720_ (.B(_18173_),
    .Y(_15355_),
    .A(_13387_));
 NOR2x1_ASAP7_75t_R _20721_ (.A(_13763_),
    .B(_15352_),
    .Y(_15356_));
 NAND2x1_ASAP7_75t_R _20722_ (.A(net389),
    .B(_00703_),
    .Y(_15357_));
 OA211x2_ASAP7_75t_R _20723_ (.A1(net389),
    .A2(_15317_),
    .B(_15357_),
    .C(net306),
    .Y(_15358_));
 NAND2x1_ASAP7_75t_R _20724_ (.A(net389),
    .B(_00702_),
    .Y(_15359_));
 OA211x2_ASAP7_75t_R _20725_ (.A1(net389),
    .A2(_15322_),
    .B(_15359_),
    .C(net409),
    .Y(_15360_));
 OR3x1_ASAP7_75t_R _20726_ (.A(_13397_),
    .B(_15358_),
    .C(_15360_),
    .Y(_15361_));
 NAND2x1_ASAP7_75t_R _20727_ (.A(net389),
    .B(_00707_),
    .Y(_15362_));
 OA211x2_ASAP7_75t_R _20728_ (.A1(net389),
    .A2(_15327_),
    .B(_15362_),
    .C(_13424_),
    .Y(_15363_));
 NAND2x1_ASAP7_75t_R _20729_ (.A(net389),
    .B(_00706_),
    .Y(_15364_));
 OA211x2_ASAP7_75t_R _20730_ (.A1(net389),
    .A2(_15331_),
    .B(_15364_),
    .C(net409),
    .Y(_15365_));
 OR3x1_ASAP7_75t_R _20731_ (.A(net370),
    .B(_15363_),
    .C(_15365_),
    .Y(_15366_));
 NAND2x1_ASAP7_75t_R _20732_ (.A(net391),
    .B(_00690_),
    .Y(_15367_));
 OA211x2_ASAP7_75t_R _20733_ (.A1(net391),
    .A2(_15296_),
    .B(_15367_),
    .C(net409),
    .Y(_15368_));
 NAND2x1_ASAP7_75t_R _20734_ (.A(net391),
    .B(_00691_),
    .Y(_15369_));
 OA211x2_ASAP7_75t_R _20735_ (.A1(net391),
    .A2(_15292_),
    .B(_15369_),
    .C(net306),
    .Y(_15370_));
 OR3x1_ASAP7_75t_R _20736_ (.A(_13814_),
    .B(_15368_),
    .C(_15370_),
    .Y(_15371_));
 NAND2x1_ASAP7_75t_R _20737_ (.A(net391),
    .B(_01696_),
    .Y(_15372_));
 OA211x2_ASAP7_75t_R _20738_ (.A1(net391),
    .A2(_15302_),
    .B(_15372_),
    .C(net306),
    .Y(_15373_));
 AND3x1_ASAP7_75t_R _20739_ (.A(net409),
    .B(net302),
    .C(_15301_),
    .Y(_15374_));
 OA31x2_ASAP7_75t_R _20740_ (.A1(_13828_),
    .A2(_15373_),
    .A3(_15374_),
    .B1(net362),
    .Y(_15375_));
 AO32x1_ASAP7_75t_R _20741_ (.A1(_13392_),
    .A2(_15361_),
    .A3(_15366_),
    .B1(_15371_),
    .B2(_15375_),
    .Y(_15376_));
 NOR2x1_ASAP7_75t_R _20742_ (.A(net391),
    .B(_00700_),
    .Y(_15377_));
 AO21x1_ASAP7_75t_R _20743_ (.A1(net391),
    .A2(_15276_),
    .B(_15377_),
    .Y(_15378_));
 BUFx16f_ASAP7_75t_R max_length311 (.A(_13145_),
    .Y(net311));
 NAND2x1_ASAP7_75t_R _20745_ (.A(net391),
    .B(_00699_),
    .Y(_15380_));
 OA211x2_ASAP7_75t_R _20746_ (.A1(net391),
    .A2(_15281_),
    .B(_15380_),
    .C(net306),
    .Y(_15381_));
 AO21x1_ASAP7_75t_R _20747_ (.A1(net409),
    .A2(_15378_),
    .B(_15381_),
    .Y(_15382_));
 NAND2x1_ASAP7_75t_R _20748_ (.A(net391),
    .B(_00695_),
    .Y(_15383_));
 OA211x2_ASAP7_75t_R _20749_ (.A1(net391),
    .A2(_15307_),
    .B(_15383_),
    .C(net306),
    .Y(_15384_));
 NAND2x1_ASAP7_75t_R _20750_ (.A(net391),
    .B(_00694_),
    .Y(_15385_));
 OA211x2_ASAP7_75t_R _20751_ (.A1(net391),
    .A2(_15310_),
    .B(_15385_),
    .C(net409),
    .Y(_15386_));
 OA21x2_ASAP7_75t_R _20752_ (.A1(_15384_),
    .A2(_15386_),
    .B(net370),
    .Y(_15387_));
 AO21x1_ASAP7_75t_R _20753_ (.A1(_13397_),
    .A2(_15382_),
    .B(_15387_),
    .Y(_15388_));
 AND2x2_ASAP7_75t_R _20754_ (.A(_15371_),
    .B(_15375_),
    .Y(_15389_));
 NAND2x1_ASAP7_75t_R _20755_ (.A(net390),
    .B(_00715_),
    .Y(_15390_));
 OA211x2_ASAP7_75t_R _20756_ (.A1(net390),
    .A2(_15343_),
    .B(_15390_),
    .C(_13424_),
    .Y(_15391_));
 NAND2x1_ASAP7_75t_R _20757_ (.A(net389),
    .B(_00714_),
    .Y(_15392_));
 OA211x2_ASAP7_75t_R _20758_ (.A1(net389),
    .A2(_15346_),
    .B(_15392_),
    .C(net409),
    .Y(_15393_));
 OR3x1_ASAP7_75t_R _20759_ (.A(net370),
    .B(_15391_),
    .C(_15393_),
    .Y(_15394_));
 NAND2x1_ASAP7_75t_R _20760_ (.A(net389),
    .B(_00711_),
    .Y(_15395_));
 OA211x2_ASAP7_75t_R _20761_ (.A1(net389),
    .A2(_15339_),
    .B(_15395_),
    .C(_13424_),
    .Y(_15396_));
 NAND2x1_ASAP7_75t_R _20762_ (.A(net389),
    .B(_00710_),
    .Y(_15397_));
 OA211x2_ASAP7_75t_R _20763_ (.A1(net389),
    .A2(_15336_),
    .B(_15397_),
    .C(net409),
    .Y(_15398_));
 OR3x1_ASAP7_75t_R _20764_ (.A(_13397_),
    .B(_15396_),
    .C(_15398_),
    .Y(_15399_));
 AND3x1_ASAP7_75t_R _20765_ (.A(_14571_),
    .B(_15394_),
    .C(_15399_),
    .Y(_15400_));
 AO221x2_ASAP7_75t_R _20766_ (.A1(net365),
    .A2(_15376_),
    .B1(_15388_),
    .B2(_15389_),
    .C(_15400_),
    .Y(_15401_));
 BUFx16f_ASAP7_75t_R max_length310 (.A(_13145_),
    .Y(net310));
 AOI22x1_ASAP7_75t_R _20768_ (.A1(_13530_),
    .A2(_00718_),
    .B1(_02220_),
    .B2(_13533_),
    .Y(_15403_));
 OA211x2_ASAP7_75t_R _20769_ (.A1(_00284_),
    .A2(_15401_),
    .B(_15403_),
    .C(_13763_),
    .Y(_15404_));
 OA21x2_ASAP7_75t_R _20770_ (.A1(_15356_),
    .A2(_15404_),
    .B(_13576_),
    .Y(_15405_));
 AOI21x1_ASAP7_75t_R _20771_ (.A1(net295),
    .A2(_15355_),
    .B(_15405_),
    .Y(_17561_));
 INVx1_ASAP7_75t_R _20772_ (.A(_17561_),
    .Y(_16520_));
 INVx3_ASAP7_75t_R _20773_ (.A(_00201_),
    .Y(\cs_registers_i.pc_id_i[13] ));
 NOR2x1_ASAP7_75t_R _20774_ (.A(_01628_),
    .B(_13223_),
    .Y(_15406_));
 AOI221x1_ASAP7_75t_R _20775_ (.A1(\cs_registers_i.pc_id_i[13] ),
    .A2(_14503_),
    .B1(_15401_),
    .B2(_13563_),
    .C(_15406_),
    .Y(_15407_));
 BUFx16f_ASAP7_75t_R max_length309 (.A(net310),
    .Y(net309));
 BUFx16f_ASAP7_75t_R max_length308 (.A(_13145_),
    .Y(net308));
 OA21x2_ASAP7_75t_R _20778_ (.A1(_00718_),
    .A2(_13574_),
    .B(_13576_),
    .Y(_15409_));
 AOI21x1_ASAP7_75t_R _20779_ (.A1(net295),
    .A2(_15407_),
    .B(_15409_),
    .Y(_17560_));
 INVx1_ASAP7_75t_R _20780_ (.A(_17560_),
    .Y(_16519_));
 AO21x1_ASAP7_75t_R _20781_ (.A1(_00673_),
    .A2(_00671_),
    .B(_02266_),
    .Y(_15410_));
 OR4x1_ASAP7_75t_R _20782_ (.A(_00681_),
    .B(_00685_),
    .C(_02270_),
    .D(_02272_),
    .Y(_15411_));
 OR2x2_ASAP7_75t_R _20783_ (.A(_15106_),
    .B(_15411_),
    .Y(_15412_));
 AO221x1_ASAP7_75t_R _20784_ (.A1(_16509_),
    .A2(_14993_),
    .B1(_15410_),
    .B2(_02265_),
    .C(_15412_),
    .Y(_15413_));
 OA21x2_ASAP7_75t_R _20785_ (.A1(_00683_),
    .A2(_02270_),
    .B(_02269_),
    .Y(_15414_));
 OR3x1_ASAP7_75t_R _20786_ (.A(_00685_),
    .B(_02272_),
    .C(_15414_),
    .Y(_15415_));
 OA21x2_ASAP7_75t_R _20787_ (.A1(_00687_),
    .A2(_02272_),
    .B(_02271_),
    .Y(_15416_));
 OA211x2_ASAP7_75t_R _20788_ (.A1(_15108_),
    .A2(_15411_),
    .B(_15415_),
    .C(_15416_),
    .Y(_15417_));
 AND2x2_ASAP7_75t_R _20789_ (.A(_15413_),
    .B(_15417_),
    .Y(_16521_));
 BUFx16f_ASAP7_75t_R max_length307 (.A(_13424_),
    .Y(net307));
 BUFx16f_ASAP7_75t_R max_length306 (.A(net307),
    .Y(net306));
 BUFx16f_ASAP7_75t_R wire305 (.A(net307),
    .Y(net305));
 INVx1_ASAP7_75t_R _20793_ (.A(_00729_),
    .Y(_15421_));
 BUFx16f_ASAP7_75t_R max_length304 (.A(net305),
    .Y(net304));
 NAND2x1_ASAP7_75t_R _20795_ (.A(net328),
    .B(_00727_),
    .Y(_15423_));
 BUFx16f_ASAP7_75t_R max_length303 (.A(_13433_),
    .Y(net303));
 OA211x2_ASAP7_75t_R _20797_ (.A1(net328),
    .A2(_15421_),
    .B(_15423_),
    .C(net310),
    .Y(_15425_));
 BUFx16f_ASAP7_75t_R max_length302 (.A(net303),
    .Y(net302));
 BUFx16f_ASAP7_75t_R load_slew301 (.A(_13828_),
    .Y(net301));
 INVx1_ASAP7_75t_R _20800_ (.A(_00728_),
    .Y(_15428_));
 NAND2x1_ASAP7_75t_R _20801_ (.A(net326),
    .B(_00726_),
    .Y(_15429_));
 BUFx12f_ASAP7_75t_R load_slew300 (.A(net301),
    .Y(net300));
 BUFx10_ASAP7_75t_R load_slew299 (.A(_02290_),
    .Y(net299));
 OA211x2_ASAP7_75t_R _20804_ (.A1(net326),
    .A2(_15428_),
    .B(_15429_),
    .C(_00246_),
    .Y(_15432_));
 OR3x1_ASAP7_75t_R _20805_ (.A(net321),
    .B(_15425_),
    .C(_15432_),
    .Y(_15433_));
 INVx1_ASAP7_75t_R _20806_ (.A(_00720_),
    .Y(_15434_));
 INVx1_ASAP7_75t_R _20807_ (.A(_00721_),
    .Y(_15435_));
 BUFx16f_ASAP7_75t_R load_slew298 (.A(_13814_),
    .Y(net298));
 NAND2x1_ASAP7_75t_R _20809_ (.A(net328),
    .B(_01695_),
    .Y(_15437_));
 OA21x2_ASAP7_75t_R _20810_ (.A1(net328),
    .A2(_15435_),
    .B(_15437_),
    .Y(_15438_));
 BUFx10_ASAP7_75t_R max_cap297 (.A(_12699_),
    .Y(net297));
 AO221x1_ASAP7_75t_R _20812_ (.A1(_15434_),
    .A2(_13190_),
    .B1(_15438_),
    .B2(net311),
    .C(_13598_),
    .Y(_15440_));
 AND2x2_ASAP7_75t_R _20813_ (.A(_15433_),
    .B(_15440_),
    .Y(_15441_));
 BUFx16f_ASAP7_75t_R max_cap296 (.A(_12723_),
    .Y(net296));
 BUFx16f_ASAP7_75t_R wire295 (.A(_13318_),
    .Y(net295));
 INVx1_ASAP7_75t_R _20816_ (.A(_00725_),
    .Y(_15444_));
 NAND2x1_ASAP7_75t_R _20817_ (.A(net326),
    .B(_00723_),
    .Y(_15445_));
 BUFx16f_ASAP7_75t_R load_slew294 (.A(net295),
    .Y(net294));
 OA211x2_ASAP7_75t_R _20819_ (.A1(net326),
    .A2(_15444_),
    .B(_15445_),
    .C(net310),
    .Y(_15447_));
 INVx1_ASAP7_75t_R _20820_ (.A(_00724_),
    .Y(_15448_));
 NAND2x1_ASAP7_75t_R _20821_ (.A(net326),
    .B(_00722_),
    .Y(_15449_));
 BUFx12f_ASAP7_75t_R load_slew293 (.A(_02286_),
    .Y(net293));
 OA211x2_ASAP7_75t_R _20823_ (.A1(net326),
    .A2(_15448_),
    .B(_15449_),
    .C(_00246_),
    .Y(_15451_));
 OR3x1_ASAP7_75t_R _20824_ (.A(_13598_),
    .B(_15447_),
    .C(_15451_),
    .Y(_15452_));
 INVx1_ASAP7_75t_R _20825_ (.A(_00733_),
    .Y(_15453_));
 NAND2x1_ASAP7_75t_R _20826_ (.A(net326),
    .B(_00731_),
    .Y(_15454_));
 OA211x2_ASAP7_75t_R _20827_ (.A1(net326),
    .A2(_15453_),
    .B(_15454_),
    .C(net311),
    .Y(_15455_));
 INVx1_ASAP7_75t_R _20828_ (.A(_00732_),
    .Y(_15456_));
 NAND2x1_ASAP7_75t_R _20829_ (.A(net326),
    .B(_00730_),
    .Y(_15457_));
 OA211x2_ASAP7_75t_R _20830_ (.A1(net326),
    .A2(_15456_),
    .B(_15457_),
    .C(_00246_),
    .Y(_15458_));
 OR3x1_ASAP7_75t_R _20831_ (.A(net321),
    .B(_15455_),
    .C(_15458_),
    .Y(_15459_));
 BUFx12f_ASAP7_75t_R max_cap292 (.A(net293),
    .Y(net292));
 AO21x1_ASAP7_75t_R _20833_ (.A1(_15452_),
    .A2(_15459_),
    .B(net322),
    .Y(_15461_));
 OA211x2_ASAP7_75t_R _20834_ (.A1(_13132_),
    .A2(_15441_),
    .B(_15461_),
    .C(_00244_),
    .Y(_15462_));
 BUFx12f_ASAP7_75t_R load_slew291 (.A(_02289_),
    .Y(net291));
 BUFx6f_ASAP7_75t_R load_slew290 (.A(_13656_),
    .Y(net290));
 INVx1_ASAP7_75t_R _20837_ (.A(_00741_),
    .Y(_15465_));
 NAND2x1_ASAP7_75t_R _20838_ (.A(net328),
    .B(_00739_),
    .Y(_15466_));
 BUFx16f_ASAP7_75t_R load_slew289 (.A(_13656_),
    .Y(net289));
 OA211x2_ASAP7_75t_R _20840_ (.A1(net328),
    .A2(_15465_),
    .B(_15466_),
    .C(net311),
    .Y(_15468_));
 INVx1_ASAP7_75t_R _20841_ (.A(_00740_),
    .Y(_15469_));
 BUFx12f_ASAP7_75t_R load_slew288 (.A(net290),
    .Y(net288));
 NAND2x1_ASAP7_75t_R _20843_ (.A(net328),
    .B(_00738_),
    .Y(_15471_));
 BUFx16f_ASAP7_75t_R load_slew287 (.A(_06226_),
    .Y(net287));
 OA211x2_ASAP7_75t_R _20845_ (.A1(net328),
    .A2(_15469_),
    .B(_15471_),
    .C(_00246_),
    .Y(_15473_));
 OR3x1_ASAP7_75t_R _20846_ (.A(net322),
    .B(_15468_),
    .C(_15473_),
    .Y(_15474_));
 INVx1_ASAP7_75t_R _20847_ (.A(_00737_),
    .Y(_15475_));
 NAND2x1_ASAP7_75t_R _20848_ (.A(net328),
    .B(_00735_),
    .Y(_15476_));
 OA211x2_ASAP7_75t_R _20849_ (.A1(net328),
    .A2(_15475_),
    .B(_15476_),
    .C(net311),
    .Y(_15477_));
 INVx1_ASAP7_75t_R _20850_ (.A(_00736_),
    .Y(_15478_));
 NAND2x1_ASAP7_75t_R _20851_ (.A(net328),
    .B(_00734_),
    .Y(_15479_));
 OA211x2_ASAP7_75t_R _20852_ (.A1(net328),
    .A2(_15478_),
    .B(_15479_),
    .C(_00246_),
    .Y(_15480_));
 OR3x1_ASAP7_75t_R _20853_ (.A(_13132_),
    .B(_15477_),
    .C(_15480_),
    .Y(_15481_));
 AND3x1_ASAP7_75t_R _20854_ (.A(net321),
    .B(_15474_),
    .C(_15481_),
    .Y(_15482_));
 BUFx16f_ASAP7_75t_R load_slew286 (.A(net287),
    .Y(net286));
 BUFx12f_ASAP7_75t_R max_cap285 (.A(_07206_),
    .Y(net285));
 INVx1_ASAP7_75t_R _20857_ (.A(_00744_),
    .Y(_15485_));
 BUFx16f_ASAP7_75t_R wire284 (.A(_07159_),
    .Y(net284));
 BUFx16f_ASAP7_75t_R max_cap283 (.A(net284),
    .Y(net283));
 NAND2x1_ASAP7_75t_R _20860_ (.A(net328),
    .B(_00742_),
    .Y(_15488_));
 OA211x2_ASAP7_75t_R _20861_ (.A1(net328),
    .A2(_15485_),
    .B(_15488_),
    .C(_00246_),
    .Y(_15489_));
 BUFx16f_ASAP7_75t_R load_slew282 (.A(_07162_),
    .Y(net282));
 BUFx12f_ASAP7_75t_R max_cap281 (.A(_06953_),
    .Y(net281));
 BUFx6f_ASAP7_75t_R load_slew280 (.A(\ex_block_i.alu_adder_result_ex_o[0] ),
    .Y(net280));
 AND2x2_ASAP7_75t_R _20865_ (.A(net328),
    .B(_00743_),
    .Y(_15493_));
 AO21x1_ASAP7_75t_R _20866_ (.A1(net312),
    .A2(_00745_),
    .B(_15493_),
    .Y(_15494_));
 BUFx4f_ASAP7_75t_R load_slew279 (.A(\ex_block_i.alu_adder_result_ex_o[1] ),
    .Y(net279));
 OAI21x1_ASAP7_75t_R _20868_ (.A1(_00246_),
    .A2(_15494_),
    .B(net322),
    .Y(_15496_));
 INVx1_ASAP7_75t_R _20869_ (.A(_00749_),
    .Y(_15497_));
 NAND2x1_ASAP7_75t_R _20870_ (.A(net328),
    .B(_00747_),
    .Y(_15498_));
 OA211x2_ASAP7_75t_R _20871_ (.A1(net328),
    .A2(_15497_),
    .B(_15498_),
    .C(net311),
    .Y(_15499_));
 INVx1_ASAP7_75t_R _20872_ (.A(_00748_),
    .Y(_15500_));
 NAND2x1_ASAP7_75t_R _20873_ (.A(net328),
    .B(_00746_),
    .Y(_15501_));
 OA211x2_ASAP7_75t_R _20874_ (.A1(net328),
    .A2(_15500_),
    .B(_15501_),
    .C(_00246_),
    .Y(_15502_));
 OR3x1_ASAP7_75t_R _20875_ (.A(net322),
    .B(_15499_),
    .C(_15502_),
    .Y(_15503_));
 BUFx6f_ASAP7_75t_R load_slew278 (.A(_17340_),
    .Y(net278));
 OA211x2_ASAP7_75t_R _20877_ (.A1(_15489_),
    .A2(_15496_),
    .B(_15503_),
    .C(_13598_),
    .Y(_15505_));
 OA21x2_ASAP7_75t_R _20878_ (.A1(_15482_),
    .A2(_15505_),
    .B(_13174_),
    .Y(_15506_));
 NOR2x2_ASAP7_75t_R _20879_ (.A(_15462_),
    .B(_15506_),
    .Y(_15507_));
 OA21x2_ASAP7_75t_R _20880_ (.A1(_00279_),
    .A2(_15268_),
    .B(_15269_),
    .Y(_15508_));
 AOI21x1_ASAP7_75t_R _20881_ (.A1(_13583_),
    .A2(_15507_),
    .B(_15508_),
    .Y(_18177_));
 NAND2x1_ASAP7_75t_R _20882_ (.A(net380),
    .B(_00735_),
    .Y(_15509_));
 OA211x2_ASAP7_75t_R _20883_ (.A1(net380),
    .A2(_15475_),
    .B(_15509_),
    .C(net305),
    .Y(_15510_));
 NAND2x1_ASAP7_75t_R _20884_ (.A(net380),
    .B(_00734_),
    .Y(_15511_));
 OA211x2_ASAP7_75t_R _20885_ (.A1(net380),
    .A2(_15478_),
    .B(_15511_),
    .C(net406),
    .Y(_15512_));
 OR3x1_ASAP7_75t_R _20886_ (.A(_13397_),
    .B(_15510_),
    .C(_15512_),
    .Y(_15513_));
 NAND2x1_ASAP7_75t_R _20887_ (.A(net376),
    .B(_00739_),
    .Y(_15514_));
 OA211x2_ASAP7_75t_R _20888_ (.A1(net376),
    .A2(_15465_),
    .B(_15514_),
    .C(net305),
    .Y(_15515_));
 NAND2x1_ASAP7_75t_R _20889_ (.A(net376),
    .B(_00738_),
    .Y(_15516_));
 OA211x2_ASAP7_75t_R _20890_ (.A1(net376),
    .A2(_15469_),
    .B(_15516_),
    .C(net406),
    .Y(_15517_));
 OR3x1_ASAP7_75t_R _20891_ (.A(net375),
    .B(_15515_),
    .C(_15517_),
    .Y(_15518_));
 BUFx12f_ASAP7_75t_R load_slew277 (.A(_02537_),
    .Y(net277));
 NAND2x1_ASAP7_75t_R _20893_ (.A(net377),
    .B(_00723_),
    .Y(_15520_));
 OA211x2_ASAP7_75t_R _20894_ (.A1(net377),
    .A2(_15444_),
    .B(_15520_),
    .C(net305),
    .Y(_15521_));
 NAND2x1_ASAP7_75t_R _20895_ (.A(net377),
    .B(_00722_),
    .Y(_15522_));
 OA211x2_ASAP7_75t_R _20896_ (.A1(net377),
    .A2(_15448_),
    .B(_15522_),
    .C(net412),
    .Y(_15523_));
 OR3x1_ASAP7_75t_R _20897_ (.A(net298),
    .B(_15521_),
    .C(_15523_),
    .Y(_15524_));
 NAND2x1_ASAP7_75t_R _20898_ (.A(net376),
    .B(_01695_),
    .Y(_15525_));
 OA211x2_ASAP7_75t_R _20899_ (.A1(net376),
    .A2(_15435_),
    .B(_15525_),
    .C(net305),
    .Y(_15526_));
 AND3x1_ASAP7_75t_R _20900_ (.A(net406),
    .B(net303),
    .C(_15434_),
    .Y(_15527_));
 OA31x2_ASAP7_75t_R _20901_ (.A1(net301),
    .A2(_15526_),
    .A3(_15527_),
    .B1(_00286_),
    .Y(_15528_));
 AO32x1_ASAP7_75t_R _20902_ (.A1(_13392_),
    .A2(_15513_),
    .A3(_15518_),
    .B1(_15524_),
    .B2(_15528_),
    .Y(_15529_));
 NAND2x1_ASAP7_75t_R _20903_ (.A(net377),
    .B(_00727_),
    .Y(_15530_));
 OA211x2_ASAP7_75t_R _20904_ (.A1(net377),
    .A2(_15421_),
    .B(_15530_),
    .C(net305),
    .Y(_15531_));
 NAND2x1_ASAP7_75t_R _20905_ (.A(net377),
    .B(_00726_),
    .Y(_15532_));
 OA211x2_ASAP7_75t_R _20906_ (.A1(net377),
    .A2(_15428_),
    .B(_15532_),
    .C(net412),
    .Y(_15533_));
 OR3x1_ASAP7_75t_R _20907_ (.A(_13397_),
    .B(_15531_),
    .C(_15533_),
    .Y(_15534_));
 NAND2x1_ASAP7_75t_R _20908_ (.A(net377),
    .B(_00731_),
    .Y(_15535_));
 OA211x2_ASAP7_75t_R _20909_ (.A1(net377),
    .A2(_15453_),
    .B(_15535_),
    .C(net305),
    .Y(_15536_));
 NAND2x1_ASAP7_75t_R _20910_ (.A(net377),
    .B(_00730_),
    .Y(_15537_));
 OA211x2_ASAP7_75t_R _20911_ (.A1(net377),
    .A2(_15456_),
    .B(_15537_),
    .C(net412),
    .Y(_15538_));
 OR3x1_ASAP7_75t_R _20912_ (.A(net375),
    .B(_15536_),
    .C(_15538_),
    .Y(_15539_));
 AND2x2_ASAP7_75t_R _20913_ (.A(_15534_),
    .B(_15539_),
    .Y(_15540_));
 AND2x2_ASAP7_75t_R _20914_ (.A(_15524_),
    .B(_15528_),
    .Y(_15541_));
 NAND2x1_ASAP7_75t_R _20915_ (.A(net375),
    .B(_00745_),
    .Y(_15542_));
 OA211x2_ASAP7_75t_R _20916_ (.A1(net375),
    .A2(_15497_),
    .B(_15542_),
    .C(net305),
    .Y(_15543_));
 NAND2x1_ASAP7_75t_R _20917_ (.A(net375),
    .B(_00744_),
    .Y(_15544_));
 OA211x2_ASAP7_75t_R _20918_ (.A1(net375),
    .A2(_15500_),
    .B(_15544_),
    .C(net406),
    .Y(_15545_));
 OR3x1_ASAP7_75t_R _20919_ (.A(net376),
    .B(_15543_),
    .C(_15545_),
    .Y(_15546_));
 INVx1_ASAP7_75t_R _20920_ (.A(_00747_),
    .Y(_15547_));
 NAND2x1_ASAP7_75t_R _20921_ (.A(net375),
    .B(_00743_),
    .Y(_15548_));
 OA211x2_ASAP7_75t_R _20922_ (.A1(net375),
    .A2(_15547_),
    .B(_15548_),
    .C(net305),
    .Y(_15549_));
 INVx1_ASAP7_75t_R _20923_ (.A(_00746_),
    .Y(_15550_));
 NAND2x1_ASAP7_75t_R _20924_ (.A(net375),
    .B(_00742_),
    .Y(_15551_));
 OA211x2_ASAP7_75t_R _20925_ (.A1(net375),
    .A2(_15550_),
    .B(_15551_),
    .C(net406),
    .Y(_15552_));
 OR3x1_ASAP7_75t_R _20926_ (.A(net303),
    .B(_15549_),
    .C(_15552_),
    .Y(_15553_));
 AND3x1_ASAP7_75t_R _20927_ (.A(_14571_),
    .B(_15546_),
    .C(_15553_),
    .Y(_15554_));
 AOI221x1_ASAP7_75t_R _20928_ (.A1(net368),
    .A2(_15529_),
    .B1(_15540_),
    .B2(_15541_),
    .C(_15554_),
    .Y(_15555_));
 OA222x2_ASAP7_75t_R _20929_ (.A1(_01627_),
    .A2(_13223_),
    .B1(_13782_),
    .B2(_15555_),
    .C1(_13880_),
    .C2(_00204_),
    .Y(_15556_));
 BUFx12f_ASAP7_75t_R load_slew276 (.A(_00231_),
    .Y(net276));
 XOR2x2_ASAP7_75t_R _20931_ (.A(_00751_),
    .B(_02227_),
    .Y(_15557_));
 CKINVDCx5p33_ASAP7_75t_R _20932_ (.A(_15557_),
    .Y(net155));
 AND2x2_ASAP7_75t_R _20933_ (.A(net345),
    .B(_01694_),
    .Y(_15558_));
 AO21x1_ASAP7_75t_R _20934_ (.A1(net312),
    .A2(_00754_),
    .B(_15558_),
    .Y(_15559_));
 OAI22x1_ASAP7_75t_R _20935_ (.A1(_00753_),
    .A2(_13586_),
    .B1(_15559_),
    .B2(net355),
    .Y(_15560_));
 INVx1_ASAP7_75t_R _20936_ (.A(_00762_),
    .Y(_15561_));
 NAND2x1_ASAP7_75t_R _20937_ (.A(net345),
    .B(_00760_),
    .Y(_15562_));
 OA211x2_ASAP7_75t_R _20938_ (.A1(net345),
    .A2(_15561_),
    .B(_15562_),
    .C(net310),
    .Y(_15563_));
 INVx1_ASAP7_75t_R _20939_ (.A(_00761_),
    .Y(_15564_));
 NAND2x1_ASAP7_75t_R _20940_ (.A(net345),
    .B(_00759_),
    .Y(_15565_));
 OA211x2_ASAP7_75t_R _20941_ (.A1(net345),
    .A2(_15564_),
    .B(_15565_),
    .C(net355),
    .Y(_15566_));
 OR3x1_ASAP7_75t_R _20942_ (.A(net318),
    .B(_15563_),
    .C(_15566_),
    .Y(_15567_));
 OA21x2_ASAP7_75t_R _20943_ (.A1(_13598_),
    .A2(_15560_),
    .B(_15567_),
    .Y(_15568_));
 INVx1_ASAP7_75t_R _20944_ (.A(_00758_),
    .Y(_15569_));
 NAND2x1_ASAP7_75t_R _20945_ (.A(net345),
    .B(_00756_),
    .Y(_15570_));
 OA211x2_ASAP7_75t_R _20946_ (.A1(net345),
    .A2(_15569_),
    .B(_15570_),
    .C(net310),
    .Y(_15571_));
 BUFx6f_ASAP7_75t_R load_slew275 (.A(net174),
    .Y(net275));
 INVx1_ASAP7_75t_R _20948_ (.A(_00757_),
    .Y(_15573_));
 NAND2x1_ASAP7_75t_R _20949_ (.A(net345),
    .B(_00755_),
    .Y(_15574_));
 OA211x2_ASAP7_75t_R _20950_ (.A1(net345),
    .A2(_15573_),
    .B(_15574_),
    .C(net355),
    .Y(_15575_));
 OR3x1_ASAP7_75t_R _20951_ (.A(_13598_),
    .B(_15571_),
    .C(_15575_),
    .Y(_15576_));
 INVx1_ASAP7_75t_R _20952_ (.A(_00766_),
    .Y(_15577_));
 NAND2x1_ASAP7_75t_R _20953_ (.A(net345),
    .B(_00764_),
    .Y(_15578_));
 OA211x2_ASAP7_75t_R _20954_ (.A1(net345),
    .A2(_15577_),
    .B(_15578_),
    .C(net310),
    .Y(_15579_));
 INVx1_ASAP7_75t_R _20955_ (.A(_00765_),
    .Y(_15580_));
 NAND2x1_ASAP7_75t_R _20956_ (.A(net345),
    .B(_00763_),
    .Y(_15581_));
 OA211x2_ASAP7_75t_R _20957_ (.A1(net345),
    .A2(_15580_),
    .B(_15581_),
    .C(net355),
    .Y(_15582_));
 OR3x1_ASAP7_75t_R _20958_ (.A(net318),
    .B(_15579_),
    .C(_15582_),
    .Y(_15583_));
 AND3x1_ASAP7_75t_R _20959_ (.A(_13132_),
    .B(_15576_),
    .C(_15583_),
    .Y(_15584_));
 AO21x1_ASAP7_75t_R _20960_ (.A1(net324),
    .A2(_15568_),
    .B(_15584_),
    .Y(_15585_));
 INVx1_ASAP7_75t_R _20961_ (.A(_00770_),
    .Y(_15586_));
 NAND2x1_ASAP7_75t_R _20962_ (.A(net344),
    .B(_00768_),
    .Y(_15587_));
 OA211x2_ASAP7_75t_R _20963_ (.A1(net344),
    .A2(_15586_),
    .B(_15587_),
    .C(net310),
    .Y(_15588_));
 INVx1_ASAP7_75t_R _20964_ (.A(_00769_),
    .Y(_15589_));
 NAND2x1_ASAP7_75t_R _20965_ (.A(net344),
    .B(_00767_),
    .Y(_15590_));
 OA211x2_ASAP7_75t_R _20966_ (.A1(net344),
    .A2(_15589_),
    .B(_15590_),
    .C(net355),
    .Y(_15591_));
 OR3x1_ASAP7_75t_R _20967_ (.A(_13132_),
    .B(_15588_),
    .C(_15591_),
    .Y(_15592_));
 INVx1_ASAP7_75t_R _20968_ (.A(_00774_),
    .Y(_15593_));
 NAND2x1_ASAP7_75t_R _20969_ (.A(net344),
    .B(_00772_),
    .Y(_15594_));
 OA211x2_ASAP7_75t_R _20970_ (.A1(net344),
    .A2(_15593_),
    .B(_15594_),
    .C(net310),
    .Y(_15595_));
 INVx1_ASAP7_75t_R _20971_ (.A(_00773_),
    .Y(_15596_));
 NAND2x1_ASAP7_75t_R _20972_ (.A(net344),
    .B(_00771_),
    .Y(_15597_));
 OA211x2_ASAP7_75t_R _20973_ (.A1(net344),
    .A2(_15596_),
    .B(_15597_),
    .C(net355),
    .Y(_15598_));
 OR3x1_ASAP7_75t_R _20974_ (.A(net324),
    .B(_15595_),
    .C(_15598_),
    .Y(_15599_));
 AND3x1_ASAP7_75t_R _20975_ (.A(net318),
    .B(_15592_),
    .C(_15599_),
    .Y(_15600_));
 INVx1_ASAP7_75t_R _20976_ (.A(_00782_),
    .Y(_15601_));
 NAND2x1_ASAP7_75t_R _20977_ (.A(net344),
    .B(_00780_),
    .Y(_15602_));
 OA211x2_ASAP7_75t_R _20978_ (.A1(net344),
    .A2(_15601_),
    .B(_15602_),
    .C(_13145_),
    .Y(_15603_));
 INVx1_ASAP7_75t_R _20979_ (.A(_00781_),
    .Y(_15604_));
 NAND2x1_ASAP7_75t_R _20980_ (.A(net344),
    .B(_00779_),
    .Y(_15605_));
 OA211x2_ASAP7_75t_R _20981_ (.A1(net344),
    .A2(_15604_),
    .B(_15605_),
    .C(net355),
    .Y(_15606_));
 OR3x1_ASAP7_75t_R _20982_ (.A(net324),
    .B(_15603_),
    .C(_15606_),
    .Y(_15607_));
 INVx1_ASAP7_75t_R _20983_ (.A(_00778_),
    .Y(_15608_));
 NAND2x1_ASAP7_75t_R _20984_ (.A(net344),
    .B(_00776_),
    .Y(_15609_));
 OA211x2_ASAP7_75t_R _20985_ (.A1(net344),
    .A2(_15608_),
    .B(_15609_),
    .C(_13145_),
    .Y(_15610_));
 INVx1_ASAP7_75t_R _20986_ (.A(_00777_),
    .Y(_15611_));
 NAND2x1_ASAP7_75t_R _20987_ (.A(net344),
    .B(_00775_),
    .Y(_15612_));
 OA211x2_ASAP7_75t_R _20988_ (.A1(net344),
    .A2(_15611_),
    .B(_15612_),
    .C(net355),
    .Y(_15613_));
 OR3x1_ASAP7_75t_R _20989_ (.A(_13132_),
    .B(_15610_),
    .C(_15613_),
    .Y(_15614_));
 AND3x1_ASAP7_75t_R _20990_ (.A(_13598_),
    .B(_15607_),
    .C(_15614_),
    .Y(_15615_));
 OR3x1_ASAP7_75t_R _20991_ (.A(net315),
    .B(_15600_),
    .C(_15615_),
    .Y(_15616_));
 OA21x2_ASAP7_75t_R _20992_ (.A1(_13174_),
    .A2(_15585_),
    .B(_15616_),
    .Y(_15617_));
 INVx1_ASAP7_75t_R _20993_ (.A(_15617_),
    .Y(_15618_));
 OA21x2_ASAP7_75t_R _20994_ (.A1(_00290_),
    .A2(_15268_),
    .B(_15269_),
    .Y(_15619_));
 AO21x2_ASAP7_75t_R _20995_ (.A1(_13583_),
    .A2(_15618_),
    .B(_15619_),
    .Y(_15620_));
 BUFx10_ASAP7_75t_R max_cap274 (.A(_18337_),
    .Y(net274));
 INVx1_ASAP7_75t_R _20997_ (.A(_15620_),
    .Y(_18181_));
 INVx1_ASAP7_75t_R _20998_ (.A(_00206_),
    .Y(\cs_registers_i.pc_id_i[15] ));
 INVx1_ASAP7_75t_R _20999_ (.A(_01626_),
    .Y(_15621_));
 NAND2x1_ASAP7_75t_R _21000_ (.A(net388),
    .B(_00756_),
    .Y(_15622_));
 OA211x2_ASAP7_75t_R _21001_ (.A1(net388),
    .A2(_15569_),
    .B(_15622_),
    .C(net307),
    .Y(_15623_));
 NAND2x1_ASAP7_75t_R _21002_ (.A(net388),
    .B(_00755_),
    .Y(_15624_));
 OA211x2_ASAP7_75t_R _21003_ (.A1(net388),
    .A2(_15573_),
    .B(_15624_),
    .C(net407),
    .Y(_15625_));
 OR3x1_ASAP7_75t_R _21004_ (.A(_13484_),
    .B(_15623_),
    .C(_15625_),
    .Y(_15626_));
 NAND2x1_ASAP7_75t_R _21005_ (.A(net388),
    .B(_00764_),
    .Y(_15627_));
 OA211x2_ASAP7_75t_R _21006_ (.A1(net388),
    .A2(_15577_),
    .B(_15627_),
    .C(net307),
    .Y(_15628_));
 NAND2x1_ASAP7_75t_R _21007_ (.A(net388),
    .B(_00763_),
    .Y(_15629_));
 OA211x2_ASAP7_75t_R _21008_ (.A1(net388),
    .A2(_15580_),
    .B(_15629_),
    .C(net407),
    .Y(_15630_));
 OR3x1_ASAP7_75t_R _21009_ (.A(net366),
    .B(_15628_),
    .C(_15630_),
    .Y(_15631_));
 AO21x1_ASAP7_75t_R _21010_ (.A1(_15626_),
    .A2(_15631_),
    .B(net370),
    .Y(_15632_));
 BUFx6f_ASAP7_75t_R max_cap273 (.A(net274),
    .Y(net273));
 NAND2x1_ASAP7_75t_R _21012_ (.A(net392),
    .B(_00760_),
    .Y(_15634_));
 OA211x2_ASAP7_75t_R _21013_ (.A1(net392),
    .A2(_15561_),
    .B(_15634_),
    .C(net307),
    .Y(_15635_));
 NAND2x1_ASAP7_75t_R _21014_ (.A(net392),
    .B(_00759_),
    .Y(_15636_));
 OA211x2_ASAP7_75t_R _21015_ (.A1(net392),
    .A2(_15564_),
    .B(_15636_),
    .C(net407),
    .Y(_15637_));
 OR3x1_ASAP7_75t_R _21016_ (.A(_14743_),
    .B(_15635_),
    .C(_15637_),
    .Y(_15638_));
 AND2x2_ASAP7_75t_R _21017_ (.A(net392),
    .B(_01694_),
    .Y(_15639_));
 AO21x1_ASAP7_75t_R _21018_ (.A1(net303),
    .A2(_00754_),
    .B(_15639_),
    .Y(_15640_));
 OAI22x1_ASAP7_75t_R _21019_ (.A1(_00753_),
    .A2(_13471_),
    .B1(_15640_),
    .B2(net407),
    .Y(_15641_));
 OA21x2_ASAP7_75t_R _21020_ (.A1(net301),
    .A2(_15641_),
    .B(net363),
    .Y(_15642_));
 NAND2x1_ASAP7_75t_R _21021_ (.A(net389),
    .B(_00776_),
    .Y(_15643_));
 OA211x2_ASAP7_75t_R _21022_ (.A1(net389),
    .A2(_15608_),
    .B(_15643_),
    .C(_13424_),
    .Y(_15644_));
 NAND2x1_ASAP7_75t_R _21023_ (.A(net389),
    .B(_00775_),
    .Y(_15645_));
 OA211x2_ASAP7_75t_R _21024_ (.A1(net389),
    .A2(_15611_),
    .B(_15645_),
    .C(net407),
    .Y(_15646_));
 OR3x1_ASAP7_75t_R _21025_ (.A(_13397_),
    .B(_15644_),
    .C(_15646_),
    .Y(_15647_));
 NAND2x1_ASAP7_75t_R _21026_ (.A(net388),
    .B(_00780_),
    .Y(_15648_));
 OA211x2_ASAP7_75t_R _21027_ (.A1(net388),
    .A2(_15601_),
    .B(_15648_),
    .C(_13424_),
    .Y(_15649_));
 NAND2x1_ASAP7_75t_R _21028_ (.A(net388),
    .B(_00779_),
    .Y(_15650_));
 OA211x2_ASAP7_75t_R _21029_ (.A1(net388),
    .A2(_15604_),
    .B(_15650_),
    .C(net407),
    .Y(_15651_));
 OR3x1_ASAP7_75t_R _21030_ (.A(net370),
    .B(_15649_),
    .C(_15651_),
    .Y(_15652_));
 AO21x1_ASAP7_75t_R _21031_ (.A1(_15647_),
    .A2(_15652_),
    .B(net366),
    .Y(_15653_));
 NAND2x1_ASAP7_75t_R _21032_ (.A(net388),
    .B(_00772_),
    .Y(_15654_));
 OA211x2_ASAP7_75t_R _21033_ (.A1(net388),
    .A2(_15593_),
    .B(_15654_),
    .C(net307),
    .Y(_15655_));
 NAND2x1_ASAP7_75t_R _21034_ (.A(net388),
    .B(_00771_),
    .Y(_15656_));
 OA211x2_ASAP7_75t_R _21035_ (.A1(net388),
    .A2(_15596_),
    .B(_15656_),
    .C(net407),
    .Y(_15657_));
 OR3x1_ASAP7_75t_R _21036_ (.A(_13814_),
    .B(_15655_),
    .C(_15657_),
    .Y(_15658_));
 NAND2x1_ASAP7_75t_R _21037_ (.A(net388),
    .B(_00767_),
    .Y(_15659_));
 OA211x2_ASAP7_75t_R _21038_ (.A1(net388),
    .A2(_15589_),
    .B(_15659_),
    .C(net407),
    .Y(_15660_));
 NAND2x1_ASAP7_75t_R _21039_ (.A(net388),
    .B(_00768_),
    .Y(_15661_));
 OA211x2_ASAP7_75t_R _21040_ (.A1(net388),
    .A2(_15586_),
    .B(_15661_),
    .C(net306),
    .Y(_15662_));
 OR3x1_ASAP7_75t_R _21041_ (.A(_13828_),
    .B(_15660_),
    .C(_15662_),
    .Y(_15663_));
 AND3x1_ASAP7_75t_R _21042_ (.A(_13392_),
    .B(_15658_),
    .C(_15663_),
    .Y(_15664_));
 AO32x2_ASAP7_75t_R _21043_ (.A1(_15632_),
    .A2(_15638_),
    .A3(_15642_),
    .B1(_15653_),
    .B2(_15664_),
    .Y(_15665_));
 NAND2x1_ASAP7_75t_R _21044_ (.A(_00206_),
    .B(_13553_),
    .Y(_15666_));
 OA211x2_ASAP7_75t_R _21045_ (.A1(_13553_),
    .A2(_15665_),
    .B(_15666_),
    .C(_14757_),
    .Y(_15667_));
 AO21x2_ASAP7_75t_R _21046_ (.A1(_15621_),
    .A2(_13270_),
    .B(_15667_),
    .Y(_15668_));
 BUFx16f_ASAP7_75t_R wire272 (.A(_12042_),
    .Y(net272));
 INVx2_ASAP7_75t_R _21048_ (.A(_15668_),
    .Y(_18182_));
 AO21x1_ASAP7_75t_R _21049_ (.A1(_15413_),
    .A2(_15417_),
    .B(_00719_),
    .Y(_15669_));
 AO21x1_ASAP7_75t_R _21050_ (.A1(_00752_),
    .A2(_15669_),
    .B(_00751_),
    .Y(_15670_));
 NAND2x1_ASAP7_75t_R _21051_ (.A(_02273_),
    .B(_15670_),
    .Y(_16523_));
 INVx3_ASAP7_75t_R _21052_ (.A(_00785_),
    .Y(net156));
 BUFx10_ASAP7_75t_R max_cap271 (.A(_12042_),
    .Y(net271));
 AND2x2_ASAP7_75t_R _21054_ (.A(net334),
    .B(_01693_),
    .Y(_15672_));
 AO21x1_ASAP7_75t_R _21055_ (.A1(net313),
    .A2(_00787_),
    .B(_15672_),
    .Y(_15673_));
 OAI22x1_ASAP7_75t_R _21056_ (.A1(_00786_),
    .A2(_13586_),
    .B1(_15673_),
    .B2(net357),
    .Y(_15674_));
 INVx1_ASAP7_75t_R _21057_ (.A(_00795_),
    .Y(_15675_));
 NAND2x1_ASAP7_75t_R _21058_ (.A(net335),
    .B(_00793_),
    .Y(_15676_));
 OA211x2_ASAP7_75t_R _21059_ (.A1(net335),
    .A2(_15675_),
    .B(_15676_),
    .C(net308),
    .Y(_15677_));
 INVx1_ASAP7_75t_R _21060_ (.A(_00794_),
    .Y(_15678_));
 NAND2x1_ASAP7_75t_R _21061_ (.A(net334),
    .B(_00792_),
    .Y(_15679_));
 OA211x2_ASAP7_75t_R _21062_ (.A1(net334),
    .A2(_15678_),
    .B(_15679_),
    .C(net357),
    .Y(_15680_));
 OR3x1_ASAP7_75t_R _21063_ (.A(net319),
    .B(_15677_),
    .C(_15680_),
    .Y(_15681_));
 OA211x2_ASAP7_75t_R _21064_ (.A1(_13598_),
    .A2(_15674_),
    .B(_15681_),
    .C(net324),
    .Y(_15682_));
 BUFx16f_ASAP7_75t_R load_slew270 (.A(_09780_),
    .Y(net270));
 INVx1_ASAP7_75t_R _21066_ (.A(_00791_),
    .Y(_15684_));
 NAND2x1_ASAP7_75t_R _21067_ (.A(net335),
    .B(_00789_),
    .Y(_15685_));
 OA211x2_ASAP7_75t_R _21068_ (.A1(net335),
    .A2(_15684_),
    .B(_15685_),
    .C(net308),
    .Y(_15686_));
 INVx1_ASAP7_75t_R _21069_ (.A(_00790_),
    .Y(_15687_));
 NAND2x1_ASAP7_75t_R _21070_ (.A(net335),
    .B(_00788_),
    .Y(_15688_));
 OA211x2_ASAP7_75t_R _21071_ (.A1(net335),
    .A2(_15687_),
    .B(_15688_),
    .C(net357),
    .Y(_15689_));
 OR3x1_ASAP7_75t_R _21072_ (.A(_13598_),
    .B(_15686_),
    .C(_15689_),
    .Y(_15690_));
 INVx1_ASAP7_75t_R _21073_ (.A(_00799_),
    .Y(_15691_));
 NAND2x1_ASAP7_75t_R _21074_ (.A(net335),
    .B(_00797_),
    .Y(_15692_));
 OA211x2_ASAP7_75t_R _21075_ (.A1(net335),
    .A2(_15691_),
    .B(_15692_),
    .C(net309),
    .Y(_15693_));
 INVx1_ASAP7_75t_R _21076_ (.A(_00798_),
    .Y(_15694_));
 NAND2x1_ASAP7_75t_R _21077_ (.A(net335),
    .B(_00796_),
    .Y(_15695_));
 OA211x2_ASAP7_75t_R _21078_ (.A1(net335),
    .A2(_15694_),
    .B(_15695_),
    .C(net356),
    .Y(_15696_));
 OR3x1_ASAP7_75t_R _21079_ (.A(net319),
    .B(_15693_),
    .C(_15696_),
    .Y(_15697_));
 AND3x1_ASAP7_75t_R _21080_ (.A(_13132_),
    .B(_15690_),
    .C(_15697_),
    .Y(_15698_));
 OR3x2_ASAP7_75t_R _21081_ (.A(_13174_),
    .B(_15682_),
    .C(_15698_),
    .Y(_15699_));
 INVx1_ASAP7_75t_R _21082_ (.A(_00807_),
    .Y(_15700_));
 NAND2x1_ASAP7_75t_R _21083_ (.A(net335),
    .B(_00805_),
    .Y(_15701_));
 OA211x2_ASAP7_75t_R _21084_ (.A1(net335),
    .A2(_15700_),
    .B(_15701_),
    .C(net308),
    .Y(_15702_));
 INVx1_ASAP7_75t_R _21085_ (.A(_00806_),
    .Y(_15703_));
 NAND2x1_ASAP7_75t_R _21086_ (.A(net335),
    .B(_00804_),
    .Y(_15704_));
 OA211x2_ASAP7_75t_R _21087_ (.A1(net335),
    .A2(_15703_),
    .B(_15704_),
    .C(net357),
    .Y(_15705_));
 OR3x1_ASAP7_75t_R _21088_ (.A(_13598_),
    .B(_15702_),
    .C(_15705_),
    .Y(_15706_));
 INVx1_ASAP7_75t_R _21089_ (.A(_00815_),
    .Y(_15707_));
 NAND2x1_ASAP7_75t_R _21090_ (.A(net335),
    .B(_00813_),
    .Y(_15708_));
 OA211x2_ASAP7_75t_R _21091_ (.A1(net335),
    .A2(_15707_),
    .B(_15708_),
    .C(net308),
    .Y(_15709_));
 INVx1_ASAP7_75t_R _21092_ (.A(_00814_),
    .Y(_15710_));
 NAND2x1_ASAP7_75t_R _21093_ (.A(net335),
    .B(_00812_),
    .Y(_15711_));
 OA211x2_ASAP7_75t_R _21094_ (.A1(net335),
    .A2(_15710_),
    .B(_15711_),
    .C(net356),
    .Y(_15712_));
 OR3x1_ASAP7_75t_R _21095_ (.A(net319),
    .B(_15709_),
    .C(_15712_),
    .Y(_15713_));
 AND3x1_ASAP7_75t_R _21096_ (.A(_13132_),
    .B(_15706_),
    .C(_15713_),
    .Y(_15714_));
 INVx1_ASAP7_75t_R _21097_ (.A(_00803_),
    .Y(_15715_));
 NAND2x1_ASAP7_75t_R _21098_ (.A(net335),
    .B(_00801_),
    .Y(_15716_));
 OA211x2_ASAP7_75t_R _21099_ (.A1(net335),
    .A2(_15715_),
    .B(_15716_),
    .C(net308),
    .Y(_15717_));
 INVx1_ASAP7_75t_R _21100_ (.A(_00802_),
    .Y(_15718_));
 NAND2x1_ASAP7_75t_R _21101_ (.A(net335),
    .B(_00800_),
    .Y(_15719_));
 OA211x2_ASAP7_75t_R _21102_ (.A1(net335),
    .A2(_15718_),
    .B(_15719_),
    .C(net357),
    .Y(_15720_));
 OR3x1_ASAP7_75t_R _21103_ (.A(_13598_),
    .B(_15717_),
    .C(_15720_),
    .Y(_15721_));
 INVx1_ASAP7_75t_R _21104_ (.A(_00811_),
    .Y(_15722_));
 NAND2x1_ASAP7_75t_R _21105_ (.A(net335),
    .B(_00809_),
    .Y(_15723_));
 OA211x2_ASAP7_75t_R _21106_ (.A1(net335),
    .A2(_15722_),
    .B(_15723_),
    .C(net308),
    .Y(_15724_));
 INVx1_ASAP7_75t_R _21107_ (.A(_00810_),
    .Y(_15725_));
 NAND2x1_ASAP7_75t_R _21108_ (.A(net334),
    .B(_00808_),
    .Y(_15726_));
 OA211x2_ASAP7_75t_R _21109_ (.A1(net334),
    .A2(_15725_),
    .B(_15726_),
    .C(net357),
    .Y(_15727_));
 OR3x1_ASAP7_75t_R _21110_ (.A(net319),
    .B(_15724_),
    .C(_15727_),
    .Y(_15728_));
 AND3x1_ASAP7_75t_R _21111_ (.A(net324),
    .B(_15721_),
    .C(_15728_),
    .Y(_15729_));
 OR3x4_ASAP7_75t_R _21112_ (.A(net314),
    .B(_15714_),
    .C(_15729_),
    .Y(_15730_));
 NAND2x2_ASAP7_75t_R _21113_ (.A(_15699_),
    .B(_15730_),
    .Y(_15731_));
 OA21x2_ASAP7_75t_R _21114_ (.A1(net398),
    .A2(_15268_),
    .B(_15269_),
    .Y(_15732_));
 AOI21x1_ASAP7_75t_R _21115_ (.A1(_13583_),
    .A2(_15731_),
    .B(_15732_),
    .Y(_18187_));
 INVx1_ASAP7_75t_R _21116_ (.A(_01625_),
    .Y(_15733_));
 AND2x2_ASAP7_75t_R _21117_ (.A(net394),
    .B(_01693_),
    .Y(_15734_));
 AO21x1_ASAP7_75t_R _21118_ (.A1(net302),
    .A2(_00787_),
    .B(_15734_),
    .Y(_15735_));
 OAI22x1_ASAP7_75t_R _21119_ (.A1(_00786_),
    .A2(_13471_),
    .B1(_15735_),
    .B2(net409),
    .Y(_15736_));
 NAND2x1_ASAP7_75t_R _21120_ (.A(net392),
    .B(_00801_),
    .Y(_15737_));
 OA211x2_ASAP7_75t_R _21121_ (.A1(net392),
    .A2(_15715_),
    .B(_15737_),
    .C(net306),
    .Y(_15738_));
 NAND2x1_ASAP7_75t_R _21122_ (.A(net392),
    .B(_00800_),
    .Y(_15739_));
 OA211x2_ASAP7_75t_R _21123_ (.A1(net392),
    .A2(_15718_),
    .B(_15739_),
    .C(net409),
    .Y(_15740_));
 OR3x1_ASAP7_75t_R _21124_ (.A(net362),
    .B(_15738_),
    .C(_15740_),
    .Y(_15741_));
 OA211x2_ASAP7_75t_R _21125_ (.A1(_13392_),
    .A2(_15736_),
    .B(_15741_),
    .C(net372),
    .Y(_15742_));
 NAND2x1_ASAP7_75t_R _21126_ (.A(net400),
    .B(_00789_),
    .Y(_15743_));
 OA211x2_ASAP7_75t_R _21127_ (.A1(net400),
    .A2(_15684_),
    .B(_15743_),
    .C(net306),
    .Y(_15744_));
 NAND2x1_ASAP7_75t_R _21128_ (.A(net400),
    .B(_00788_),
    .Y(_15745_));
 OA211x2_ASAP7_75t_R _21129_ (.A1(net400),
    .A2(_15687_),
    .B(_15745_),
    .C(net409),
    .Y(_15746_));
 OR3x1_ASAP7_75t_R _21130_ (.A(_13392_),
    .B(_15744_),
    .C(_15746_),
    .Y(_15747_));
 NAND2x1_ASAP7_75t_R _21131_ (.A(net392),
    .B(_00805_),
    .Y(_15748_));
 OA211x2_ASAP7_75t_R _21132_ (.A1(net392),
    .A2(_15700_),
    .B(_15748_),
    .C(net306),
    .Y(_15749_));
 NAND2x1_ASAP7_75t_R _21133_ (.A(net391),
    .B(_00804_),
    .Y(_15750_));
 OA211x2_ASAP7_75t_R _21134_ (.A1(net391),
    .A2(_15703_),
    .B(_15750_),
    .C(net409),
    .Y(_15751_));
 OR3x1_ASAP7_75t_R _21135_ (.A(net362),
    .B(_15749_),
    .C(_15751_),
    .Y(_15752_));
 AND3x1_ASAP7_75t_R _21136_ (.A(_13397_),
    .B(_15747_),
    .C(_15752_),
    .Y(_15753_));
 OR3x4_ASAP7_75t_R _21137_ (.A(_13484_),
    .B(_15742_),
    .C(_15753_),
    .Y(_15754_));
 NAND2x1_ASAP7_75t_R _21138_ (.A(net394),
    .B(_00793_),
    .Y(_15755_));
 OA211x2_ASAP7_75t_R _21139_ (.A1(net394),
    .A2(_15675_),
    .B(_15755_),
    .C(net362),
    .Y(_15756_));
 NAND2x1_ASAP7_75t_R _21140_ (.A(net394),
    .B(_00809_),
    .Y(_15757_));
 OA211x2_ASAP7_75t_R _21141_ (.A1(net394),
    .A2(_15722_),
    .B(_15757_),
    .C(_13392_),
    .Y(_15758_));
 OR3x1_ASAP7_75t_R _21142_ (.A(net409),
    .B(_15756_),
    .C(_15758_),
    .Y(_15759_));
 NAND2x1_ASAP7_75t_R _21143_ (.A(net394),
    .B(_00792_),
    .Y(_15760_));
 OA211x2_ASAP7_75t_R _21144_ (.A1(net394),
    .A2(_15678_),
    .B(_15760_),
    .C(net362),
    .Y(_15761_));
 NAND2x1_ASAP7_75t_R _21145_ (.A(net394),
    .B(_00808_),
    .Y(_15762_));
 OA211x2_ASAP7_75t_R _21146_ (.A1(net394),
    .A2(_15725_),
    .B(_15762_),
    .C(_13392_),
    .Y(_15763_));
 OR3x1_ASAP7_75t_R _21147_ (.A(net306),
    .B(_15761_),
    .C(_15763_),
    .Y(_15764_));
 AND3x1_ASAP7_75t_R _21148_ (.A(net372),
    .B(_15759_),
    .C(_15764_),
    .Y(_15765_));
 NAND2x1_ASAP7_75t_R _21149_ (.A(net392),
    .B(_00796_),
    .Y(_15766_));
 OA211x2_ASAP7_75t_R _21150_ (.A1(net392),
    .A2(_15694_),
    .B(_15766_),
    .C(net362),
    .Y(_15767_));
 NAND2x1_ASAP7_75t_R _21151_ (.A(net392),
    .B(_00812_),
    .Y(_15768_));
 OA211x2_ASAP7_75t_R _21152_ (.A1(net392),
    .A2(_15710_),
    .B(_15768_),
    .C(_13392_),
    .Y(_15769_));
 OR3x1_ASAP7_75t_R _21153_ (.A(net307),
    .B(_15767_),
    .C(_15769_),
    .Y(_15770_));
 NAND2x1_ASAP7_75t_R _21154_ (.A(net392),
    .B(_00797_),
    .Y(_15771_));
 OA211x2_ASAP7_75t_R _21155_ (.A1(net392),
    .A2(_15691_),
    .B(_15771_),
    .C(net362),
    .Y(_15772_));
 NAND2x1_ASAP7_75t_R _21156_ (.A(net392),
    .B(_00813_),
    .Y(_15773_));
 OA211x2_ASAP7_75t_R _21157_ (.A1(net392),
    .A2(_15707_),
    .B(_15773_),
    .C(_13392_),
    .Y(_15774_));
 OR3x1_ASAP7_75t_R _21158_ (.A(net409),
    .B(_15772_),
    .C(_15774_),
    .Y(_15775_));
 AND3x1_ASAP7_75t_R _21159_ (.A(_13397_),
    .B(_15770_),
    .C(_15775_),
    .Y(_15776_));
 OR3x4_ASAP7_75t_R _21160_ (.A(net365),
    .B(_15765_),
    .C(_15776_),
    .Y(_15777_));
 BUFx16f_ASAP7_75t_R load_slew269 (.A(net270),
    .Y(net269));
 NOR2x1_ASAP7_75t_R _21162_ (.A(_00208_),
    .B(_13879_),
    .Y(_15779_));
 AO31x2_ASAP7_75t_R _21163_ (.A1(_13879_),
    .A2(_15754_),
    .A3(_15777_),
    .B(_15779_),
    .Y(_15780_));
 AO22x2_ASAP7_75t_R _21164_ (.A1(_15733_),
    .A2(_13270_),
    .B1(_14757_),
    .B2(_15780_),
    .Y(_15781_));
 BUFx16f_ASAP7_75t_R load_slew268 (.A(_09941_),
    .Y(net268));
 INVx3_ASAP7_75t_R _21166_ (.A(_15781_),
    .Y(_18186_));
 INVx1_ASAP7_75t_R _21167_ (.A(_00843_),
    .Y(_15782_));
 NAND2x1_ASAP7_75t_R _21168_ (.A(net342),
    .B(_00841_),
    .Y(_15783_));
 OA211x2_ASAP7_75t_R _21169_ (.A1(net342),
    .A2(_15782_),
    .B(_15783_),
    .C(net356),
    .Y(_15784_));
 AND2x2_ASAP7_75t_R _21170_ (.A(net342),
    .B(_00842_),
    .Y(_15785_));
 AO21x1_ASAP7_75t_R _21171_ (.A1(net312),
    .A2(_00844_),
    .B(_15785_),
    .Y(_15786_));
 OAI21x1_ASAP7_75t_R _21172_ (.A1(net356),
    .A2(_15786_),
    .B(net323),
    .Y(_15787_));
 INVx1_ASAP7_75t_R _21173_ (.A(_00848_),
    .Y(_15788_));
 NAND2x1_ASAP7_75t_R _21174_ (.A(net342),
    .B(_00846_),
    .Y(_15789_));
 OA211x2_ASAP7_75t_R _21175_ (.A1(net342),
    .A2(_15788_),
    .B(_15789_),
    .C(net311),
    .Y(_15790_));
 INVx1_ASAP7_75t_R _21176_ (.A(_00847_),
    .Y(_15791_));
 NAND2x1_ASAP7_75t_R _21177_ (.A(net342),
    .B(_00845_),
    .Y(_15792_));
 OA211x2_ASAP7_75t_R _21178_ (.A1(net342),
    .A2(_15791_),
    .B(_15792_),
    .C(net356),
    .Y(_15793_));
 OR3x1_ASAP7_75t_R _21179_ (.A(net323),
    .B(_15790_),
    .C(_15793_),
    .Y(_15794_));
 OA21x2_ASAP7_75t_R _21180_ (.A1(_15784_),
    .A2(_15787_),
    .B(_15794_),
    .Y(_15795_));
 INVx1_ASAP7_75t_R _21181_ (.A(_00840_),
    .Y(_15796_));
 NAND2x1_ASAP7_75t_R _21182_ (.A(net342),
    .B(_00838_),
    .Y(_15797_));
 OA211x2_ASAP7_75t_R _21183_ (.A1(net342),
    .A2(_15796_),
    .B(_15797_),
    .C(net311),
    .Y(_15798_));
 INVx1_ASAP7_75t_R _21184_ (.A(_00839_),
    .Y(_15799_));
 NAND2x1_ASAP7_75t_R _21185_ (.A(net342),
    .B(_00837_),
    .Y(_15800_));
 OA211x2_ASAP7_75t_R _21186_ (.A1(net342),
    .A2(_15799_),
    .B(_15800_),
    .C(net356),
    .Y(_15801_));
 OR3x1_ASAP7_75t_R _21187_ (.A(net323),
    .B(_15798_),
    .C(_15801_),
    .Y(_15802_));
 INVx1_ASAP7_75t_R _21188_ (.A(_00836_),
    .Y(_15803_));
 NAND2x1_ASAP7_75t_R _21189_ (.A(net342),
    .B(_00834_),
    .Y(_15804_));
 OA211x2_ASAP7_75t_R _21190_ (.A1(net342),
    .A2(_15803_),
    .B(_15804_),
    .C(net311),
    .Y(_15805_));
 INVx1_ASAP7_75t_R _21191_ (.A(_00835_),
    .Y(_15806_));
 NAND2x1_ASAP7_75t_R _21192_ (.A(net342),
    .B(_00833_),
    .Y(_15807_));
 OA211x2_ASAP7_75t_R _21193_ (.A1(net342),
    .A2(_15806_),
    .B(_15807_),
    .C(net356),
    .Y(_15808_));
 OR3x1_ASAP7_75t_R _21194_ (.A(_13132_),
    .B(_15805_),
    .C(_15808_),
    .Y(_15809_));
 AND3x1_ASAP7_75t_R _21195_ (.A(net318),
    .B(_15802_),
    .C(_15809_),
    .Y(_15810_));
 AO21x1_ASAP7_75t_R _21196_ (.A1(_13598_),
    .A2(_15795_),
    .B(_15810_),
    .Y(_15811_));
 INVx1_ASAP7_75t_R _21197_ (.A(_00819_),
    .Y(_15812_));
 INVx1_ASAP7_75t_R _21198_ (.A(_00820_),
    .Y(_15813_));
 NAND2x1_ASAP7_75t_R _21199_ (.A(net343),
    .B(_01692_),
    .Y(_15814_));
 OA211x2_ASAP7_75t_R _21200_ (.A1(net343),
    .A2(_15813_),
    .B(_15814_),
    .C(net311),
    .Y(_15815_));
 AO21x1_ASAP7_75t_R _21201_ (.A1(_15812_),
    .A2(_13190_),
    .B(_15815_),
    .Y(_15816_));
 INVx1_ASAP7_75t_R _21202_ (.A(_00828_),
    .Y(_15817_));
 NAND2x1_ASAP7_75t_R _21203_ (.A(net343),
    .B(_00826_),
    .Y(_15818_));
 OA211x2_ASAP7_75t_R _21204_ (.A1(net343),
    .A2(_15817_),
    .B(_15818_),
    .C(net311),
    .Y(_15819_));
 INVx1_ASAP7_75t_R _21205_ (.A(_00827_),
    .Y(_15820_));
 NAND2x1_ASAP7_75t_R _21206_ (.A(net343),
    .B(_00825_),
    .Y(_15821_));
 OA211x2_ASAP7_75t_R _21207_ (.A1(net343),
    .A2(_15820_),
    .B(_15821_),
    .C(net356),
    .Y(_15822_));
 OR3x1_ASAP7_75t_R _21208_ (.A(net317),
    .B(_15819_),
    .C(_15822_),
    .Y(_15823_));
 OA211x2_ASAP7_75t_R _21209_ (.A1(_13598_),
    .A2(_15816_),
    .B(_15823_),
    .C(net323),
    .Y(_15824_));
 INVx1_ASAP7_75t_R _21210_ (.A(_00829_),
    .Y(_15825_));
 NOR2x1_ASAP7_75t_R _21211_ (.A(net343),
    .B(_00831_),
    .Y(_15826_));
 AO21x1_ASAP7_75t_R _21212_ (.A1(net343),
    .A2(_15825_),
    .B(_15826_),
    .Y(_15827_));
 INVx1_ASAP7_75t_R _21213_ (.A(_00832_),
    .Y(_15828_));
 NAND2x1_ASAP7_75t_R _21214_ (.A(net343),
    .B(_00830_),
    .Y(_15829_));
 OA211x2_ASAP7_75t_R _21215_ (.A1(net343),
    .A2(_15828_),
    .B(_15829_),
    .C(net311),
    .Y(_15830_));
 AO21x1_ASAP7_75t_R _21216_ (.A1(net356),
    .A2(_15827_),
    .B(_15830_),
    .Y(_15831_));
 INVx1_ASAP7_75t_R _21217_ (.A(_00824_),
    .Y(_15832_));
 NAND2x1_ASAP7_75t_R _21218_ (.A(net343),
    .B(_00822_),
    .Y(_15833_));
 OA211x2_ASAP7_75t_R _21219_ (.A1(net343),
    .A2(_15832_),
    .B(_15833_),
    .C(net311),
    .Y(_15834_));
 INVx1_ASAP7_75t_R _21220_ (.A(_00823_),
    .Y(_15835_));
 NAND2x1_ASAP7_75t_R _21221_ (.A(net343),
    .B(_00821_),
    .Y(_15836_));
 OA211x2_ASAP7_75t_R _21222_ (.A1(net343),
    .A2(_15835_),
    .B(_15836_),
    .C(net356),
    .Y(_15837_));
 OR3x1_ASAP7_75t_R _21223_ (.A(_13598_),
    .B(_15834_),
    .C(_15837_),
    .Y(_15838_));
 OA211x2_ASAP7_75t_R _21224_ (.A1(net317),
    .A2(_15831_),
    .B(_15838_),
    .C(_13132_),
    .Y(_15839_));
 OA21x2_ASAP7_75t_R _21225_ (.A1(_15824_),
    .A2(_15839_),
    .B(net314),
    .Y(_15840_));
 AO21x2_ASAP7_75t_R _21226_ (.A1(_13174_),
    .A2(_15811_),
    .B(_15840_),
    .Y(_15841_));
 INVx2_ASAP7_75t_R _21227_ (.A(_15841_),
    .Y(_15842_));
 OA21x2_ASAP7_75t_R _21228_ (.A1(net371),
    .A2(_15268_),
    .B(_15269_),
    .Y(_15843_));
 AO21x2_ASAP7_75t_R _21229_ (.A1(_13583_),
    .A2(_15842_),
    .B(_15843_),
    .Y(_18190_));
 INVx1_ASAP7_75t_R _21230_ (.A(_18190_),
    .Y(_18192_));
 XNOR2x1_ASAP7_75t_R _21231_ (.B(_18190_),
    .Y(_15844_),
    .A(_13387_));
 NAND2x1_ASAP7_75t_R _21232_ (.A(net387),
    .B(_00838_),
    .Y(_15845_));
 OA211x2_ASAP7_75t_R _21233_ (.A1(net387),
    .A2(_15796_),
    .B(_15845_),
    .C(net307),
    .Y(_15846_));
 NAND2x1_ASAP7_75t_R _21234_ (.A(net387),
    .B(_00837_),
    .Y(_15847_));
 OA211x2_ASAP7_75t_R _21235_ (.A1(net387),
    .A2(_15799_),
    .B(_15847_),
    .C(net407),
    .Y(_15848_));
 OR3x1_ASAP7_75t_R _21236_ (.A(net369),
    .B(_15846_),
    .C(_15848_),
    .Y(_15849_));
 NAND2x1_ASAP7_75t_R _21237_ (.A(net387),
    .B(_00834_),
    .Y(_15850_));
 OA211x2_ASAP7_75t_R _21238_ (.A1(net387),
    .A2(_15803_),
    .B(_15850_),
    .C(net307),
    .Y(_15851_));
 NAND2x1_ASAP7_75t_R _21239_ (.A(net387),
    .B(_00833_),
    .Y(_15852_));
 OA211x2_ASAP7_75t_R _21240_ (.A1(net387),
    .A2(_15806_),
    .B(_15852_),
    .C(net407),
    .Y(_15853_));
 OR3x1_ASAP7_75t_R _21241_ (.A(_13397_),
    .B(_15851_),
    .C(_15853_),
    .Y(_15854_));
 NAND2x1_ASAP7_75t_R _21242_ (.A(net387),
    .B(_00822_),
    .Y(_15855_));
 OA211x2_ASAP7_75t_R _21243_ (.A1(net387),
    .A2(_15832_),
    .B(_15855_),
    .C(net307),
    .Y(_15856_));
 NAND2x1_ASAP7_75t_R _21244_ (.A(net387),
    .B(_00821_),
    .Y(_15857_));
 OA211x2_ASAP7_75t_R _21245_ (.A1(net387),
    .A2(_15835_),
    .B(_15857_),
    .C(net407),
    .Y(_15858_));
 OR3x1_ASAP7_75t_R _21246_ (.A(net298),
    .B(_15856_),
    .C(_15858_),
    .Y(_15859_));
 NAND2x1_ASAP7_75t_R _21247_ (.A(net395),
    .B(_01692_),
    .Y(_15860_));
 OA211x2_ASAP7_75t_R _21248_ (.A1(net395),
    .A2(_15813_),
    .B(_15860_),
    .C(net307),
    .Y(_15861_));
 AND3x1_ASAP7_75t_R _21249_ (.A(net409),
    .B(net303),
    .C(_15812_),
    .Y(_15862_));
 OA31x2_ASAP7_75t_R _21250_ (.A1(net301),
    .A2(_15861_),
    .A3(_15862_),
    .B1(net363),
    .Y(_15863_));
 AO32x1_ASAP7_75t_R _21251_ (.A1(_13392_),
    .A2(_15849_),
    .A3(_15854_),
    .B1(_15859_),
    .B2(_15863_),
    .Y(_15864_));
 NOR2x1_ASAP7_75t_R _21252_ (.A(net387),
    .B(_00831_),
    .Y(_15865_));
 AO21x1_ASAP7_75t_R _21253_ (.A1(net387),
    .A2(_15825_),
    .B(_15865_),
    .Y(_15866_));
 NAND2x1_ASAP7_75t_R _21254_ (.A(net387),
    .B(_00830_),
    .Y(_15867_));
 OA211x2_ASAP7_75t_R _21255_ (.A1(net387),
    .A2(_15828_),
    .B(_15867_),
    .C(net307),
    .Y(_15868_));
 AO21x1_ASAP7_75t_R _21256_ (.A1(net409),
    .A2(_15866_),
    .B(_15868_),
    .Y(_15869_));
 NAND2x1_ASAP7_75t_R _21257_ (.A(net387),
    .B(_00826_),
    .Y(_15870_));
 OA211x2_ASAP7_75t_R _21258_ (.A1(net387),
    .A2(_15817_),
    .B(_15870_),
    .C(net305),
    .Y(_15871_));
 NAND2x1_ASAP7_75t_R _21259_ (.A(net395),
    .B(_00825_),
    .Y(_15872_));
 OA211x2_ASAP7_75t_R _21260_ (.A1(net387),
    .A2(_15820_),
    .B(_15872_),
    .C(net409),
    .Y(_15873_));
 OA21x2_ASAP7_75t_R _21261_ (.A1(_15871_),
    .A2(_15873_),
    .B(net369),
    .Y(_15874_));
 AO21x1_ASAP7_75t_R _21262_ (.A1(_13397_),
    .A2(_15869_),
    .B(_15874_),
    .Y(_15875_));
 AND2x2_ASAP7_75t_R _21263_ (.A(_15859_),
    .B(_15863_),
    .Y(_15876_));
 NAND2x1_ASAP7_75t_R _21264_ (.A(net369),
    .B(_00844_),
    .Y(_15877_));
 OA211x2_ASAP7_75t_R _21265_ (.A1(net369),
    .A2(_15788_),
    .B(_15877_),
    .C(net307),
    .Y(_15878_));
 NAND2x1_ASAP7_75t_R _21266_ (.A(net369),
    .B(_00843_),
    .Y(_15879_));
 OA211x2_ASAP7_75t_R _21267_ (.A1(net369),
    .A2(_15791_),
    .B(_15879_),
    .C(net407),
    .Y(_15880_));
 OR3x1_ASAP7_75t_R _21268_ (.A(net387),
    .B(_15878_),
    .C(_15880_),
    .Y(_15881_));
 INVx1_ASAP7_75t_R _21269_ (.A(_00846_),
    .Y(_15882_));
 NAND2x1_ASAP7_75t_R _21270_ (.A(net369),
    .B(_00842_),
    .Y(_15883_));
 OA211x2_ASAP7_75t_R _21271_ (.A1(net369),
    .A2(_15882_),
    .B(_15883_),
    .C(net307),
    .Y(_15884_));
 INVx1_ASAP7_75t_R _21272_ (.A(_00845_),
    .Y(_15885_));
 NAND2x1_ASAP7_75t_R _21273_ (.A(net369),
    .B(_00841_),
    .Y(_15886_));
 OA211x2_ASAP7_75t_R _21274_ (.A1(net369),
    .A2(_15885_),
    .B(_15886_),
    .C(net407),
    .Y(_15887_));
 OR3x1_ASAP7_75t_R _21275_ (.A(net303),
    .B(_15884_),
    .C(_15887_),
    .Y(_15888_));
 AND3x1_ASAP7_75t_R _21276_ (.A(_14571_),
    .B(_15881_),
    .C(_15888_),
    .Y(_15889_));
 AO221x2_ASAP7_75t_R _21277_ (.A1(net366),
    .A2(_15864_),
    .B1(_15875_),
    .B2(_15876_),
    .C(_15889_),
    .Y(_15890_));
 NOR2x1_ASAP7_75t_R _21278_ (.A(_00284_),
    .B(_15890_),
    .Y(_15891_));
 BUFx16f_ASAP7_75t_R load_slew267 (.A(_09941_),
    .Y(net267));
 AO221x1_ASAP7_75t_R _21280_ (.A1(_13530_),
    .A2(_00849_),
    .B1(_02216_),
    .B2(_13533_),
    .C(_13528_),
    .Y(_15893_));
 OA22x2_ASAP7_75t_R _21281_ (.A1(_13763_),
    .A2(_15842_),
    .B1(_15891_),
    .B2(_15893_),
    .Y(_15894_));
 NOR2x1_ASAP7_75t_R _21282_ (.A(net295),
    .B(_15894_),
    .Y(_15895_));
 AOI21x1_ASAP7_75t_R _21283_ (.A1(net295),
    .A2(_15844_),
    .B(_15895_),
    .Y(_17566_));
 INVx1_ASAP7_75t_R _21284_ (.A(_17566_),
    .Y(_16525_));
 INVx3_ASAP7_75t_R _21285_ (.A(_00209_),
    .Y(\cs_registers_i.pc_id_i[17] ));
 NOR2x1_ASAP7_75t_R _21286_ (.A(_01624_),
    .B(_13223_),
    .Y(_15896_));
 AOI221x1_ASAP7_75t_R _21287_ (.A1(\cs_registers_i.pc_id_i[17] ),
    .A2(_14503_),
    .B1(_15890_),
    .B2(_13563_),
    .C(_15896_),
    .Y(_15897_));
 BUFx12f_ASAP7_75t_R load_slew266 (.A(_10103_),
    .Y(net266));
 OA21x2_ASAP7_75t_R _21289_ (.A1(_00849_),
    .A2(_13574_),
    .B(_13576_),
    .Y(_15898_));
 AOI21x1_ASAP7_75t_R _21290_ (.A1(net294),
    .A2(_15897_),
    .B(_15898_),
    .Y(_17567_));
 INVx1_ASAP7_75t_R _21291_ (.A(_17567_),
    .Y(_16526_));
 AO21x1_ASAP7_75t_R _21292_ (.A1(_02273_),
    .A2(_15670_),
    .B(_00784_),
    .Y(_15899_));
 AO21x1_ASAP7_75t_R _21293_ (.A1(_00817_),
    .A2(_15899_),
    .B(_02275_),
    .Y(_15900_));
 AND2x2_ASAP7_75t_R _21294_ (.A(_02274_),
    .B(_15900_),
    .Y(_16527_));
 AND2x2_ASAP7_75t_R _21295_ (.A(net338),
    .B(_01691_),
    .Y(_15901_));
 AO21x1_ASAP7_75t_R _21296_ (.A1(net313),
    .A2(_00852_),
    .B(_15901_),
    .Y(_15902_));
 OAI22x1_ASAP7_75t_R _21297_ (.A1(_00851_),
    .A2(_13586_),
    .B1(_15902_),
    .B2(net359),
    .Y(_15903_));
 BUFx16f_ASAP7_75t_R load_slew265 (.A(net266),
    .Y(net265));
 INVx1_ASAP7_75t_R _21299_ (.A(_00860_),
    .Y(_15905_));
 NAND2x1_ASAP7_75t_R _21300_ (.A(net339),
    .B(_00858_),
    .Y(_15906_));
 OA211x2_ASAP7_75t_R _21301_ (.A1(net339),
    .A2(_15905_),
    .B(_15906_),
    .C(net308),
    .Y(_15907_));
 INVx1_ASAP7_75t_R _21302_ (.A(_00859_),
    .Y(_15908_));
 NAND2x1_ASAP7_75t_R _21303_ (.A(net339),
    .B(_00857_),
    .Y(_15909_));
 BUFx16f_ASAP7_75t_R load_slew264 (.A(net265),
    .Y(net264));
 OA211x2_ASAP7_75t_R _21305_ (.A1(net339),
    .A2(_15908_),
    .B(_15909_),
    .C(net359),
    .Y(_15911_));
 OR3x1_ASAP7_75t_R _21306_ (.A(net319),
    .B(_15907_),
    .C(_15911_),
    .Y(_15912_));
 OA211x2_ASAP7_75t_R _21307_ (.A1(_13598_),
    .A2(_15903_),
    .B(_15912_),
    .C(net325),
    .Y(_15913_));
 BUFx16f_ASAP7_75t_R load_slew263 (.A(_10456_),
    .Y(net263));
 INVx1_ASAP7_75t_R _21309_ (.A(_00856_),
    .Y(_15915_));
 NAND2x1_ASAP7_75t_R _21310_ (.A(net339),
    .B(_00854_),
    .Y(_15916_));
 BUFx16f_ASAP7_75t_R load_slew262 (.A(net263),
    .Y(net262));
 OA211x2_ASAP7_75t_R _21312_ (.A1(net339),
    .A2(_15915_),
    .B(_15916_),
    .C(net308),
    .Y(_15918_));
 BUFx16f_ASAP7_75t_R load_slew261 (.A(_10648_),
    .Y(net261));
 INVx1_ASAP7_75t_R _21314_ (.A(_00855_),
    .Y(_15920_));
 NAND2x1_ASAP7_75t_R _21315_ (.A(net339),
    .B(_00853_),
    .Y(_15921_));
 BUFx16f_ASAP7_75t_R load_slew260 (.A(_10648_),
    .Y(net260));
 OA211x2_ASAP7_75t_R _21317_ (.A1(net339),
    .A2(_15920_),
    .B(_15921_),
    .C(net359),
    .Y(_15923_));
 OR3x1_ASAP7_75t_R _21318_ (.A(_13598_),
    .B(_15918_),
    .C(_15923_),
    .Y(_15924_));
 INVx1_ASAP7_75t_R _21319_ (.A(_00864_),
    .Y(_15925_));
 NAND2x1_ASAP7_75t_R _21320_ (.A(net339),
    .B(_00862_),
    .Y(_15926_));
 OA211x2_ASAP7_75t_R _21321_ (.A1(net339),
    .A2(_15925_),
    .B(_15926_),
    .C(net308),
    .Y(_15927_));
 BUFx16f_ASAP7_75t_R load_slew259 (.A(_10808_),
    .Y(net259));
 INVx1_ASAP7_75t_R _21323_ (.A(_00863_),
    .Y(_15929_));
 BUFx16f_ASAP7_75t_R load_slew258 (.A(net259),
    .Y(net258));
 NAND2x1_ASAP7_75t_R _21325_ (.A(net339),
    .B(_00861_),
    .Y(_15931_));
 OA211x2_ASAP7_75t_R _21326_ (.A1(net339),
    .A2(_15929_),
    .B(_15931_),
    .C(net359),
    .Y(_15932_));
 OR3x1_ASAP7_75t_R _21327_ (.A(net319),
    .B(_15927_),
    .C(_15932_),
    .Y(_15933_));
 AND3x1_ASAP7_75t_R _21328_ (.A(_13132_),
    .B(_15924_),
    .C(_15933_),
    .Y(_15934_));
 OR3x2_ASAP7_75t_R _21329_ (.A(_13174_),
    .B(_15913_),
    .C(_15934_),
    .Y(_15935_));
 BUFx6f_ASAP7_75t_R load_slew257 (.A(net160),
    .Y(net257));
 INVx1_ASAP7_75t_R _21331_ (.A(_00872_),
    .Y(_15937_));
 NAND2x1_ASAP7_75t_R _21332_ (.A(net336),
    .B(_00870_),
    .Y(_15938_));
 OA211x2_ASAP7_75t_R _21333_ (.A1(net336),
    .A2(_15937_),
    .B(_15938_),
    .C(_13145_),
    .Y(_15939_));
 INVx1_ASAP7_75t_R _21334_ (.A(_00871_),
    .Y(_15940_));
 NAND2x1_ASAP7_75t_R _21335_ (.A(net336),
    .B(_00869_),
    .Y(_15941_));
 OA211x2_ASAP7_75t_R _21336_ (.A1(net336),
    .A2(_15940_),
    .B(_15941_),
    .C(net358),
    .Y(_15942_));
 OR3x1_ASAP7_75t_R _21337_ (.A(_13598_),
    .B(_15939_),
    .C(_15942_),
    .Y(_15943_));
 INVx1_ASAP7_75t_R _21338_ (.A(_00880_),
    .Y(_15944_));
 NAND2x1_ASAP7_75t_R _21339_ (.A(net336),
    .B(_00878_),
    .Y(_15945_));
 OA211x2_ASAP7_75t_R _21340_ (.A1(net336),
    .A2(_15944_),
    .B(_15945_),
    .C(_13145_),
    .Y(_15946_));
 INVx1_ASAP7_75t_R _21341_ (.A(_00879_),
    .Y(_15947_));
 NAND2x1_ASAP7_75t_R _21342_ (.A(net336),
    .B(_00877_),
    .Y(_15948_));
 OA211x2_ASAP7_75t_R _21343_ (.A1(net336),
    .A2(_15947_),
    .B(_15948_),
    .C(net358),
    .Y(_15949_));
 OR3x1_ASAP7_75t_R _21344_ (.A(net318),
    .B(_15946_),
    .C(_15949_),
    .Y(_15950_));
 AND3x1_ASAP7_75t_R _21345_ (.A(_13132_),
    .B(_15943_),
    .C(_15950_),
    .Y(_15951_));
 INVx1_ASAP7_75t_R _21346_ (.A(_00873_),
    .Y(_15952_));
 BUFx4f_ASAP7_75t_R load_slew256 (.A(_00785_),
    .Y(net256));
 NOR2x1_ASAP7_75t_R _21348_ (.A(net336),
    .B(_00875_),
    .Y(_15954_));
 AO21x1_ASAP7_75t_R _21349_ (.A1(net336),
    .A2(_15952_),
    .B(_15954_),
    .Y(_15955_));
 BUFx6f_ASAP7_75t_R load_slew255 (.A(net162),
    .Y(net255));
 BUFx12f_ASAP7_75t_R max_cap254 (.A(_11601_),
    .Y(net254));
 INVx1_ASAP7_75t_R _21352_ (.A(_00876_),
    .Y(_15958_));
 NAND2x1_ASAP7_75t_R _21353_ (.A(net336),
    .B(_00874_),
    .Y(_15959_));
 OA211x2_ASAP7_75t_R _21354_ (.A1(net336),
    .A2(_15958_),
    .B(_15959_),
    .C(_13145_),
    .Y(_15960_));
 AO21x1_ASAP7_75t_R _21355_ (.A1(net358),
    .A2(_15955_),
    .B(_15960_),
    .Y(_15961_));
 INVx1_ASAP7_75t_R _21356_ (.A(_00868_),
    .Y(_15962_));
 NAND2x1_ASAP7_75t_R _21357_ (.A(net336),
    .B(_00866_),
    .Y(_15963_));
 OA211x2_ASAP7_75t_R _21358_ (.A1(net336),
    .A2(_15962_),
    .B(_15963_),
    .C(_13145_),
    .Y(_15964_));
 INVx1_ASAP7_75t_R _21359_ (.A(_00867_),
    .Y(_15965_));
 NAND2x1_ASAP7_75t_R _21360_ (.A(net336),
    .B(_00865_),
    .Y(_15966_));
 OA211x2_ASAP7_75t_R _21361_ (.A1(net336),
    .A2(_15965_),
    .B(_15966_),
    .C(net358),
    .Y(_15967_));
 OR3x1_ASAP7_75t_R _21362_ (.A(_13598_),
    .B(_15964_),
    .C(_15967_),
    .Y(_15968_));
 OA211x2_ASAP7_75t_R _21363_ (.A1(net319),
    .A2(_15961_),
    .B(_15968_),
    .C(net325),
    .Y(_15969_));
 OR3x4_ASAP7_75t_R _21364_ (.A(net315),
    .B(_15951_),
    .C(_15969_),
    .Y(_15970_));
 NAND2x2_ASAP7_75t_R _21365_ (.A(_15935_),
    .B(_15970_),
    .Y(_15971_));
 OA21x2_ASAP7_75t_R _21366_ (.A1(net367),
    .A2(_15268_),
    .B(_15269_),
    .Y(_15972_));
 AOI21x1_ASAP7_75t_R _21367_ (.A1(_13583_),
    .A2(_15971_),
    .B(_15972_),
    .Y(_18197_));
 AND2x2_ASAP7_75t_R _21368_ (.A(net399),
    .B(_01691_),
    .Y(_15973_));
 AO21x1_ASAP7_75t_R _21369_ (.A1(net302),
    .A2(_00852_),
    .B(_15973_),
    .Y(_15974_));
 OAI22x1_ASAP7_75t_R _21370_ (.A1(_00851_),
    .A2(_13471_),
    .B1(_15974_),
    .B2(net410),
    .Y(_15975_));
 NAND2x1_ASAP7_75t_R _21371_ (.A(net398),
    .B(_00858_),
    .Y(_15976_));
 OA211x2_ASAP7_75t_R _21372_ (.A1(net398),
    .A2(_15905_),
    .B(_15976_),
    .C(net306),
    .Y(_15977_));
 NAND2x1_ASAP7_75t_R _21373_ (.A(net398),
    .B(_00857_),
    .Y(_15978_));
 OA211x2_ASAP7_75t_R _21374_ (.A1(net398),
    .A2(_15908_),
    .B(_15978_),
    .C(_00290_),
    .Y(_15979_));
 OR3x1_ASAP7_75t_R _21375_ (.A(net367),
    .B(_15977_),
    .C(_15979_),
    .Y(_15980_));
 OA211x2_ASAP7_75t_R _21376_ (.A1(_13484_),
    .A2(_15975_),
    .B(_15980_),
    .C(net371),
    .Y(_15981_));
 NAND2x1_ASAP7_75t_R _21377_ (.A(net398),
    .B(_00853_),
    .Y(_15982_));
 OA211x2_ASAP7_75t_R _21378_ (.A1(net398),
    .A2(_15920_),
    .B(_15982_),
    .C(net367),
    .Y(_15983_));
 NAND2x1_ASAP7_75t_R _21379_ (.A(net398),
    .B(_00861_),
    .Y(_15984_));
 OA211x2_ASAP7_75t_R _21380_ (.A1(net398),
    .A2(_15929_),
    .B(_15984_),
    .C(_13484_),
    .Y(_15985_));
 OR3x1_ASAP7_75t_R _21381_ (.A(net306),
    .B(_15983_),
    .C(_15985_),
    .Y(_15986_));
 NAND2x1_ASAP7_75t_R _21382_ (.A(net367),
    .B(_00856_),
    .Y(_15987_));
 OA211x2_ASAP7_75t_R _21383_ (.A1(net367),
    .A2(_15925_),
    .B(_15987_),
    .C(net302),
    .Y(_15988_));
 INVx1_ASAP7_75t_R _21384_ (.A(_00862_),
    .Y(_15989_));
 NAND2x1_ASAP7_75t_R _21385_ (.A(net367),
    .B(_00854_),
    .Y(_15990_));
 OA211x2_ASAP7_75t_R _21386_ (.A1(net367),
    .A2(_15989_),
    .B(_15990_),
    .C(net398),
    .Y(_15991_));
 OR3x1_ASAP7_75t_R _21387_ (.A(_00290_),
    .B(_15988_),
    .C(_15991_),
    .Y(_15992_));
 AND3x1_ASAP7_75t_R _21388_ (.A(_13397_),
    .B(_15986_),
    .C(_15992_),
    .Y(_15993_));
 OR3x2_ASAP7_75t_R _21389_ (.A(_13392_),
    .B(_15981_),
    .C(_15993_),
    .Y(_15994_));
 NOR2x1_ASAP7_75t_R _21390_ (.A(net397),
    .B(_00875_),
    .Y(_15995_));
 AO21x1_ASAP7_75t_R _21391_ (.A1(net397),
    .A2(_15952_),
    .B(_15995_),
    .Y(_15996_));
 NAND2x1_ASAP7_75t_R _21392_ (.A(net397),
    .B(_00874_),
    .Y(_15997_));
 OA211x2_ASAP7_75t_R _21393_ (.A1(net397),
    .A2(_15958_),
    .B(_15997_),
    .C(net306),
    .Y(_15998_));
 AO21x1_ASAP7_75t_R _21394_ (.A1(net410),
    .A2(_15996_),
    .B(_15998_),
    .Y(_15999_));
 NAND2x1_ASAP7_75t_R _21395_ (.A(net397),
    .B(_00878_),
    .Y(_16000_));
 OA211x2_ASAP7_75t_R _21396_ (.A1(net397),
    .A2(_15944_),
    .B(_16000_),
    .C(_13424_),
    .Y(_16001_));
 NAND2x1_ASAP7_75t_R _21397_ (.A(net397),
    .B(_00877_),
    .Y(_16002_));
 OA211x2_ASAP7_75t_R _21398_ (.A1(net397),
    .A2(_15947_),
    .B(_16002_),
    .C(net410),
    .Y(_16003_));
 OR3x1_ASAP7_75t_R _21399_ (.A(net371),
    .B(_16001_),
    .C(_16003_),
    .Y(_16004_));
 OA211x2_ASAP7_75t_R _21400_ (.A1(_13397_),
    .A2(_15999_),
    .B(_16004_),
    .C(_13484_),
    .Y(_16005_));
 NAND2x1_ASAP7_75t_R _21401_ (.A(net397),
    .B(_00866_),
    .Y(_16006_));
 OA211x2_ASAP7_75t_R _21402_ (.A1(net397),
    .A2(_15962_),
    .B(_16006_),
    .C(net306),
    .Y(_16007_));
 NAND2x1_ASAP7_75t_R _21403_ (.A(net397),
    .B(_00865_),
    .Y(_16008_));
 OA211x2_ASAP7_75t_R _21404_ (.A1(net397),
    .A2(_15965_),
    .B(_16008_),
    .C(net410),
    .Y(_16009_));
 OR3x1_ASAP7_75t_R _21405_ (.A(_13397_),
    .B(_16007_),
    .C(_16009_),
    .Y(_16010_));
 NAND2x1_ASAP7_75t_R _21406_ (.A(net397),
    .B(_00870_),
    .Y(_16011_));
 OA211x2_ASAP7_75t_R _21407_ (.A1(net397),
    .A2(_15937_),
    .B(_16011_),
    .C(_13424_),
    .Y(_16012_));
 NAND2x1_ASAP7_75t_R _21408_ (.A(net397),
    .B(_00869_),
    .Y(_16013_));
 OA211x2_ASAP7_75t_R _21409_ (.A1(net397),
    .A2(_15940_),
    .B(_16013_),
    .C(net410),
    .Y(_16014_));
 OR3x1_ASAP7_75t_R _21410_ (.A(net371),
    .B(_16012_),
    .C(_16014_),
    .Y(_16015_));
 AND3x1_ASAP7_75t_R _21411_ (.A(net365),
    .B(_16010_),
    .C(_16015_),
    .Y(_16016_));
 OR3x4_ASAP7_75t_R _21412_ (.A(net364),
    .B(_16005_),
    .C(_16016_),
    .Y(_16017_));
 NAND2x2_ASAP7_75t_R _21413_ (.A(_15994_),
    .B(_16017_),
    .Y(_16018_));
 OA22x2_ASAP7_75t_R _21414_ (.A1(_01623_),
    .A2(_13223_),
    .B1(_13880_),
    .B2(_00211_),
    .Y(_16019_));
 OAI21x1_ASAP7_75t_R _21415_ (.A1(_13782_),
    .A2(_16018_),
    .B(_16019_),
    .Y(_18198_));
 INVx3_ASAP7_75t_R _21416_ (.A(_18198_),
    .Y(_18196_));
 XOR2x2_ASAP7_75t_R _21417_ (.A(_00882_),
    .B(_02228_),
    .Y(_16020_));
 INVx4_ASAP7_75t_R _21418_ (.A(_16020_),
    .Y(net159));
 INVx1_ASAP7_75t_R _21419_ (.A(_00893_),
    .Y(_16021_));
 NAND2x1_ASAP7_75t_R _21420_ (.A(net338),
    .B(_00891_),
    .Y(_16022_));
 OA211x2_ASAP7_75t_R _21421_ (.A1(net338),
    .A2(_16021_),
    .B(_16022_),
    .C(net308),
    .Y(_16023_));
 INVx1_ASAP7_75t_R _21422_ (.A(_00892_),
    .Y(_16024_));
 NAND2x1_ASAP7_75t_R _21423_ (.A(net338),
    .B(_00890_),
    .Y(_16025_));
 OA211x2_ASAP7_75t_R _21424_ (.A1(net338),
    .A2(_16024_),
    .B(_16025_),
    .C(net358),
    .Y(_16026_));
 OR3x1_ASAP7_75t_R _21425_ (.A(net319),
    .B(_16023_),
    .C(_16026_),
    .Y(_16027_));
 INVx1_ASAP7_75t_R _21426_ (.A(_00884_),
    .Y(_16028_));
 INVx1_ASAP7_75t_R _21427_ (.A(_00885_),
    .Y(_16029_));
 NAND2x1_ASAP7_75t_R _21428_ (.A(net334),
    .B(_01690_),
    .Y(_16030_));
 OA21x2_ASAP7_75t_R _21429_ (.A1(net334),
    .A2(_16029_),
    .B(_16030_),
    .Y(_16031_));
 BUFx16f_ASAP7_75t_R max_cap253 (.A(_07620_),
    .Y(net253));
 AO221x1_ASAP7_75t_R _21431_ (.A1(_16028_),
    .A2(_13190_),
    .B1(_16031_),
    .B2(net308),
    .C(_13598_),
    .Y(_16033_));
 AO21x1_ASAP7_75t_R _21432_ (.A1(_16027_),
    .A2(_16033_),
    .B(_13132_),
    .Y(_16034_));
 INVx1_ASAP7_75t_R _21433_ (.A(_00889_),
    .Y(_16035_));
 NAND2x1_ASAP7_75t_R _21434_ (.A(net333),
    .B(_00887_),
    .Y(_16036_));
 OA211x2_ASAP7_75t_R _21435_ (.A1(net333),
    .A2(_16035_),
    .B(_16036_),
    .C(net308),
    .Y(_16037_));
 INVx1_ASAP7_75t_R _21436_ (.A(_00888_),
    .Y(_16038_));
 NAND2x1_ASAP7_75t_R _21437_ (.A(net333),
    .B(_00886_),
    .Y(_16039_));
 OA211x2_ASAP7_75t_R _21438_ (.A1(net333),
    .A2(_16038_),
    .B(_16039_),
    .C(net358),
    .Y(_16040_));
 OR3x1_ASAP7_75t_R _21439_ (.A(_13598_),
    .B(_16037_),
    .C(_16040_),
    .Y(_16041_));
 INVx1_ASAP7_75t_R _21440_ (.A(_00897_),
    .Y(_16042_));
 NAND2x1_ASAP7_75t_R _21441_ (.A(net337),
    .B(_00895_),
    .Y(_16043_));
 OA211x2_ASAP7_75t_R _21442_ (.A1(net337),
    .A2(_16042_),
    .B(_16043_),
    .C(_13145_),
    .Y(_16044_));
 INVx1_ASAP7_75t_R _21443_ (.A(_00896_),
    .Y(_16045_));
 NAND2x1_ASAP7_75t_R _21444_ (.A(net337),
    .B(_00894_),
    .Y(_16046_));
 OA211x2_ASAP7_75t_R _21445_ (.A1(net337),
    .A2(_16045_),
    .B(_16046_),
    .C(net358),
    .Y(_16047_));
 OR3x1_ASAP7_75t_R _21446_ (.A(net319),
    .B(_16044_),
    .C(_16047_),
    .Y(_16048_));
 AO21x1_ASAP7_75t_R _21447_ (.A1(_16041_),
    .A2(_16048_),
    .B(net325),
    .Y(_16049_));
 AO21x2_ASAP7_75t_R _21448_ (.A1(_16034_),
    .A2(_16049_),
    .B(_13174_),
    .Y(_16050_));
 INVx1_ASAP7_75t_R _21449_ (.A(_00901_),
    .Y(_16051_));
 NAND2x1_ASAP7_75t_R _21450_ (.A(net334),
    .B(_00899_),
    .Y(_16052_));
 OA211x2_ASAP7_75t_R _21451_ (.A1(net334),
    .A2(_16051_),
    .B(_16052_),
    .C(_13145_),
    .Y(_16053_));
 INVx1_ASAP7_75t_R _21452_ (.A(_00900_),
    .Y(_16054_));
 NAND2x1_ASAP7_75t_R _21453_ (.A(net334),
    .B(_00898_),
    .Y(_16055_));
 OA211x2_ASAP7_75t_R _21454_ (.A1(net334),
    .A2(_16054_),
    .B(_16055_),
    .C(net358),
    .Y(_16056_));
 OR3x1_ASAP7_75t_R _21455_ (.A(_13132_),
    .B(_16053_),
    .C(_16056_),
    .Y(_16057_));
 INVx1_ASAP7_75t_R _21456_ (.A(_00905_),
    .Y(_16058_));
 NAND2x1_ASAP7_75t_R _21457_ (.A(net334),
    .B(_00903_),
    .Y(_16059_));
 OA211x2_ASAP7_75t_R _21458_ (.A1(net334),
    .A2(_16058_),
    .B(_16059_),
    .C(_13145_),
    .Y(_16060_));
 INVx1_ASAP7_75t_R _21459_ (.A(_00904_),
    .Y(_16061_));
 NAND2x1_ASAP7_75t_R _21460_ (.A(net334),
    .B(_00902_),
    .Y(_16062_));
 OA211x2_ASAP7_75t_R _21461_ (.A1(net334),
    .A2(_16061_),
    .B(_16062_),
    .C(net358),
    .Y(_16063_));
 OR3x1_ASAP7_75t_R _21462_ (.A(net325),
    .B(_16060_),
    .C(_16063_),
    .Y(_16064_));
 AND3x1_ASAP7_75t_R _21463_ (.A(net318),
    .B(_16057_),
    .C(_16064_),
    .Y(_16065_));
 INVx1_ASAP7_75t_R _21464_ (.A(_00906_),
    .Y(_16066_));
 NOR2x1_ASAP7_75t_R _21465_ (.A(net336),
    .B(_00908_),
    .Y(_16067_));
 AO21x1_ASAP7_75t_R _21466_ (.A1(net336),
    .A2(_16066_),
    .B(_16067_),
    .Y(_16068_));
 INVx1_ASAP7_75t_R _21467_ (.A(_00909_),
    .Y(_16069_));
 NAND2x1_ASAP7_75t_R _21468_ (.A(net336),
    .B(_00907_),
    .Y(_16070_));
 OA211x2_ASAP7_75t_R _21469_ (.A1(net336),
    .A2(_16069_),
    .B(_16070_),
    .C(_13145_),
    .Y(_16071_));
 AO21x1_ASAP7_75t_R _21470_ (.A1(net358),
    .A2(_16068_),
    .B(_16071_),
    .Y(_16072_));
 INVx1_ASAP7_75t_R _21471_ (.A(_00913_),
    .Y(_16073_));
 BUFx10_ASAP7_75t_R max_cap252 (.A(_07738_),
    .Y(net252));
 NAND2x1_ASAP7_75t_R _21473_ (.A(net336),
    .B(_00911_),
    .Y(_16075_));
 OA211x2_ASAP7_75t_R _21474_ (.A1(net336),
    .A2(_16073_),
    .B(_16075_),
    .C(_13145_),
    .Y(_16076_));
 INVx1_ASAP7_75t_R _21475_ (.A(_00912_),
    .Y(_16077_));
 NAND2x1_ASAP7_75t_R _21476_ (.A(net336),
    .B(_00910_),
    .Y(_16078_));
 OA211x2_ASAP7_75t_R _21477_ (.A1(net336),
    .A2(_16077_),
    .B(_16078_),
    .C(net358),
    .Y(_16079_));
 OR3x1_ASAP7_75t_R _21478_ (.A(net325),
    .B(_16076_),
    .C(_16079_),
    .Y(_16080_));
 OA211x2_ASAP7_75t_R _21479_ (.A1(_13132_),
    .A2(_16072_),
    .B(_16080_),
    .C(_13598_),
    .Y(_16081_));
 OR3x4_ASAP7_75t_R _21480_ (.A(net315),
    .B(_16065_),
    .C(_16081_),
    .Y(_16082_));
 NAND2x2_ASAP7_75t_R _21481_ (.A(_16050_),
    .B(_16082_),
    .Y(_16083_));
 OA21x2_ASAP7_75t_R _21482_ (.A1(net364),
    .A2(_15268_),
    .B(_15269_),
    .Y(_16084_));
 AO21x2_ASAP7_75t_R _21483_ (.A1(_13583_),
    .A2(_16083_),
    .B(_16084_),
    .Y(_18203_));
 INVx1_ASAP7_75t_R _21484_ (.A(_18203_),
    .Y(_18201_));
 XNOR2x1_ASAP7_75t_R _21485_ (.B(_18203_),
    .Y(_16085_),
    .A(_13387_));
 AND3x1_ASAP7_75t_R _21486_ (.A(_13528_),
    .B(_16050_),
    .C(_16082_),
    .Y(_16086_));
 INVx1_ASAP7_75t_R _21487_ (.A(_00914_),
    .Y(_16087_));
 INVx1_ASAP7_75t_R _21488_ (.A(_02214_),
    .Y(_16088_));
 NAND2x1_ASAP7_75t_R _21489_ (.A(net394),
    .B(_00898_),
    .Y(_16089_));
 OA211x2_ASAP7_75t_R _21490_ (.A1(net394),
    .A2(_16054_),
    .B(_16089_),
    .C(net372),
    .Y(_16090_));
 NAND2x1_ASAP7_75t_R _21491_ (.A(net394),
    .B(_00902_),
    .Y(_16091_));
 OA211x2_ASAP7_75t_R _21492_ (.A1(net394),
    .A2(_16061_),
    .B(_16091_),
    .C(_13397_),
    .Y(_16092_));
 OR3x1_ASAP7_75t_R _21493_ (.A(_13424_),
    .B(_16090_),
    .C(_16092_),
    .Y(_16093_));
 NAND2x1_ASAP7_75t_R _21494_ (.A(net394),
    .B(_00899_),
    .Y(_16094_));
 OA211x2_ASAP7_75t_R _21495_ (.A1(net394),
    .A2(_16051_),
    .B(_16094_),
    .C(net372),
    .Y(_16095_));
 NAND2x1_ASAP7_75t_R _21496_ (.A(net394),
    .B(_00903_),
    .Y(_16096_));
 OA211x2_ASAP7_75t_R _21497_ (.A1(net394),
    .A2(_16058_),
    .B(_16096_),
    .C(_13397_),
    .Y(_16097_));
 OR3x1_ASAP7_75t_R _21498_ (.A(net408),
    .B(_16095_),
    .C(_16097_),
    .Y(_16098_));
 NAND2x1_ASAP7_75t_R _21499_ (.A(net393),
    .B(_00887_),
    .Y(_16099_));
 OA211x2_ASAP7_75t_R _21500_ (.A1(net393),
    .A2(_16035_),
    .B(_16099_),
    .C(net306),
    .Y(_16100_));
 NAND2x1_ASAP7_75t_R _21501_ (.A(net393),
    .B(_00886_),
    .Y(_16101_));
 OA211x2_ASAP7_75t_R _21502_ (.A1(net393),
    .A2(_16038_),
    .B(_16101_),
    .C(net408),
    .Y(_16102_));
 OR3x1_ASAP7_75t_R _21503_ (.A(_13814_),
    .B(_16100_),
    .C(_16102_),
    .Y(_16103_));
 NAND2x1_ASAP7_75t_R _21504_ (.A(net394),
    .B(_01690_),
    .Y(_16104_));
 OA211x2_ASAP7_75t_R _21505_ (.A1(net394),
    .A2(_16029_),
    .B(_16104_),
    .C(net306),
    .Y(_16105_));
 AND3x1_ASAP7_75t_R _21506_ (.A(net408),
    .B(net302),
    .C(_16028_),
    .Y(_16106_));
 OA31x2_ASAP7_75t_R _21507_ (.A1(_13828_),
    .A2(_16105_),
    .A3(_16106_),
    .B1(net364),
    .Y(_16107_));
 AO32x1_ASAP7_75t_R _21508_ (.A1(_13392_),
    .A2(_16093_),
    .A3(_16098_),
    .B1(_16103_),
    .B2(_16107_),
    .Y(_16108_));
 NAND2x1_ASAP7_75t_R _21509_ (.A(net396),
    .B(_00895_),
    .Y(_16109_));
 OA211x2_ASAP7_75t_R _21510_ (.A1(net396),
    .A2(_16042_),
    .B(_16109_),
    .C(net306),
    .Y(_16110_));
 NAND2x1_ASAP7_75t_R _21511_ (.A(net397),
    .B(_00894_),
    .Y(_16111_));
 OA211x2_ASAP7_75t_R _21512_ (.A1(net396),
    .A2(_16045_),
    .B(_16111_),
    .C(net410),
    .Y(_16112_));
 OR3x1_ASAP7_75t_R _21513_ (.A(net371),
    .B(_16110_),
    .C(_16112_),
    .Y(_16113_));
 NAND2x1_ASAP7_75t_R _21514_ (.A(net399),
    .B(_00891_),
    .Y(_16114_));
 OA211x2_ASAP7_75t_R _21515_ (.A1(net399),
    .A2(_16021_),
    .B(_16114_),
    .C(net306),
    .Y(_16115_));
 NAND2x1_ASAP7_75t_R _21516_ (.A(net399),
    .B(_00890_),
    .Y(_16116_));
 OA211x2_ASAP7_75t_R _21517_ (.A1(net399),
    .A2(_16024_),
    .B(_16116_),
    .C(net408),
    .Y(_16117_));
 OR3x1_ASAP7_75t_R _21518_ (.A(_13397_),
    .B(_16115_),
    .C(_16117_),
    .Y(_16118_));
 AND2x2_ASAP7_75t_R _21519_ (.A(_16113_),
    .B(_16118_),
    .Y(_16119_));
 AND2x2_ASAP7_75t_R _21520_ (.A(_16103_),
    .B(_16107_),
    .Y(_16120_));
 NOR2x1_ASAP7_75t_R _21521_ (.A(net371),
    .B(_00910_),
    .Y(_16121_));
 AO21x1_ASAP7_75t_R _21522_ (.A1(net371),
    .A2(_16066_),
    .B(_16121_),
    .Y(_16122_));
 NAND2x1_ASAP7_75t_R _21523_ (.A(net371),
    .B(_00908_),
    .Y(_16123_));
 OA211x2_ASAP7_75t_R _21524_ (.A1(net371),
    .A2(_16077_),
    .B(_16123_),
    .C(net302),
    .Y(_16124_));
 AO21x1_ASAP7_75t_R _21525_ (.A1(net397),
    .A2(_16122_),
    .B(_16124_),
    .Y(_16125_));
 NAND2x1_ASAP7_75t_R _21526_ (.A(net397),
    .B(_00907_),
    .Y(_16126_));
 OA211x2_ASAP7_75t_R _21527_ (.A1(net397),
    .A2(_16069_),
    .B(_16126_),
    .C(net371),
    .Y(_16127_));
 NAND2x1_ASAP7_75t_R _21528_ (.A(net397),
    .B(_00911_),
    .Y(_16128_));
 OA211x2_ASAP7_75t_R _21529_ (.A1(net397),
    .A2(_16073_),
    .B(_16128_),
    .C(_13397_),
    .Y(_16129_));
 OR3x1_ASAP7_75t_R _21530_ (.A(net410),
    .B(_16127_),
    .C(_16129_),
    .Y(_16130_));
 OA211x2_ASAP7_75t_R _21531_ (.A1(net306),
    .A2(_16125_),
    .B(_16130_),
    .C(_14571_),
    .Y(_16131_));
 AO221x2_ASAP7_75t_R _21532_ (.A1(net365),
    .A2(_16108_),
    .B1(_16119_),
    .B2(_16120_),
    .C(_16131_),
    .Y(_16132_));
 OA222x2_ASAP7_75t_R _21533_ (.A1(_00285_),
    .A2(_16087_),
    .B1(_16088_),
    .B2(_13574_),
    .C1(_16132_),
    .C2(_00284_),
    .Y(_16133_));
 AND2x2_ASAP7_75t_R _21534_ (.A(_13763_),
    .B(_16133_),
    .Y(_16134_));
 OA21x2_ASAP7_75t_R _21535_ (.A1(_16086_),
    .A2(_16134_),
    .B(_13576_),
    .Y(_16135_));
 AOI21x1_ASAP7_75t_R _21536_ (.A1(net295),
    .A2(_16085_),
    .B(_16135_),
    .Y(_17570_));
 INVx1_ASAP7_75t_R _21537_ (.A(_17570_),
    .Y(_16528_));
 INVx4_ASAP7_75t_R _21538_ (.A(_00212_),
    .Y(\cs_registers_i.pc_id_i[19] ));
 NOR2x1_ASAP7_75t_R _21539_ (.A(_01622_),
    .B(_13223_),
    .Y(_16136_));
 AOI221x1_ASAP7_75t_R _21540_ (.A1(\cs_registers_i.pc_id_i[19] ),
    .A2(_14503_),
    .B1(_16132_),
    .B2(_13563_),
    .C(_16136_),
    .Y(_16137_));
 BUFx10_ASAP7_75t_R max_cap251 (.A(_08150_),
    .Y(net251));
 OA21x2_ASAP7_75t_R _21542_ (.A1(_00914_),
    .A2(_13574_),
    .B(_13576_),
    .Y(_16138_));
 AOI21x1_ASAP7_75t_R _21543_ (.A1(net295),
    .A2(_16137_),
    .B(_16138_),
    .Y(_17571_));
 INVx1_ASAP7_75t_R _21544_ (.A(_17571_),
    .Y(_16530_));
 OR4x1_ASAP7_75t_R _21545_ (.A(_00784_),
    .B(_00882_),
    .C(_00850_),
    .D(_02275_),
    .Y(_16139_));
 OR3x1_ASAP7_75t_R _21546_ (.A(_00751_),
    .B(_00719_),
    .C(_16139_),
    .Y(_16140_));
 OA21x2_ASAP7_75t_R _21547_ (.A1(_00817_),
    .A2(_02275_),
    .B(_02274_),
    .Y(_16141_));
 OA21x2_ASAP7_75t_R _21548_ (.A1(_00850_),
    .A2(_16141_),
    .B(_00883_),
    .Y(_16142_));
 OA21x2_ASAP7_75t_R _21549_ (.A1(_00751_),
    .A2(_00752_),
    .B(_02273_),
    .Y(_16143_));
 OA21x2_ASAP7_75t_R _21550_ (.A1(_16139_),
    .A2(_16143_),
    .B(_02276_),
    .Y(_16144_));
 OA21x2_ASAP7_75t_R _21551_ (.A1(_00882_),
    .A2(_16142_),
    .B(_16144_),
    .Y(_16145_));
 OA21x2_ASAP7_75t_R _21552_ (.A1(_16521_),
    .A2(_16140_),
    .B(_16145_),
    .Y(_16529_));
 AND2x2_ASAP7_75t_R _21553_ (.A(net346),
    .B(_01689_),
    .Y(_16146_));
 AO21x1_ASAP7_75t_R _21554_ (.A1(net312),
    .A2(_00917_),
    .B(_16146_),
    .Y(_16147_));
 OAI22x1_ASAP7_75t_R _21555_ (.A1(_00916_),
    .A2(_13586_),
    .B1(_16147_),
    .B2(net357),
    .Y(_16148_));
 INVx1_ASAP7_75t_R _21556_ (.A(_00925_),
    .Y(_16149_));
 NAND2x1_ASAP7_75t_R _21557_ (.A(net346),
    .B(_00923_),
    .Y(_16150_));
 OA211x2_ASAP7_75t_R _21558_ (.A1(net346),
    .A2(_16149_),
    .B(_16150_),
    .C(net310),
    .Y(_16151_));
 INVx1_ASAP7_75t_R _21559_ (.A(_00924_),
    .Y(_16152_));
 NAND2x1_ASAP7_75t_R _21560_ (.A(net346),
    .B(_00922_),
    .Y(_16153_));
 OA211x2_ASAP7_75t_R _21561_ (.A1(net346),
    .A2(_16152_),
    .B(_16153_),
    .C(net357),
    .Y(_16154_));
 OR3x1_ASAP7_75t_R _21562_ (.A(net317),
    .B(_16151_),
    .C(_16154_),
    .Y(_16155_));
 OA21x2_ASAP7_75t_R _21563_ (.A1(_13598_),
    .A2(_16148_),
    .B(_16155_),
    .Y(_16156_));
 INVx1_ASAP7_75t_R _21564_ (.A(_00921_),
    .Y(_16157_));
 NAND2x1_ASAP7_75t_R _21565_ (.A(net347),
    .B(_00919_),
    .Y(_16158_));
 OA211x2_ASAP7_75t_R _21566_ (.A1(net347),
    .A2(_16157_),
    .B(_16158_),
    .C(net311),
    .Y(_16159_));
 INVx1_ASAP7_75t_R _21567_ (.A(_00920_),
    .Y(_16160_));
 NAND2x1_ASAP7_75t_R _21568_ (.A(net347),
    .B(_00918_),
    .Y(_16161_));
 OA211x2_ASAP7_75t_R _21569_ (.A1(net347),
    .A2(_16160_),
    .B(_16161_),
    .C(net357),
    .Y(_16162_));
 OR3x1_ASAP7_75t_R _21570_ (.A(_13598_),
    .B(_16159_),
    .C(_16162_),
    .Y(_16163_));
 INVx1_ASAP7_75t_R _21571_ (.A(_00929_),
    .Y(_16164_));
 NAND2x1_ASAP7_75t_R _21572_ (.A(net347),
    .B(_00927_),
    .Y(_16165_));
 OA211x2_ASAP7_75t_R _21573_ (.A1(net347),
    .A2(_16164_),
    .B(_16165_),
    .C(net311),
    .Y(_16166_));
 INVx1_ASAP7_75t_R _21574_ (.A(_00928_),
    .Y(_16167_));
 NAND2x1_ASAP7_75t_R _21575_ (.A(net347),
    .B(_00926_),
    .Y(_16168_));
 OA211x2_ASAP7_75t_R _21576_ (.A1(net347),
    .A2(_16167_),
    .B(_16168_),
    .C(net357),
    .Y(_16169_));
 OR3x1_ASAP7_75t_R _21577_ (.A(net317),
    .B(_16166_),
    .C(_16169_),
    .Y(_16170_));
 AND3x1_ASAP7_75t_R _21578_ (.A(_13132_),
    .B(_16163_),
    .C(_16170_),
    .Y(_16171_));
 AO21x1_ASAP7_75t_R _21579_ (.A1(net324),
    .A2(_16156_),
    .B(_16171_),
    .Y(_16172_));
 INVx1_ASAP7_75t_R _21580_ (.A(_00945_),
    .Y(_16173_));
 NAND2x1_ASAP7_75t_R _21581_ (.A(net343),
    .B(_00943_),
    .Y(_16174_));
 OA211x2_ASAP7_75t_R _21582_ (.A1(net343),
    .A2(_16173_),
    .B(_16174_),
    .C(net311),
    .Y(_16175_));
 INVx1_ASAP7_75t_R _21583_ (.A(_00944_),
    .Y(_16176_));
 NAND2x1_ASAP7_75t_R _21584_ (.A(net343),
    .B(_00942_),
    .Y(_16177_));
 OA211x2_ASAP7_75t_R _21585_ (.A1(net343),
    .A2(_16176_),
    .B(_16177_),
    .C(net357),
    .Y(_16178_));
 OR3x1_ASAP7_75t_R _21586_ (.A(net323),
    .B(_16175_),
    .C(_16178_),
    .Y(_16179_));
 INVx1_ASAP7_75t_R _21587_ (.A(_00941_),
    .Y(_16180_));
 NAND2x1_ASAP7_75t_R _21588_ (.A(net343),
    .B(_00939_),
    .Y(_16181_));
 OA211x2_ASAP7_75t_R _21589_ (.A1(net343),
    .A2(_16180_),
    .B(_16181_),
    .C(net311),
    .Y(_16182_));
 INVx1_ASAP7_75t_R _21590_ (.A(_00940_),
    .Y(_16183_));
 NAND2x1_ASAP7_75t_R _21591_ (.A(net343),
    .B(_00938_),
    .Y(_16184_));
 OA211x2_ASAP7_75t_R _21592_ (.A1(net343),
    .A2(_16183_),
    .B(_16184_),
    .C(net357),
    .Y(_16185_));
 OR3x1_ASAP7_75t_R _21593_ (.A(_13132_),
    .B(_16182_),
    .C(_16185_),
    .Y(_16186_));
 AND3x1_ASAP7_75t_R _21594_ (.A(_13598_),
    .B(_16179_),
    .C(_16186_),
    .Y(_16187_));
 INVx1_ASAP7_75t_R _21595_ (.A(_00933_),
    .Y(_16188_));
 NAND2x1_ASAP7_75t_R _21596_ (.A(net343),
    .B(_00931_),
    .Y(_16189_));
 OA211x2_ASAP7_75t_R _21597_ (.A1(net343),
    .A2(_16188_),
    .B(_16189_),
    .C(net311),
    .Y(_16190_));
 INVx1_ASAP7_75t_R _21598_ (.A(_00932_),
    .Y(_16191_));
 NAND2x1_ASAP7_75t_R _21599_ (.A(net343),
    .B(_00930_),
    .Y(_16192_));
 OA211x2_ASAP7_75t_R _21600_ (.A1(net343),
    .A2(_16191_),
    .B(_16192_),
    .C(net357),
    .Y(_16193_));
 OR3x1_ASAP7_75t_R _21601_ (.A(_13132_),
    .B(_16190_),
    .C(_16193_),
    .Y(_16194_));
 INVx1_ASAP7_75t_R _21602_ (.A(_00937_),
    .Y(_16195_));
 NAND2x1_ASAP7_75t_R _21603_ (.A(net343),
    .B(_00935_),
    .Y(_16196_));
 OA211x2_ASAP7_75t_R _21604_ (.A1(net343),
    .A2(_16195_),
    .B(_16196_),
    .C(net311),
    .Y(_16197_));
 INVx1_ASAP7_75t_R _21605_ (.A(_00936_),
    .Y(_16198_));
 NAND2x1_ASAP7_75t_R _21606_ (.A(net343),
    .B(_00934_),
    .Y(_16199_));
 OA211x2_ASAP7_75t_R _21607_ (.A1(net343),
    .A2(_16198_),
    .B(_16199_),
    .C(net357),
    .Y(_16200_));
 OR3x1_ASAP7_75t_R _21608_ (.A(net323),
    .B(_16197_),
    .C(_16200_),
    .Y(_16201_));
 AND3x1_ASAP7_75t_R _21609_ (.A(net317),
    .B(_16194_),
    .C(_16201_),
    .Y(_16202_));
 OR3x1_ASAP7_75t_R _21610_ (.A(net314),
    .B(_16187_),
    .C(_16202_),
    .Y(_16203_));
 OA21x2_ASAP7_75t_R _21611_ (.A1(_13174_),
    .A2(_16172_),
    .B(_16203_),
    .Y(_16204_));
 INVx3_ASAP7_75t_R _21612_ (.A(_16204_),
    .Y(_16205_));
 BUFx12f_ASAP7_75t_R max_cap250 (.A(_08287_),
    .Y(net250));
 OA21x2_ASAP7_75t_R _21614_ (.A1(_00280_),
    .A2(_14437_),
    .B(_13299_),
    .Y(_16207_));
 BUFx2_ASAP7_75t_R output249 (.A(net249),
    .Y(instr_req_o));
 OA21x2_ASAP7_75t_R _21616_ (.A1(net360),
    .A2(_15267_),
    .B(_16207_),
    .Y(_16209_));
 AO21x2_ASAP7_75t_R _21617_ (.A1(_13583_),
    .A2(_16205_),
    .B(_16209_),
    .Y(_18205_));
 INVx1_ASAP7_75t_R _21618_ (.A(_18205_),
    .Y(_18207_));
 AND2x2_ASAP7_75t_R _21619_ (.A(net395),
    .B(_01689_),
    .Y(_16210_));
 AO21x1_ASAP7_75t_R _21620_ (.A1(net302),
    .A2(_00917_),
    .B(_16210_),
    .Y(_16211_));
 OAI22x1_ASAP7_75t_R _21621_ (.A1(_00916_),
    .A2(_13471_),
    .B1(_16211_),
    .B2(net405),
    .Y(_16212_));
 NAND2x1_ASAP7_75t_R _21622_ (.A(net395),
    .B(_00923_),
    .Y(_16213_));
 OA211x2_ASAP7_75t_R _21623_ (.A1(net395),
    .A2(_16149_),
    .B(_16213_),
    .C(net305),
    .Y(_16214_));
 NAND2x1_ASAP7_75t_R _21624_ (.A(net395),
    .B(_00922_),
    .Y(_16215_));
 OA211x2_ASAP7_75t_R _21625_ (.A1(net395),
    .A2(_16152_),
    .B(_16215_),
    .C(net405),
    .Y(_16216_));
 OR3x1_ASAP7_75t_R _21626_ (.A(_14743_),
    .B(_16214_),
    .C(_16216_),
    .Y(_16217_));
 OA21x2_ASAP7_75t_R _21627_ (.A1(net300),
    .A2(_16212_),
    .B(_16217_),
    .Y(_16218_));
 NAND2x1_ASAP7_75t_R _21628_ (.A(net385),
    .B(_00919_),
    .Y(_16219_));
 OA211x2_ASAP7_75t_R _21629_ (.A1(net385),
    .A2(_16157_),
    .B(_16219_),
    .C(net305),
    .Y(_16220_));
 NAND2x1_ASAP7_75t_R _21630_ (.A(net385),
    .B(_00918_),
    .Y(_16221_));
 OA211x2_ASAP7_75t_R _21631_ (.A1(net385),
    .A2(_16160_),
    .B(_16221_),
    .C(net405),
    .Y(_16222_));
 OR3x1_ASAP7_75t_R _21632_ (.A(_13484_),
    .B(_16220_),
    .C(_16222_),
    .Y(_16223_));
 NAND2x1_ASAP7_75t_R _21633_ (.A(net385),
    .B(_00927_),
    .Y(_16224_));
 OA211x2_ASAP7_75t_R _21634_ (.A1(net385),
    .A2(_16164_),
    .B(_16224_),
    .C(net305),
    .Y(_16225_));
 NAND2x1_ASAP7_75t_R _21635_ (.A(net385),
    .B(_00926_),
    .Y(_16226_));
 OA211x2_ASAP7_75t_R _21636_ (.A1(net385),
    .A2(_16167_),
    .B(_16226_),
    .C(net405),
    .Y(_16227_));
 OR3x1_ASAP7_75t_R _21637_ (.A(net366),
    .B(_16225_),
    .C(_16227_),
    .Y(_16228_));
 AO21x1_ASAP7_75t_R _21638_ (.A1(_16223_),
    .A2(_16228_),
    .B(net373),
    .Y(_16229_));
 AO21x2_ASAP7_75t_R _21639_ (.A1(_16218_),
    .A2(_16229_),
    .B(_13392_),
    .Y(_16230_));
 NAND2x1_ASAP7_75t_R _21640_ (.A(net385),
    .B(_00942_),
    .Y(_16231_));
 OA211x2_ASAP7_75t_R _21641_ (.A1(net385),
    .A2(_16176_),
    .B(_16231_),
    .C(_13397_),
    .Y(_16232_));
 NAND2x1_ASAP7_75t_R _21642_ (.A(net385),
    .B(_00938_),
    .Y(_16233_));
 OA211x2_ASAP7_75t_R _21643_ (.A1(net385),
    .A2(_16183_),
    .B(_16233_),
    .C(net369),
    .Y(_16234_));
 OR3x1_ASAP7_75t_R _21644_ (.A(net305),
    .B(_16232_),
    .C(_16234_),
    .Y(_16235_));
 NAND2x1_ASAP7_75t_R _21645_ (.A(net385),
    .B(_00939_),
    .Y(_16236_));
 OA211x2_ASAP7_75t_R _21646_ (.A1(net385),
    .A2(_16180_),
    .B(_16236_),
    .C(net369),
    .Y(_16237_));
 NAND2x1_ASAP7_75t_R _21647_ (.A(net385),
    .B(_00943_),
    .Y(_16238_));
 OA211x2_ASAP7_75t_R _21648_ (.A1(net385),
    .A2(_16173_),
    .B(_16238_),
    .C(_13397_),
    .Y(_16239_));
 OR3x1_ASAP7_75t_R _21649_ (.A(net404),
    .B(_16237_),
    .C(_16239_),
    .Y(_16240_));
 AND3x1_ASAP7_75t_R _21650_ (.A(_13484_),
    .B(_16235_),
    .C(_16240_),
    .Y(_16241_));
 NAND2x1_ASAP7_75t_R _21651_ (.A(net369),
    .B(_00932_),
    .Y(_16242_));
 OA211x2_ASAP7_75t_R _21652_ (.A1(net369),
    .A2(_16198_),
    .B(_16242_),
    .C(net303),
    .Y(_16243_));
 INVx1_ASAP7_75t_R _21653_ (.A(_00934_),
    .Y(_16244_));
 NAND2x1_ASAP7_75t_R _21654_ (.A(net369),
    .B(_00930_),
    .Y(_16245_));
 OA211x2_ASAP7_75t_R _21655_ (.A1(net369),
    .A2(_16244_),
    .B(_16245_),
    .C(net387),
    .Y(_16246_));
 OR3x1_ASAP7_75t_R _21656_ (.A(net305),
    .B(_16243_),
    .C(_16246_),
    .Y(_16247_));
 NAND2x1_ASAP7_75t_R _21657_ (.A(net369),
    .B(_00933_),
    .Y(_16248_));
 OA211x2_ASAP7_75t_R _21658_ (.A1(net369),
    .A2(_16195_),
    .B(_16248_),
    .C(net303),
    .Y(_16249_));
 INVx1_ASAP7_75t_R _21659_ (.A(_00935_),
    .Y(_16250_));
 NAND2x1_ASAP7_75t_R _21660_ (.A(net369),
    .B(_00931_),
    .Y(_16251_));
 OA211x2_ASAP7_75t_R _21661_ (.A1(net369),
    .A2(_16250_),
    .B(_16251_),
    .C(net385),
    .Y(_16252_));
 OR3x1_ASAP7_75t_R _21662_ (.A(net404),
    .B(_16249_),
    .C(_16252_),
    .Y(_16253_));
 AND3x1_ASAP7_75t_R _21663_ (.A(net366),
    .B(_16247_),
    .C(_16253_),
    .Y(_16254_));
 OR3x4_ASAP7_75t_R _21664_ (.A(net363),
    .B(_16241_),
    .C(_16254_),
    .Y(_16255_));
 AND2x4_ASAP7_75t_R _21665_ (.A(_16230_),
    .B(_16255_),
    .Y(_16256_));
 BUFx2_ASAP7_75t_R output248 (.A(net248),
    .Y(instr_addr_o[9]));
 OAI22x1_ASAP7_75t_R _21667_ (.A1(_01621_),
    .A2(_13223_),
    .B1(_13880_),
    .B2(_00214_),
    .Y(_16258_));
 AO21x2_ASAP7_75t_R _21668_ (.A1(_13563_),
    .A2(_16256_),
    .B(_16258_),
    .Y(_16259_));
 BUFx2_ASAP7_75t_R output247 (.A(net247),
    .Y(instr_addr_o[8]));
 INVx2_ASAP7_75t_R _21670_ (.A(_16259_),
    .Y(_18206_));
 XOR2x2_ASAP7_75t_R _21671_ (.A(_00947_),
    .B(_02229_),
    .Y(_16260_));
 INVx4_ASAP7_75t_R _21672_ (.A(_16260_),
    .Y(net161));
 BUFx2_ASAP7_75t_R output246 (.A(net246),
    .Y(instr_addr_o[7]));
 INVx1_ASAP7_75t_R _21674_ (.A(_00958_),
    .Y(_16262_));
 NAND2x1_ASAP7_75t_R _21675_ (.A(net334),
    .B(_00956_),
    .Y(_16263_));
 OA211x2_ASAP7_75t_R _21676_ (.A1(net334),
    .A2(_16262_),
    .B(_16263_),
    .C(net308),
    .Y(_16264_));
 INVx1_ASAP7_75t_R _21677_ (.A(_00957_),
    .Y(_16265_));
 NAND2x1_ASAP7_75t_R _21678_ (.A(net334),
    .B(_00955_),
    .Y(_16266_));
 OA211x2_ASAP7_75t_R _21679_ (.A1(net334),
    .A2(_16265_),
    .B(_16266_),
    .C(net358),
    .Y(_16267_));
 OR3x1_ASAP7_75t_R _21680_ (.A(net319),
    .B(_16264_),
    .C(_16267_),
    .Y(_16268_));
 INVx1_ASAP7_75t_R _21681_ (.A(_00949_),
    .Y(_16269_));
 INVx1_ASAP7_75t_R _21682_ (.A(_00950_),
    .Y(_16270_));
 BUFx2_ASAP7_75t_R output245 (.A(net245),
    .Y(instr_addr_o[6]));
 NAND2x1_ASAP7_75t_R _21684_ (.A(net334),
    .B(_01688_),
    .Y(_16272_));
 OA21x2_ASAP7_75t_R _21685_ (.A1(net334),
    .A2(_16270_),
    .B(_16272_),
    .Y(_16273_));
 AO221x1_ASAP7_75t_R _21686_ (.A1(_16269_),
    .A2(_13190_),
    .B1(_16273_),
    .B2(net308),
    .C(_13598_),
    .Y(_16274_));
 AO21x1_ASAP7_75t_R _21687_ (.A1(_16268_),
    .A2(_16274_),
    .B(_13132_),
    .Y(_16275_));
 INVx1_ASAP7_75t_R _21688_ (.A(_00954_),
    .Y(_16276_));
 NAND2x1_ASAP7_75t_R _21689_ (.A(net337),
    .B(_00952_),
    .Y(_16277_));
 OA211x2_ASAP7_75t_R _21690_ (.A1(net337),
    .A2(_16276_),
    .B(_16277_),
    .C(_13145_),
    .Y(_16278_));
 INVx1_ASAP7_75t_R _21691_ (.A(_00953_),
    .Y(_16279_));
 NAND2x1_ASAP7_75t_R _21692_ (.A(net337),
    .B(_00951_),
    .Y(_16280_));
 OA211x2_ASAP7_75t_R _21693_ (.A1(net337),
    .A2(_16279_),
    .B(_16280_),
    .C(net358),
    .Y(_16281_));
 OR3x1_ASAP7_75t_R _21694_ (.A(_13598_),
    .B(_16278_),
    .C(_16281_),
    .Y(_16282_));
 INVx1_ASAP7_75t_R _21695_ (.A(_00962_),
    .Y(_16283_));
 NAND2x1_ASAP7_75t_R _21696_ (.A(net337),
    .B(_00960_),
    .Y(_16284_));
 OA211x2_ASAP7_75t_R _21697_ (.A1(net337),
    .A2(_16283_),
    .B(_16284_),
    .C(_13145_),
    .Y(_16285_));
 BUFx2_ASAP7_75t_R output244 (.A(net244),
    .Y(instr_addr_o[5]));
 INVx1_ASAP7_75t_R _21699_ (.A(_00961_),
    .Y(_16287_));
 NAND2x1_ASAP7_75t_R _21700_ (.A(net337),
    .B(_00959_),
    .Y(_16288_));
 OA211x2_ASAP7_75t_R _21701_ (.A1(net337),
    .A2(_16287_),
    .B(_16288_),
    .C(net358),
    .Y(_16289_));
 OR3x1_ASAP7_75t_R _21702_ (.A(net319),
    .B(_16285_),
    .C(_16289_),
    .Y(_16290_));
 AO21x1_ASAP7_75t_R _21703_ (.A1(_16282_),
    .A2(_16290_),
    .B(net325),
    .Y(_16291_));
 AO21x1_ASAP7_75t_R _21704_ (.A1(_16275_),
    .A2(_16291_),
    .B(_13174_),
    .Y(_16292_));
 INVx1_ASAP7_75t_R _21705_ (.A(_00970_),
    .Y(_16293_));
 NAND2x1_ASAP7_75t_R _21706_ (.A(net334),
    .B(_00968_),
    .Y(_16294_));
 OA211x2_ASAP7_75t_R _21707_ (.A1(net334),
    .A2(_16293_),
    .B(_16294_),
    .C(_13145_),
    .Y(_16295_));
 INVx1_ASAP7_75t_R _21708_ (.A(_00969_),
    .Y(_16296_));
 NAND2x1_ASAP7_75t_R _21709_ (.A(net334),
    .B(_00967_),
    .Y(_16297_));
 OA211x2_ASAP7_75t_R _21710_ (.A1(net334),
    .A2(_16296_),
    .B(_16297_),
    .C(net358),
    .Y(_16298_));
 OR3x1_ASAP7_75t_R _21711_ (.A(_13598_),
    .B(_16295_),
    .C(_16298_),
    .Y(_16299_));
 INVx1_ASAP7_75t_R _21712_ (.A(_00978_),
    .Y(_16300_));
 NAND2x1_ASAP7_75t_R _21713_ (.A(net334),
    .B(_00976_),
    .Y(_16301_));
 OA211x2_ASAP7_75t_R _21714_ (.A1(net334),
    .A2(_16300_),
    .B(_16301_),
    .C(_13145_),
    .Y(_16302_));
 INVx1_ASAP7_75t_R _21715_ (.A(_00977_),
    .Y(_16303_));
 NAND2x1_ASAP7_75t_R _21716_ (.A(net334),
    .B(_00975_),
    .Y(_16304_));
 OA211x2_ASAP7_75t_R _21717_ (.A1(net334),
    .A2(_16303_),
    .B(_16304_),
    .C(net358),
    .Y(_16305_));
 OR3x1_ASAP7_75t_R _21718_ (.A(net318),
    .B(_16302_),
    .C(_16305_),
    .Y(_16306_));
 AND3x1_ASAP7_75t_R _21719_ (.A(_13132_),
    .B(_16299_),
    .C(_16306_),
    .Y(_16307_));
 INVx1_ASAP7_75t_R _21720_ (.A(_00966_),
    .Y(_16308_));
 NAND2x1_ASAP7_75t_R _21721_ (.A(net337),
    .B(_00964_),
    .Y(_16309_));
 OA211x2_ASAP7_75t_R _21722_ (.A1(net337),
    .A2(_16308_),
    .B(_16309_),
    .C(_13145_),
    .Y(_16310_));
 INVx1_ASAP7_75t_R _21723_ (.A(_00965_),
    .Y(_16311_));
 NAND2x1_ASAP7_75t_R _21724_ (.A(net337),
    .B(_00963_),
    .Y(_16312_));
 OA211x2_ASAP7_75t_R _21725_ (.A1(net337),
    .A2(_16311_),
    .B(_16312_),
    .C(net358),
    .Y(_16313_));
 OR3x1_ASAP7_75t_R _21726_ (.A(_13598_),
    .B(_16310_),
    .C(_16313_),
    .Y(_16314_));
 INVx1_ASAP7_75t_R _21727_ (.A(_00974_),
    .Y(_16315_));
 NAND2x1_ASAP7_75t_R _21728_ (.A(net337),
    .B(_00972_),
    .Y(_16316_));
 OA211x2_ASAP7_75t_R _21729_ (.A1(net337),
    .A2(_16315_),
    .B(_16316_),
    .C(_13145_),
    .Y(_16317_));
 INVx1_ASAP7_75t_R _21730_ (.A(_00973_),
    .Y(_16318_));
 NAND2x1_ASAP7_75t_R _21731_ (.A(net337),
    .B(_00971_),
    .Y(_16319_));
 OA211x2_ASAP7_75t_R _21732_ (.A1(net337),
    .A2(_16318_),
    .B(_16319_),
    .C(net358),
    .Y(_16320_));
 OR3x1_ASAP7_75t_R _21733_ (.A(net318),
    .B(_16317_),
    .C(_16320_),
    .Y(_16321_));
 AND3x1_ASAP7_75t_R _21734_ (.A(net325),
    .B(_16314_),
    .C(_16321_),
    .Y(_16322_));
 OR3x4_ASAP7_75t_R _21735_ (.A(net315),
    .B(_16307_),
    .C(_16322_),
    .Y(_16323_));
 NAND2x2_ASAP7_75t_R _21736_ (.A(_16292_),
    .B(_16323_),
    .Y(_16324_));
 OA21x2_ASAP7_75t_R _21737_ (.A1(_01745_),
    .A2(_15267_),
    .B(_16207_),
    .Y(_16325_));
 AO21x2_ASAP7_75t_R _21738_ (.A1(_13583_),
    .A2(_16324_),
    .B(_16325_),
    .Y(_16326_));
 BUFx2_ASAP7_75t_R output243 (.A(net243),
    .Y(instr_addr_o[4]));
 INVx1_ASAP7_75t_R _21740_ (.A(_16326_),
    .Y(_18212_));
 INVx2_ASAP7_75t_R _21741_ (.A(_00215_),
    .Y(\cs_registers_i.pc_id_i[21] ));
 NOR2x1_ASAP7_75t_R _21742_ (.A(_01620_),
    .B(_13223_),
    .Y(_16327_));
 AOI21x1_ASAP7_75t_R _21743_ (.A1(_00215_),
    .A2(_13553_),
    .B(_13561_),
    .Y(_16328_));
 NAND2x1_ASAP7_75t_R _21744_ (.A(net396),
    .B(_00968_),
    .Y(_16329_));
 OA211x2_ASAP7_75t_R _21745_ (.A1(net396),
    .A2(_16293_),
    .B(_16329_),
    .C(_13424_),
    .Y(_16330_));
 NAND2x1_ASAP7_75t_R _21746_ (.A(net396),
    .B(_00967_),
    .Y(_16331_));
 OA211x2_ASAP7_75t_R _21747_ (.A1(net396),
    .A2(_16296_),
    .B(_16331_),
    .C(net408),
    .Y(_16332_));
 OR3x1_ASAP7_75t_R _21748_ (.A(net372),
    .B(_16330_),
    .C(_16332_),
    .Y(_16333_));
 NAND2x1_ASAP7_75t_R _21749_ (.A(net396),
    .B(_00964_),
    .Y(_16334_));
 OA211x2_ASAP7_75t_R _21750_ (.A1(net396),
    .A2(_16308_),
    .B(_16334_),
    .C(_13424_),
    .Y(_16335_));
 NAND2x1_ASAP7_75t_R _21751_ (.A(net396),
    .B(_00963_),
    .Y(_16336_));
 OA211x2_ASAP7_75t_R _21752_ (.A1(net396),
    .A2(_16311_),
    .B(_16336_),
    .C(net408),
    .Y(_16337_));
 OR3x1_ASAP7_75t_R _21753_ (.A(_13397_),
    .B(_16335_),
    .C(_16337_),
    .Y(_16338_));
 NAND2x1_ASAP7_75t_R _21754_ (.A(net396),
    .B(_00951_),
    .Y(_16339_));
 OA211x2_ASAP7_75t_R _21755_ (.A1(net396),
    .A2(_16279_),
    .B(_16339_),
    .C(net408),
    .Y(_16340_));
 NAND2x1_ASAP7_75t_R _21756_ (.A(net396),
    .B(_00952_),
    .Y(_16341_));
 OA211x2_ASAP7_75t_R _21757_ (.A1(net396),
    .A2(_16276_),
    .B(_16341_),
    .C(net306),
    .Y(_16342_));
 OR3x1_ASAP7_75t_R _21758_ (.A(_13814_),
    .B(_16340_),
    .C(_16342_),
    .Y(_16343_));
 NAND2x1_ASAP7_75t_R _21759_ (.A(net394),
    .B(_01688_),
    .Y(_16344_));
 OA211x2_ASAP7_75t_R _21760_ (.A1(net394),
    .A2(_16270_),
    .B(_16344_),
    .C(net306),
    .Y(_16345_));
 AND3x1_ASAP7_75t_R _21761_ (.A(net408),
    .B(net302),
    .C(_16269_),
    .Y(_16346_));
 OA31x2_ASAP7_75t_R _21762_ (.A1(_13828_),
    .A2(_16345_),
    .A3(_16346_),
    .B1(net364),
    .Y(_16347_));
 AO32x1_ASAP7_75t_R _21763_ (.A1(_13392_),
    .A2(_16333_),
    .A3(_16338_),
    .B1(_16343_),
    .B2(_16347_),
    .Y(_16348_));
 NAND2x1_ASAP7_75t_R _21764_ (.A(net396),
    .B(_00960_),
    .Y(_16349_));
 OA211x2_ASAP7_75t_R _21765_ (.A1(net396),
    .A2(_16283_),
    .B(_16349_),
    .C(net306),
    .Y(_16350_));
 NAND2x1_ASAP7_75t_R _21766_ (.A(net396),
    .B(_00959_),
    .Y(_16351_));
 OA211x2_ASAP7_75t_R _21767_ (.A1(net396),
    .A2(_16287_),
    .B(_16351_),
    .C(net410),
    .Y(_16352_));
 OR3x1_ASAP7_75t_R _21768_ (.A(net371),
    .B(_16350_),
    .C(_16352_),
    .Y(_16353_));
 NAND2x1_ASAP7_75t_R _21769_ (.A(net394),
    .B(_00956_),
    .Y(_16354_));
 OA211x2_ASAP7_75t_R _21770_ (.A1(net394),
    .A2(_16262_),
    .B(_16354_),
    .C(net306),
    .Y(_16355_));
 NAND2x1_ASAP7_75t_R _21771_ (.A(net394),
    .B(_00955_),
    .Y(_16356_));
 OA211x2_ASAP7_75t_R _21772_ (.A1(net394),
    .A2(_16265_),
    .B(_16356_),
    .C(net408),
    .Y(_16357_));
 OR3x1_ASAP7_75t_R _21773_ (.A(_13397_),
    .B(_16355_),
    .C(_16357_),
    .Y(_16358_));
 AND2x2_ASAP7_75t_R _21774_ (.A(_16353_),
    .B(_16358_),
    .Y(_16359_));
 AND2x2_ASAP7_75t_R _21775_ (.A(_16343_),
    .B(_16347_),
    .Y(_16360_));
 NAND2x1_ASAP7_75t_R _21776_ (.A(net396),
    .B(_00972_),
    .Y(_16361_));
 OA211x2_ASAP7_75t_R _21777_ (.A1(net396),
    .A2(_16315_),
    .B(_16361_),
    .C(_13424_),
    .Y(_16362_));
 NAND2x1_ASAP7_75t_R _21778_ (.A(net396),
    .B(_00971_),
    .Y(_16363_));
 OA211x2_ASAP7_75t_R _21779_ (.A1(net396),
    .A2(_16318_),
    .B(_16363_),
    .C(net408),
    .Y(_16364_));
 OR3x1_ASAP7_75t_R _21780_ (.A(_13397_),
    .B(_16362_),
    .C(_16364_),
    .Y(_16365_));
 NAND2x1_ASAP7_75t_R _21781_ (.A(net396),
    .B(_00976_),
    .Y(_16366_));
 OA211x2_ASAP7_75t_R _21782_ (.A1(net396),
    .A2(_16300_),
    .B(_16366_),
    .C(_13424_),
    .Y(_16367_));
 NAND2x1_ASAP7_75t_R _21783_ (.A(net396),
    .B(_00975_),
    .Y(_16368_));
 OA211x2_ASAP7_75t_R _21784_ (.A1(net396),
    .A2(_16303_),
    .B(_16368_),
    .C(net408),
    .Y(_16369_));
 OR3x1_ASAP7_75t_R _21785_ (.A(net372),
    .B(_16367_),
    .C(_16369_),
    .Y(_16370_));
 AND3x1_ASAP7_75t_R _21786_ (.A(_14571_),
    .B(_16365_),
    .C(_16370_),
    .Y(_16371_));
 AO221x2_ASAP7_75t_R _21787_ (.A1(net365),
    .A2(_16348_),
    .B1(_16359_),
    .B2(_16360_),
    .C(_16371_),
    .Y(_16372_));
 OAI22x1_ASAP7_75t_R _21788_ (.A1(_16327_),
    .A2(_16328_),
    .B1(_16372_),
    .B2(_13782_),
    .Y(_18211_));
 AND2x2_ASAP7_75t_R _21789_ (.A(net330),
    .B(_01687_),
    .Y(_16373_));
 AO21x1_ASAP7_75t_R _21790_ (.A1(net312),
    .A2(_00982_),
    .B(_16373_),
    .Y(_16374_));
 OAI22x1_ASAP7_75t_R _21791_ (.A1(_00981_),
    .A2(_13586_),
    .B1(_16374_),
    .B2(net361),
    .Y(_16375_));
 INVx1_ASAP7_75t_R _21792_ (.A(_00990_),
    .Y(_16376_));
 NAND2x1_ASAP7_75t_R _21793_ (.A(net330),
    .B(_00988_),
    .Y(_16377_));
 OA211x2_ASAP7_75t_R _21794_ (.A1(net330),
    .A2(_16376_),
    .B(_16377_),
    .C(net310),
    .Y(_16378_));
 INVx1_ASAP7_75t_R _21795_ (.A(_00989_),
    .Y(_16379_));
 NAND2x1_ASAP7_75t_R _21796_ (.A(net330),
    .B(_00987_),
    .Y(_16380_));
 OA211x2_ASAP7_75t_R _21797_ (.A1(net330),
    .A2(_16379_),
    .B(_16380_),
    .C(net354),
    .Y(_16381_));
 OR3x1_ASAP7_75t_R _21798_ (.A(net321),
    .B(_16378_),
    .C(_16381_),
    .Y(_16382_));
 OA211x2_ASAP7_75t_R _21799_ (.A1(_13598_),
    .A2(_16375_),
    .B(_16382_),
    .C(net322),
    .Y(_16383_));
 INVx1_ASAP7_75t_R _21800_ (.A(_00986_),
    .Y(_16384_));
 NAND2x1_ASAP7_75t_R _21801_ (.A(net326),
    .B(_00984_),
    .Y(_16385_));
 OA211x2_ASAP7_75t_R _21802_ (.A1(net326),
    .A2(_16384_),
    .B(_16385_),
    .C(net310),
    .Y(_16386_));
 INVx1_ASAP7_75t_R _21803_ (.A(_00985_),
    .Y(_16387_));
 NAND2x1_ASAP7_75t_R _21804_ (.A(net326),
    .B(_00983_),
    .Y(_16388_));
 OA211x2_ASAP7_75t_R _21805_ (.A1(net326),
    .A2(_16387_),
    .B(_16388_),
    .C(_00246_),
    .Y(_16389_));
 OR3x1_ASAP7_75t_R _21806_ (.A(_13598_),
    .B(_16386_),
    .C(_16389_),
    .Y(_16390_));
 INVx1_ASAP7_75t_R _21807_ (.A(_00994_),
    .Y(_16391_));
 NAND2x1_ASAP7_75t_R _21808_ (.A(net326),
    .B(_00992_),
    .Y(_16392_));
 OA211x2_ASAP7_75t_R _21809_ (.A1(net326),
    .A2(_16391_),
    .B(_16392_),
    .C(net310),
    .Y(_16393_));
 INVx1_ASAP7_75t_R _21810_ (.A(_00993_),
    .Y(_16394_));
 NAND2x1_ASAP7_75t_R _21811_ (.A(net326),
    .B(_00991_),
    .Y(_16395_));
 OA211x2_ASAP7_75t_R _21812_ (.A1(net326),
    .A2(_16394_),
    .B(_16395_),
    .C(_00246_),
    .Y(_16396_));
 OR3x1_ASAP7_75t_R _21813_ (.A(net321),
    .B(_16393_),
    .C(_16396_),
    .Y(_16397_));
 AND3x1_ASAP7_75t_R _21814_ (.A(_13132_),
    .B(_16390_),
    .C(_16397_),
    .Y(_16398_));
 OR3x4_ASAP7_75t_R _21815_ (.A(_13174_),
    .B(_16383_),
    .C(_16398_),
    .Y(_16399_));
 INVx1_ASAP7_75t_R _21816_ (.A(_01002_),
    .Y(_16400_));
 NAND2x1_ASAP7_75t_R _21817_ (.A(net329),
    .B(_01000_),
    .Y(_16401_));
 OA211x2_ASAP7_75t_R _21818_ (.A1(net329),
    .A2(_16400_),
    .B(_16401_),
    .C(net310),
    .Y(_16402_));
 INVx1_ASAP7_75t_R _21819_ (.A(_01001_),
    .Y(_16403_));
 BUFx2_ASAP7_75t_R output242 (.A(net242),
    .Y(instr_addr_o[3]));
 NAND2x1_ASAP7_75t_R _21821_ (.A(net329),
    .B(_00999_),
    .Y(_16405_));
 OA211x2_ASAP7_75t_R _21822_ (.A1(net329),
    .A2(_16403_),
    .B(_16405_),
    .C(net354),
    .Y(_16406_));
 OR3x1_ASAP7_75t_R _21823_ (.A(net322),
    .B(_16402_),
    .C(_16406_),
    .Y(_16407_));
 INVx1_ASAP7_75t_R _21824_ (.A(_00998_),
    .Y(_16408_));
 NAND2x1_ASAP7_75t_R _21825_ (.A(net330),
    .B(_00996_),
    .Y(_16409_));
 OA211x2_ASAP7_75t_R _21826_ (.A1(net330),
    .A2(_16408_),
    .B(_16409_),
    .C(net310),
    .Y(_16410_));
 INVx1_ASAP7_75t_R _21827_ (.A(_00997_),
    .Y(_16411_));
 NAND2x1_ASAP7_75t_R _21828_ (.A(net330),
    .B(_00995_),
    .Y(_16412_));
 OA211x2_ASAP7_75t_R _21829_ (.A1(net330),
    .A2(_16411_),
    .B(_16412_),
    .C(net361),
    .Y(_16413_));
 OR3x1_ASAP7_75t_R _21830_ (.A(_13132_),
    .B(_16410_),
    .C(_16413_),
    .Y(_16414_));
 AND3x1_ASAP7_75t_R _21831_ (.A(net321),
    .B(_16407_),
    .C(_16414_),
    .Y(_16415_));
 INVx1_ASAP7_75t_R _21832_ (.A(_01010_),
    .Y(_16416_));
 NAND2x1_ASAP7_75t_R _21833_ (.A(net330),
    .B(_01008_),
    .Y(_16417_));
 OA211x2_ASAP7_75t_R _21834_ (.A1(net330),
    .A2(_16416_),
    .B(_16417_),
    .C(net310),
    .Y(_16418_));
 BUFx2_ASAP7_75t_R output241 (.A(net241),
    .Y(instr_addr_o[31]));
 INVx1_ASAP7_75t_R _21836_ (.A(_01009_),
    .Y(_16420_));
 NAND2x1_ASAP7_75t_R _21837_ (.A(net330),
    .B(_01007_),
    .Y(_16421_));
 OA211x2_ASAP7_75t_R _21838_ (.A1(net330),
    .A2(_16420_),
    .B(_16421_),
    .C(net354),
    .Y(_16422_));
 OR3x1_ASAP7_75t_R _21839_ (.A(net322),
    .B(_16418_),
    .C(_16422_),
    .Y(_16423_));
 INVx1_ASAP7_75t_R _21840_ (.A(_01006_),
    .Y(_16424_));
 NAND2x1_ASAP7_75t_R _21841_ (.A(net330),
    .B(_01004_),
    .Y(_16425_));
 OA211x2_ASAP7_75t_R _21842_ (.A1(net330),
    .A2(_16424_),
    .B(_16425_),
    .C(net310),
    .Y(_16426_));
 INVx1_ASAP7_75t_R _21843_ (.A(_01005_),
    .Y(_16427_));
 NAND2x1_ASAP7_75t_R _21844_ (.A(net330),
    .B(_01003_),
    .Y(_16428_));
 OA211x2_ASAP7_75t_R _21845_ (.A1(net330),
    .A2(_16427_),
    .B(_16428_),
    .C(net354),
    .Y(_16429_));
 OR3x1_ASAP7_75t_R _21846_ (.A(_13132_),
    .B(_16426_),
    .C(_16429_),
    .Y(_16430_));
 AND3x1_ASAP7_75t_R _21847_ (.A(_13598_),
    .B(_16423_),
    .C(_16430_),
    .Y(_16431_));
 OR3x4_ASAP7_75t_R _21848_ (.A(net316),
    .B(_16415_),
    .C(_16431_),
    .Y(_16432_));
 NAND2x2_ASAP7_75t_R _21849_ (.A(_16399_),
    .B(_16432_),
    .Y(_16433_));
 OA21x2_ASAP7_75t_R _21850_ (.A1(_01744_),
    .A2(_15267_),
    .B(_16207_),
    .Y(_16434_));
 AO21x2_ASAP7_75t_R _21851_ (.A1(_13583_),
    .A2(_16433_),
    .B(_16434_),
    .Y(_18218_));
 INVx1_ASAP7_75t_R _21852_ (.A(_18218_),
    .Y(_18216_));
 AND2x2_ASAP7_75t_R _21853_ (.A(_00217_),
    .B(_13553_),
    .Y(_16435_));
 NAND2x1_ASAP7_75t_R _21854_ (.A(net377),
    .B(_00984_),
    .Y(_16436_));
 OA211x2_ASAP7_75t_R _21855_ (.A1(net377),
    .A2(_16384_),
    .B(_16436_),
    .C(net304),
    .Y(_16437_));
 NAND2x1_ASAP7_75t_R _21856_ (.A(net377),
    .B(_00983_),
    .Y(_16438_));
 OA211x2_ASAP7_75t_R _21857_ (.A1(net377),
    .A2(_16387_),
    .B(_16438_),
    .C(net412),
    .Y(_16439_));
 OR3x1_ASAP7_75t_R _21858_ (.A(_13484_),
    .B(_16437_),
    .C(_16439_),
    .Y(_16440_));
 NAND2x1_ASAP7_75t_R _21859_ (.A(net377),
    .B(_00992_),
    .Y(_16441_));
 OA211x2_ASAP7_75t_R _21860_ (.A1(net377),
    .A2(_16391_),
    .B(_16441_),
    .C(net304),
    .Y(_16442_));
 NAND2x1_ASAP7_75t_R _21861_ (.A(net379),
    .B(_00991_),
    .Y(_16443_));
 OA211x2_ASAP7_75t_R _21862_ (.A1(net377),
    .A2(_16394_),
    .B(_16443_),
    .C(net412),
    .Y(_16444_));
 OR3x1_ASAP7_75t_R _21863_ (.A(net368),
    .B(_16442_),
    .C(_16444_),
    .Y(_16445_));
 AO21x1_ASAP7_75t_R _21864_ (.A1(_16440_),
    .A2(_16445_),
    .B(net375),
    .Y(_16446_));
 AND2x2_ASAP7_75t_R _21865_ (.A(net384),
    .B(_01687_),
    .Y(_16447_));
 AO21x1_ASAP7_75t_R _21866_ (.A1(net303),
    .A2(_00982_),
    .B(_16447_),
    .Y(_16448_));
 OAI22x1_ASAP7_75t_R _21867_ (.A1(_00981_),
    .A2(_13471_),
    .B1(_16448_),
    .B2(net412),
    .Y(_16449_));
 NAND2x1_ASAP7_75t_R _21868_ (.A(net378),
    .B(_00987_),
    .Y(_16450_));
 OA211x2_ASAP7_75t_R _21869_ (.A1(net378),
    .A2(_16379_),
    .B(_16450_),
    .C(net412),
    .Y(_16451_));
 NAND2x1_ASAP7_75t_R _21870_ (.A(net378),
    .B(_00988_),
    .Y(_16452_));
 OA211x2_ASAP7_75t_R _21871_ (.A1(net378),
    .A2(_16376_),
    .B(_16452_),
    .C(net304),
    .Y(_16453_));
 OR3x1_ASAP7_75t_R _21872_ (.A(_14743_),
    .B(_16451_),
    .C(_16453_),
    .Y(_16454_));
 OA211x2_ASAP7_75t_R _21873_ (.A1(net301),
    .A2(_16449_),
    .B(_16454_),
    .C(net363),
    .Y(_16455_));
 NAND2x1_ASAP7_75t_R _21874_ (.A(net376),
    .B(_01004_),
    .Y(_16456_));
 OA211x2_ASAP7_75t_R _21875_ (.A1(net376),
    .A2(_16424_),
    .B(_16456_),
    .C(net304),
    .Y(_16457_));
 NAND2x1_ASAP7_75t_R _21876_ (.A(net376),
    .B(_01003_),
    .Y(_16458_));
 OA211x2_ASAP7_75t_R _21877_ (.A1(net376),
    .A2(_16427_),
    .B(_16458_),
    .C(net406),
    .Y(_16459_));
 OR3x1_ASAP7_75t_R _21878_ (.A(_13397_),
    .B(_16457_),
    .C(_16459_),
    .Y(_16460_));
 NAND2x1_ASAP7_75t_R _21879_ (.A(net378),
    .B(_01008_),
    .Y(_16461_));
 OA211x2_ASAP7_75t_R _21880_ (.A1(net378),
    .A2(_16416_),
    .B(_16461_),
    .C(net304),
    .Y(_16462_));
 NAND2x1_ASAP7_75t_R _21881_ (.A(net376),
    .B(_01007_),
    .Y(_16463_));
 OA211x2_ASAP7_75t_R _21882_ (.A1(net376),
    .A2(_16420_),
    .B(_16463_),
    .C(net406),
    .Y(_16464_));
 OR3x1_ASAP7_75t_R _21883_ (.A(net374),
    .B(_16462_),
    .C(_16464_),
    .Y(_16465_));
 AO21x1_ASAP7_75t_R _21884_ (.A1(_16460_),
    .A2(_16465_),
    .B(net368),
    .Y(_16466_));
 NAND2x1_ASAP7_75t_R _21885_ (.A(net376),
    .B(_00999_),
    .Y(_16467_));
 OA211x2_ASAP7_75t_R _21886_ (.A1(net376),
    .A2(_16403_),
    .B(_16467_),
    .C(net406),
    .Y(_16468_));
 NAND2x1_ASAP7_75t_R _21887_ (.A(net376),
    .B(_01000_),
    .Y(_16469_));
 OA211x2_ASAP7_75t_R _21888_ (.A1(net376),
    .A2(_16400_),
    .B(_16469_),
    .C(net304),
    .Y(_16470_));
 OR3x1_ASAP7_75t_R _21889_ (.A(net298),
    .B(_16468_),
    .C(_16470_),
    .Y(_16471_));
 NAND2x1_ASAP7_75t_R _21890_ (.A(net384),
    .B(_00996_),
    .Y(_16472_));
 OA211x2_ASAP7_75t_R _21891_ (.A1(net384),
    .A2(_16408_),
    .B(_16472_),
    .C(net304),
    .Y(_16473_));
 NAND2x1_ASAP7_75t_R _21892_ (.A(net384),
    .B(_00995_),
    .Y(_16474_));
 OA211x2_ASAP7_75t_R _21893_ (.A1(net384),
    .A2(_16411_),
    .B(_16474_),
    .C(net412),
    .Y(_16475_));
 OR3x1_ASAP7_75t_R _21894_ (.A(net301),
    .B(_16473_),
    .C(_16475_),
    .Y(_16476_));
 AND3x1_ASAP7_75t_R _21895_ (.A(_13392_),
    .B(_16471_),
    .C(_16476_),
    .Y(_16477_));
 AOI221x1_ASAP7_75t_R _21896_ (.A1(_16446_),
    .A2(_16455_),
    .B1(_16466_),
    .B2(_16477_),
    .C(_13553_),
    .Y(_16478_));
 AO21x1_ASAP7_75t_R _21897_ (.A1(_13219_),
    .A2(_13222_),
    .B(_01619_),
    .Y(_16479_));
 OA31x2_ASAP7_75t_R _21898_ (.A1(_13561_),
    .A2(_16435_),
    .A3(_16478_),
    .B1(_16479_),
    .Y(_16480_));
 BUFx2_ASAP7_75t_R output240 (.A(net240),
    .Y(instr_addr_o[30]));
 XOR2x2_ASAP7_75t_R _21900_ (.A(_01014_),
    .B(_01012_),
    .Y(net163));
 AND2x2_ASAP7_75t_R _21901_ (.A(net339),
    .B(_01686_),
    .Y(_16481_));
 AO21x1_ASAP7_75t_R _21902_ (.A1(net313),
    .A2(_01016_),
    .B(_16481_),
    .Y(_16482_));
 OAI22x1_ASAP7_75t_R _21903_ (.A1(_01015_),
    .A2(_13586_),
    .B1(_16482_),
    .B2(net359),
    .Y(_16483_));
 INVx1_ASAP7_75t_R _21904_ (.A(_01024_),
    .Y(_16484_));
 NAND2x1_ASAP7_75t_R _21905_ (.A(net338),
    .B(_01022_),
    .Y(_16485_));
 OA211x2_ASAP7_75t_R _21906_ (.A1(net338),
    .A2(_16484_),
    .B(_16485_),
    .C(net308),
    .Y(_16486_));
 INVx1_ASAP7_75t_R _21907_ (.A(_01023_),
    .Y(_16487_));
 NAND2x1_ASAP7_75t_R _21908_ (.A(net338),
    .B(_01021_),
    .Y(_16488_));
 OA211x2_ASAP7_75t_R _21909_ (.A1(net338),
    .A2(_16487_),
    .B(_16488_),
    .C(net359),
    .Y(_16489_));
 OR3x1_ASAP7_75t_R _21910_ (.A(net319),
    .B(_16486_),
    .C(_16489_),
    .Y(_16490_));
 OA21x2_ASAP7_75t_R _21911_ (.A1(_13598_),
    .A2(_16483_),
    .B(_16490_),
    .Y(_16491_));
 INVx1_ASAP7_75t_R _21912_ (.A(_01020_),
    .Y(_16492_));
 NAND2x1_ASAP7_75t_R _21913_ (.A(net339),
    .B(_01018_),
    .Y(_16493_));
 OA211x2_ASAP7_75t_R _21914_ (.A1(net339),
    .A2(_16492_),
    .B(_16493_),
    .C(net309),
    .Y(_16494_));
 INVx1_ASAP7_75t_R _21915_ (.A(_01019_),
    .Y(_16495_));
 NAND2x1_ASAP7_75t_R _21916_ (.A(net340),
    .B(_01017_),
    .Y(_04504_));
 OA211x2_ASAP7_75t_R _21917_ (.A1(net339),
    .A2(_16495_),
    .B(_04504_),
    .C(net359),
    .Y(_04505_));
 OR3x1_ASAP7_75t_R _21918_ (.A(_13598_),
    .B(_16494_),
    .C(_04505_),
    .Y(_04506_));
 INVx1_ASAP7_75t_R _21919_ (.A(_01028_),
    .Y(_04507_));
 NAND2x1_ASAP7_75t_R _21920_ (.A(net338),
    .B(_01026_),
    .Y(_04508_));
 OA211x2_ASAP7_75t_R _21921_ (.A1(net338),
    .A2(_04507_),
    .B(_04508_),
    .C(net308),
    .Y(_04509_));
 INVx1_ASAP7_75t_R _21922_ (.A(_01027_),
    .Y(_04510_));
 NAND2x1_ASAP7_75t_R _21923_ (.A(net338),
    .B(_01025_),
    .Y(_04511_));
 OA211x2_ASAP7_75t_R _21924_ (.A1(net339),
    .A2(_04510_),
    .B(_04511_),
    .C(net359),
    .Y(_04512_));
 OR3x1_ASAP7_75t_R _21925_ (.A(net319),
    .B(_04509_),
    .C(_04512_),
    .Y(_04513_));
 AND3x1_ASAP7_75t_R _21926_ (.A(_13132_),
    .B(_04506_),
    .C(_04513_),
    .Y(_04514_));
 AO21x1_ASAP7_75t_R _21927_ (.A1(_01744_),
    .A2(_16491_),
    .B(_04514_),
    .Y(_04515_));
 INVx1_ASAP7_75t_R _21928_ (.A(_01036_),
    .Y(_04516_));
 NAND2x1_ASAP7_75t_R _21929_ (.A(net339),
    .B(_01034_),
    .Y(_04517_));
 OA211x2_ASAP7_75t_R _21930_ (.A1(net339),
    .A2(_04516_),
    .B(_04517_),
    .C(net308),
    .Y(_04518_));
 INVx1_ASAP7_75t_R _21931_ (.A(_01035_),
    .Y(_04519_));
 NAND2x1_ASAP7_75t_R _21932_ (.A(net339),
    .B(_01033_),
    .Y(_04520_));
 OA211x2_ASAP7_75t_R _21933_ (.A1(net339),
    .A2(_04519_),
    .B(_04520_),
    .C(net359),
    .Y(_04521_));
 OR3x1_ASAP7_75t_R _21934_ (.A(_13598_),
    .B(_04518_),
    .C(_04521_),
    .Y(_04522_));
 INVx1_ASAP7_75t_R _21935_ (.A(_01044_),
    .Y(_04523_));
 NAND2x1_ASAP7_75t_R _21936_ (.A(net339),
    .B(_01042_),
    .Y(_04524_));
 OA211x2_ASAP7_75t_R _21937_ (.A1(net339),
    .A2(_04523_),
    .B(_04524_),
    .C(net308),
    .Y(_04525_));
 INVx1_ASAP7_75t_R _21938_ (.A(_01043_),
    .Y(_04526_));
 NAND2x1_ASAP7_75t_R _21939_ (.A(net339),
    .B(_01041_),
    .Y(_04527_));
 OA211x2_ASAP7_75t_R _21940_ (.A1(net339),
    .A2(_04526_),
    .B(_04527_),
    .C(net359),
    .Y(_04528_));
 OR3x1_ASAP7_75t_R _21941_ (.A(net319),
    .B(_04525_),
    .C(_04528_),
    .Y(_04529_));
 AND3x1_ASAP7_75t_R _21942_ (.A(_13132_),
    .B(_04522_),
    .C(_04529_),
    .Y(_04530_));
 INVx1_ASAP7_75t_R _21943_ (.A(_01032_),
    .Y(_04531_));
 NAND2x1_ASAP7_75t_R _21944_ (.A(net339),
    .B(_01030_),
    .Y(_04532_));
 OA211x2_ASAP7_75t_R _21945_ (.A1(net339),
    .A2(_04531_),
    .B(_04532_),
    .C(net308),
    .Y(_04533_));
 INVx1_ASAP7_75t_R _21946_ (.A(_01031_),
    .Y(_04534_));
 NAND2x1_ASAP7_75t_R _21947_ (.A(net339),
    .B(_01029_),
    .Y(_04535_));
 OA211x2_ASAP7_75t_R _21948_ (.A1(net339),
    .A2(_04534_),
    .B(_04535_),
    .C(net359),
    .Y(_04536_));
 OR3x1_ASAP7_75t_R _21949_ (.A(_13598_),
    .B(_04533_),
    .C(_04536_),
    .Y(_04537_));
 INVx1_ASAP7_75t_R _21950_ (.A(_01040_),
    .Y(_04538_));
 NAND2x1_ASAP7_75t_R _21951_ (.A(net339),
    .B(_01038_),
    .Y(_04539_));
 OA211x2_ASAP7_75t_R _21952_ (.A1(net339),
    .A2(_04538_),
    .B(_04539_),
    .C(net308),
    .Y(_04540_));
 INVx1_ASAP7_75t_R _21953_ (.A(_01039_),
    .Y(_04541_));
 NAND2x1_ASAP7_75t_R _21954_ (.A(net339),
    .B(_01037_),
    .Y(_04542_));
 OA211x2_ASAP7_75t_R _21955_ (.A1(net339),
    .A2(_04541_),
    .B(_04542_),
    .C(net359),
    .Y(_04543_));
 OR3x1_ASAP7_75t_R _21956_ (.A(net319),
    .B(_04540_),
    .C(_04543_),
    .Y(_04544_));
 AND3x1_ASAP7_75t_R _21957_ (.A(_01744_),
    .B(_04537_),
    .C(_04544_),
    .Y(_04545_));
 OR3x1_ASAP7_75t_R _21958_ (.A(net315),
    .B(_04530_),
    .C(_04545_),
    .Y(_04546_));
 OA21x2_ASAP7_75t_R _21959_ (.A1(_13174_),
    .A2(_04515_),
    .B(_04546_),
    .Y(_04547_));
 INVx1_ASAP7_75t_R _21960_ (.A(_04547_),
    .Y(_04548_));
 OA21x2_ASAP7_75t_R _21961_ (.A1(_00245_),
    .A2(_15267_),
    .B(_16207_),
    .Y(_04549_));
 AO21x2_ASAP7_75t_R _21962_ (.A1(_13583_),
    .A2(_04548_),
    .B(_04549_),
    .Y(_18223_));
 INVx1_ASAP7_75t_R _21963_ (.A(_18223_),
    .Y(_18221_));
 XNOR2x1_ASAP7_75t_R _21964_ (.B(_18223_),
    .Y(_04550_),
    .A(_13387_));
 NAND2x1_ASAP7_75t_R _21965_ (.A(net398),
    .B(_01033_),
    .Y(_04551_));
 OA211x2_ASAP7_75t_R _21966_ (.A1(net398),
    .A2(_04519_),
    .B(_04551_),
    .C(_13397_),
    .Y(_04552_));
 NAND2x1_ASAP7_75t_R _21967_ (.A(net398),
    .B(_01029_),
    .Y(_04553_));
 OA211x2_ASAP7_75t_R _21968_ (.A1(net398),
    .A2(_04534_),
    .B(_04553_),
    .C(net371),
    .Y(_04554_));
 OR3x1_ASAP7_75t_R _21969_ (.A(net306),
    .B(_04552_),
    .C(_04554_),
    .Y(_04555_));
 NAND2x1_ASAP7_75t_R _21970_ (.A(net398),
    .B(_01034_),
    .Y(_04556_));
 OA211x2_ASAP7_75t_R _21971_ (.A1(net398),
    .A2(_04516_),
    .B(_04556_),
    .C(_13397_),
    .Y(_04557_));
 NAND2x1_ASAP7_75t_R _21972_ (.A(net398),
    .B(_01030_),
    .Y(_04558_));
 OA211x2_ASAP7_75t_R _21973_ (.A1(net398),
    .A2(_04531_),
    .B(_04558_),
    .C(net371),
    .Y(_04559_));
 OR3x1_ASAP7_75t_R _21974_ (.A(_00290_),
    .B(_04557_),
    .C(_04559_),
    .Y(_04560_));
 AND3x1_ASAP7_75t_R _21975_ (.A(net367),
    .B(_04555_),
    .C(_04560_),
    .Y(_04561_));
 NAND2x1_ASAP7_75t_R _21976_ (.A(net398),
    .B(_01041_),
    .Y(_04562_));
 OA211x2_ASAP7_75t_R _21977_ (.A1(net398),
    .A2(_04526_),
    .B(_04562_),
    .C(_13397_),
    .Y(_04563_));
 NAND2x1_ASAP7_75t_R _21978_ (.A(net398),
    .B(_01037_),
    .Y(_04564_));
 OA211x2_ASAP7_75t_R _21979_ (.A1(net398),
    .A2(_04541_),
    .B(_04564_),
    .C(net371),
    .Y(_04565_));
 OR3x1_ASAP7_75t_R _21980_ (.A(net306),
    .B(_04563_),
    .C(_04565_),
    .Y(_04566_));
 NAND2x1_ASAP7_75t_R _21981_ (.A(net398),
    .B(_01042_),
    .Y(_04567_));
 OA211x2_ASAP7_75t_R _21982_ (.A1(net398),
    .A2(_04523_),
    .B(_04567_),
    .C(_13397_),
    .Y(_04568_));
 NAND2x1_ASAP7_75t_R _21983_ (.A(net398),
    .B(_01038_),
    .Y(_04569_));
 OA211x2_ASAP7_75t_R _21984_ (.A1(net398),
    .A2(_04538_),
    .B(_04569_),
    .C(net371),
    .Y(_04570_));
 OR3x1_ASAP7_75t_R _21985_ (.A(_00290_),
    .B(_04568_),
    .C(_04570_),
    .Y(_04571_));
 AND3x1_ASAP7_75t_R _21986_ (.A(_13484_),
    .B(_04566_),
    .C(_04571_),
    .Y(_04572_));
 OR2x2_ASAP7_75t_R _21987_ (.A(_04561_),
    .B(_04572_),
    .Y(_04573_));
 NAND2x1_ASAP7_75t_R _21988_ (.A(net399),
    .B(_01018_),
    .Y(_04574_));
 OA211x2_ASAP7_75t_R _21989_ (.A1(net399),
    .A2(_16492_),
    .B(_04574_),
    .C(net306),
    .Y(_04575_));
 NAND2x1_ASAP7_75t_R _21990_ (.A(net399),
    .B(_01017_),
    .Y(_04576_));
 OA211x2_ASAP7_75t_R _21991_ (.A1(net399),
    .A2(_16495_),
    .B(_04576_),
    .C(net410),
    .Y(_04577_));
 INVx1_ASAP7_75t_R _21992_ (.A(_01016_),
    .Y(_04578_));
 NAND2x1_ASAP7_75t_R _21993_ (.A(net399),
    .B(_01686_),
    .Y(_04579_));
 OA211x2_ASAP7_75t_R _21994_ (.A1(net399),
    .A2(_04578_),
    .B(_04579_),
    .C(net306),
    .Y(_04580_));
 NOR2x1_ASAP7_75t_R _21995_ (.A(_01015_),
    .B(_13471_),
    .Y(_04581_));
 OA33x2_ASAP7_75t_R _21996_ (.A1(_13814_),
    .A2(_04575_),
    .A3(_04577_),
    .B1(_04580_),
    .B2(_04581_),
    .B3(_13828_),
    .Y(_04582_));
 NAND2x1_ASAP7_75t_R _21997_ (.A(net399),
    .B(_01022_),
    .Y(_04583_));
 OA211x2_ASAP7_75t_R _21998_ (.A1(net399),
    .A2(_16484_),
    .B(_04583_),
    .C(net306),
    .Y(_04584_));
 NAND2x1_ASAP7_75t_R _21999_ (.A(net399),
    .B(_01021_),
    .Y(_04585_));
 OA211x2_ASAP7_75t_R _22000_ (.A1(net399),
    .A2(_16487_),
    .B(_04585_),
    .C(net410),
    .Y(_04586_));
 OR3x1_ASAP7_75t_R _22001_ (.A(_13397_),
    .B(_04584_),
    .C(_04586_),
    .Y(_04587_));
 NAND2x1_ASAP7_75t_R _22002_ (.A(net399),
    .B(_01026_),
    .Y(_04588_));
 OA211x2_ASAP7_75t_R _22003_ (.A1(net399),
    .A2(_04507_),
    .B(_04588_),
    .C(net306),
    .Y(_04589_));
 NAND2x1_ASAP7_75t_R _22004_ (.A(net399),
    .B(_01025_),
    .Y(_04590_));
 OA211x2_ASAP7_75t_R _22005_ (.A1(net399),
    .A2(_04510_),
    .B(_04590_),
    .C(net410),
    .Y(_04591_));
 OR3x1_ASAP7_75t_R _22006_ (.A(net371),
    .B(_04589_),
    .C(_04591_),
    .Y(_04592_));
 AO21x1_ASAP7_75t_R _22007_ (.A1(_04587_),
    .A2(_04592_),
    .B(net367),
    .Y(_04593_));
 AO21x1_ASAP7_75t_R _22008_ (.A1(_04582_),
    .A2(_04593_),
    .B(_13392_),
    .Y(_04594_));
 OA21x2_ASAP7_75t_R _22009_ (.A1(net364),
    .A2(_04573_),
    .B(_04594_),
    .Y(_04595_));
 BUFx2_ASAP7_75t_R output239 (.A(net239),
    .Y(instr_addr_o[2]));
 AOI22x1_ASAP7_75t_R _22011_ (.A1(_13530_),
    .A2(_01045_),
    .B1(_02210_),
    .B2(_13533_),
    .Y(_04597_));
 OA211x2_ASAP7_75t_R _22012_ (.A1(_00284_),
    .A2(_04595_),
    .B(_04597_),
    .C(_13763_),
    .Y(_04598_));
 AO21x1_ASAP7_75t_R _22013_ (.A1(_13528_),
    .A2(_04547_),
    .B(_04598_),
    .Y(_04599_));
 AND2x2_ASAP7_75t_R _22014_ (.A(_13576_),
    .B(_04599_),
    .Y(_04600_));
 AOI21x1_ASAP7_75t_R _22015_ (.A1(net295),
    .A2(_04550_),
    .B(_04600_),
    .Y(_17577_));
 INVx1_ASAP7_75t_R _22016_ (.A(_17577_),
    .Y(_16536_));
 INVx2_ASAP7_75t_R _22017_ (.A(_00218_),
    .Y(\cs_registers_i.pc_id_i[23] ));
 OA211x2_ASAP7_75t_R _22018_ (.A1(net364),
    .A2(_04573_),
    .B(_04594_),
    .C(_13563_),
    .Y(_04601_));
 OAI22x1_ASAP7_75t_R _22019_ (.A1(_01618_),
    .A2(_13223_),
    .B1(_13880_),
    .B2(_00218_),
    .Y(_04602_));
 OR2x4_ASAP7_75t_R _22020_ (.A(_04601_),
    .B(_04602_),
    .Y(_04603_));
 BUFx2_ASAP7_75t_R output238 (.A(net238),
    .Y(instr_addr_o[29]));
 INVx2_ASAP7_75t_R _22022_ (.A(_04603_),
    .Y(_18222_));
 OA21x2_ASAP7_75t_R _22023_ (.A1(_01045_),
    .A2(_13574_),
    .B(_13576_),
    .Y(_04604_));
 AOI21x1_ASAP7_75t_R _22024_ (.A1(net295),
    .A2(_18222_),
    .B(_04604_),
    .Y(_17576_));
 INVx1_ASAP7_75t_R _22025_ (.A(_17576_),
    .Y(_16535_));
 OR4x2_ASAP7_75t_R _22026_ (.A(_00947_),
    .B(_00915_),
    .C(_01012_),
    .D(_00980_),
    .Y(_04605_));
 OA21x2_ASAP7_75t_R _22027_ (.A1(_00947_),
    .A2(_00948_),
    .B(_02277_),
    .Y(_04606_));
 OA21x2_ASAP7_75t_R _22028_ (.A1(_00980_),
    .A2(_04606_),
    .B(_01013_),
    .Y(_04607_));
 OA21x2_ASAP7_75t_R _22029_ (.A1(_01012_),
    .A2(_04607_),
    .B(_02278_),
    .Y(_04608_));
 OA21x2_ASAP7_75t_R _22030_ (.A1(_16529_),
    .A2(_04605_),
    .B(_04608_),
    .Y(_16534_));
 AND2x2_ASAP7_75t_R _22031_ (.A(net332),
    .B(_01685_),
    .Y(_04609_));
 AO21x1_ASAP7_75t_R _22032_ (.A1(net313),
    .A2(_01048_),
    .B(_04609_),
    .Y(_04610_));
 OAI22x1_ASAP7_75t_R _22033_ (.A1(_01047_),
    .A2(_13586_),
    .B1(_04610_),
    .B2(net357),
    .Y(_04611_));
 INVx1_ASAP7_75t_R _22034_ (.A(_01056_),
    .Y(_04612_));
 NAND2x1_ASAP7_75t_R _22035_ (.A(net331),
    .B(_01054_),
    .Y(_04613_));
 OA211x2_ASAP7_75t_R _22036_ (.A1(net331),
    .A2(_04612_),
    .B(_04613_),
    .C(net308),
    .Y(_04614_));
 INVx1_ASAP7_75t_R _22037_ (.A(_01055_),
    .Y(_04615_));
 NAND2x1_ASAP7_75t_R _22038_ (.A(net331),
    .B(_01053_),
    .Y(_04616_));
 OA211x2_ASAP7_75t_R _22039_ (.A1(net331),
    .A2(_04615_),
    .B(_04616_),
    .C(net357),
    .Y(_04617_));
 OR3x1_ASAP7_75t_R _22040_ (.A(net318),
    .B(_04614_),
    .C(_04617_),
    .Y(_04618_));
 OA211x2_ASAP7_75t_R _22041_ (.A1(_13598_),
    .A2(_04611_),
    .B(_04618_),
    .C(net325),
    .Y(_04619_));
 INVx1_ASAP7_75t_R _22042_ (.A(_01052_),
    .Y(_04620_));
 NAND2x1_ASAP7_75t_R _22043_ (.A(net332),
    .B(_01050_),
    .Y(_04621_));
 OA211x2_ASAP7_75t_R _22044_ (.A1(net332),
    .A2(_04620_),
    .B(_04621_),
    .C(net308),
    .Y(_04622_));
 INVx1_ASAP7_75t_R _22045_ (.A(_01051_),
    .Y(_04623_));
 NAND2x1_ASAP7_75t_R _22046_ (.A(net332),
    .B(_01049_),
    .Y(_04624_));
 OA211x2_ASAP7_75t_R _22047_ (.A1(net332),
    .A2(_04623_),
    .B(_04624_),
    .C(net357),
    .Y(_04625_));
 OR3x1_ASAP7_75t_R _22048_ (.A(_13598_),
    .B(_04622_),
    .C(_04625_),
    .Y(_04626_));
 INVx1_ASAP7_75t_R _22049_ (.A(_01060_),
    .Y(_04627_));
 NAND2x1_ASAP7_75t_R _22050_ (.A(net332),
    .B(_01058_),
    .Y(_04628_));
 OA211x2_ASAP7_75t_R _22051_ (.A1(net332),
    .A2(_04627_),
    .B(_04628_),
    .C(net308),
    .Y(_04629_));
 INVx1_ASAP7_75t_R _22052_ (.A(_01059_),
    .Y(_04630_));
 NAND2x1_ASAP7_75t_R _22053_ (.A(net335),
    .B(_01057_),
    .Y(_04631_));
 OA211x2_ASAP7_75t_R _22054_ (.A1(net335),
    .A2(_04630_),
    .B(_04631_),
    .C(net357),
    .Y(_04632_));
 OR3x1_ASAP7_75t_R _22055_ (.A(net318),
    .B(_04629_),
    .C(_04632_),
    .Y(_04633_));
 AND3x1_ASAP7_75t_R _22056_ (.A(_13132_),
    .B(_04626_),
    .C(_04633_),
    .Y(_04634_));
 OR3x1_ASAP7_75t_R _22057_ (.A(_13174_),
    .B(_04619_),
    .C(_04634_),
    .Y(_04635_));
 INVx1_ASAP7_75t_R _22058_ (.A(_01061_),
    .Y(_04636_));
 NOR2x1_ASAP7_75t_R _22059_ (.A(net331),
    .B(_01063_),
    .Y(_04637_));
 AO21x1_ASAP7_75t_R _22060_ (.A1(net331),
    .A2(_04636_),
    .B(_04637_),
    .Y(_04638_));
 INVx1_ASAP7_75t_R _22061_ (.A(_01064_),
    .Y(_04639_));
 NAND2x1_ASAP7_75t_R _22062_ (.A(net331),
    .B(_01062_),
    .Y(_04640_));
 OA211x2_ASAP7_75t_R _22063_ (.A1(net331),
    .A2(_04639_),
    .B(_04640_),
    .C(net308),
    .Y(_04641_));
 AO21x1_ASAP7_75t_R _22064_ (.A1(net357),
    .A2(_04638_),
    .B(_04641_),
    .Y(_04642_));
 INVx1_ASAP7_75t_R _22065_ (.A(_01068_),
    .Y(_04643_));
 NAND2x1_ASAP7_75t_R _22066_ (.A(net331),
    .B(_01066_),
    .Y(_04644_));
 OA211x2_ASAP7_75t_R _22067_ (.A1(net331),
    .A2(_04643_),
    .B(_04644_),
    .C(net308),
    .Y(_04645_));
 INVx1_ASAP7_75t_R _22068_ (.A(_01067_),
    .Y(_04646_));
 NAND2x1_ASAP7_75t_R _22069_ (.A(net331),
    .B(_01065_),
    .Y(_04647_));
 OA211x2_ASAP7_75t_R _22070_ (.A1(net331),
    .A2(_04646_),
    .B(_04647_),
    .C(net357),
    .Y(_04648_));
 OR3x1_ASAP7_75t_R _22071_ (.A(net325),
    .B(_04645_),
    .C(_04648_),
    .Y(_04649_));
 OA211x2_ASAP7_75t_R _22072_ (.A1(_13132_),
    .A2(_04642_),
    .B(_04649_),
    .C(net318),
    .Y(_04650_));
 INVx1_ASAP7_75t_R _22073_ (.A(_01076_),
    .Y(_04651_));
 NAND2x1_ASAP7_75t_R _22074_ (.A(net331),
    .B(_01074_),
    .Y(_04652_));
 OA211x2_ASAP7_75t_R _22075_ (.A1(net331),
    .A2(_04651_),
    .B(_04652_),
    .C(_13145_),
    .Y(_04653_));
 INVx1_ASAP7_75t_R _22076_ (.A(_01075_),
    .Y(_04654_));
 NAND2x1_ASAP7_75t_R _22077_ (.A(net331),
    .B(_01073_),
    .Y(_04655_));
 OA211x2_ASAP7_75t_R _22078_ (.A1(net331),
    .A2(_04654_),
    .B(_04655_),
    .C(net356),
    .Y(_04656_));
 OR3x1_ASAP7_75t_R _22079_ (.A(net325),
    .B(_04653_),
    .C(_04656_),
    .Y(_04657_));
 INVx1_ASAP7_75t_R _22080_ (.A(_01072_),
    .Y(_04658_));
 NAND2x1_ASAP7_75t_R _22081_ (.A(net331),
    .B(_01070_),
    .Y(_04659_));
 OA211x2_ASAP7_75t_R _22082_ (.A1(net331),
    .A2(_04658_),
    .B(_04659_),
    .C(_13145_),
    .Y(_04660_));
 INVx1_ASAP7_75t_R _22083_ (.A(_01071_),
    .Y(_04661_));
 NAND2x1_ASAP7_75t_R _22084_ (.A(net331),
    .B(_01069_),
    .Y(_04662_));
 OA211x2_ASAP7_75t_R _22085_ (.A1(net331),
    .A2(_04661_),
    .B(_04662_),
    .C(net356),
    .Y(_04663_));
 OR3x1_ASAP7_75t_R _22086_ (.A(_13132_),
    .B(_04660_),
    .C(_04663_),
    .Y(_04664_));
 AND3x1_ASAP7_75t_R _22087_ (.A(_13598_),
    .B(_04657_),
    .C(_04664_),
    .Y(_04665_));
 OR3x2_ASAP7_75t_R _22088_ (.A(net315),
    .B(_04650_),
    .C(_04665_),
    .Y(_04666_));
 AND2x6_ASAP7_75t_R _22089_ (.A(_04635_),
    .B(_04666_),
    .Y(_04667_));
 INVx4_ASAP7_75t_R _22090_ (.A(_04667_),
    .Y(_04668_));
 OA21x2_ASAP7_75t_R _22091_ (.A1(net316),
    .A2(_15267_),
    .B(_16207_),
    .Y(_04669_));
 AO21x1_ASAP7_75t_R _22092_ (.A1(_13583_),
    .A2(_04668_),
    .B(_04669_),
    .Y(_18225_));
 INVx1_ASAP7_75t_R _22093_ (.A(_18225_),
    .Y(_18227_));
 NAND2x1_ASAP7_75t_R _22094_ (.A(net391),
    .B(_01049_),
    .Y(_04670_));
 OA211x2_ASAP7_75t_R _22095_ (.A1(net391),
    .A2(_04623_),
    .B(_04670_),
    .C(net409),
    .Y(_04671_));
 NAND2x1_ASAP7_75t_R _22096_ (.A(net391),
    .B(_01050_),
    .Y(_04672_));
 OA211x2_ASAP7_75t_R _22097_ (.A1(net391),
    .A2(_04620_),
    .B(_04672_),
    .C(net306),
    .Y(_04673_));
 INVx1_ASAP7_75t_R _22098_ (.A(_01048_),
    .Y(_04674_));
 NAND2x1_ASAP7_75t_R _22099_ (.A(net391),
    .B(_01685_),
    .Y(_04675_));
 OA211x2_ASAP7_75t_R _22100_ (.A1(net391),
    .A2(_04674_),
    .B(_04675_),
    .C(net306),
    .Y(_04676_));
 NOR2x1_ASAP7_75t_R _22101_ (.A(_01047_),
    .B(_13471_),
    .Y(_04677_));
 OA33x2_ASAP7_75t_R _22102_ (.A1(_13814_),
    .A2(_04671_),
    .A3(_04673_),
    .B1(_04676_),
    .B2(_04677_),
    .B3(_13828_),
    .Y(_04678_));
 NAND2x1_ASAP7_75t_R _22103_ (.A(net390),
    .B(_01065_),
    .Y(_04679_));
 OA211x2_ASAP7_75t_R _22104_ (.A1(net390),
    .A2(_04646_),
    .B(_04679_),
    .C(_13397_),
    .Y(_04680_));
 NAND2x1_ASAP7_75t_R _22105_ (.A(net302),
    .B(_01063_),
    .Y(_04681_));
 OA211x2_ASAP7_75t_R _22106_ (.A1(net302),
    .A2(_04636_),
    .B(_04681_),
    .C(net370),
    .Y(_04682_));
 OR3x1_ASAP7_75t_R _22107_ (.A(net306),
    .B(_04680_),
    .C(_04682_),
    .Y(_04683_));
 NAND2x1_ASAP7_75t_R _22108_ (.A(net390),
    .B(_01066_),
    .Y(_04684_));
 OA211x2_ASAP7_75t_R _22109_ (.A1(net390),
    .A2(_04643_),
    .B(_04684_),
    .C(_13397_),
    .Y(_04685_));
 NAND2x1_ASAP7_75t_R _22110_ (.A(net390),
    .B(_01062_),
    .Y(_04686_));
 OA211x2_ASAP7_75t_R _22111_ (.A1(net390),
    .A2(_04639_),
    .B(_04686_),
    .C(net370),
    .Y(_04687_));
 OR3x1_ASAP7_75t_R _22112_ (.A(net408),
    .B(_04685_),
    .C(_04687_),
    .Y(_04688_));
 AND2x2_ASAP7_75t_R _22113_ (.A(net366),
    .B(_13392_),
    .Y(_04689_));
 INVx2_ASAP7_75t_R _22114_ (.A(_04689_),
    .Y(_04690_));
 AO21x1_ASAP7_75t_R _22115_ (.A1(_04683_),
    .A2(_04688_),
    .B(_04690_),
    .Y(_04691_));
 NAND2x1_ASAP7_75t_R _22116_ (.A(net391),
    .B(_01054_),
    .Y(_04692_));
 OA211x2_ASAP7_75t_R _22117_ (.A1(net390),
    .A2(_04612_),
    .B(_04692_),
    .C(net306),
    .Y(_04693_));
 NAND2x1_ASAP7_75t_R _22118_ (.A(net390),
    .B(_01053_),
    .Y(_04694_));
 OA211x2_ASAP7_75t_R _22119_ (.A1(net390),
    .A2(_04615_),
    .B(_04694_),
    .C(net408),
    .Y(_04695_));
 OR3x1_ASAP7_75t_R _22120_ (.A(_13397_),
    .B(_04693_),
    .C(_04695_),
    .Y(_04696_));
 NAND2x1_ASAP7_75t_R _22121_ (.A(net391),
    .B(_01058_),
    .Y(_04697_));
 OA211x2_ASAP7_75t_R _22122_ (.A1(net391),
    .A2(_04627_),
    .B(_04697_),
    .C(net306),
    .Y(_04698_));
 NAND2x1_ASAP7_75t_R _22123_ (.A(net391),
    .B(_01057_),
    .Y(_04699_));
 OA211x2_ASAP7_75t_R _22124_ (.A1(net391),
    .A2(_04630_),
    .B(_04699_),
    .C(net409),
    .Y(_04700_));
 OR3x1_ASAP7_75t_R _22125_ (.A(net372),
    .B(_04698_),
    .C(_04700_),
    .Y(_04701_));
 AND3x1_ASAP7_75t_R _22126_ (.A(net362),
    .B(_04696_),
    .C(_04701_),
    .Y(_04702_));
 NAND2x1_ASAP7_75t_R _22127_ (.A(net390),
    .B(_01073_),
    .Y(_04703_));
 OA211x2_ASAP7_75t_R _22128_ (.A1(net390),
    .A2(_04654_),
    .B(_04703_),
    .C(_13397_),
    .Y(_04704_));
 NAND2x1_ASAP7_75t_R _22129_ (.A(net390),
    .B(_01069_),
    .Y(_04705_));
 OA211x2_ASAP7_75t_R _22130_ (.A1(net390),
    .A2(_04661_),
    .B(_04705_),
    .C(net370),
    .Y(_04706_));
 OR3x1_ASAP7_75t_R _22131_ (.A(_13424_),
    .B(_04704_),
    .C(_04706_),
    .Y(_04707_));
 NAND2x1_ASAP7_75t_R _22132_ (.A(net390),
    .B(_01074_),
    .Y(_04708_));
 OA211x2_ASAP7_75t_R _22133_ (.A1(net390),
    .A2(_04651_),
    .B(_04708_),
    .C(_13397_),
    .Y(_04709_));
 NAND2x1_ASAP7_75t_R _22134_ (.A(net390),
    .B(_01070_),
    .Y(_04710_));
 OA211x2_ASAP7_75t_R _22135_ (.A1(net390),
    .A2(_04658_),
    .B(_04710_),
    .C(net370),
    .Y(_04711_));
 OR3x1_ASAP7_75t_R _22136_ (.A(net408),
    .B(_04709_),
    .C(_04711_),
    .Y(_04712_));
 AND3x1_ASAP7_75t_R _22137_ (.A(_13392_),
    .B(_04707_),
    .C(_04712_),
    .Y(_04713_));
 OR3x1_ASAP7_75t_R _22138_ (.A(net365),
    .B(_04702_),
    .C(_04713_),
    .Y(_04714_));
 OA211x2_ASAP7_75t_R _22139_ (.A1(_13392_),
    .A2(_04678_),
    .B(_04691_),
    .C(_04714_),
    .Y(_04715_));
 BUFx2_ASAP7_75t_R output237 (.A(net237),
    .Y(instr_addr_o[28]));
 OAI22x1_ASAP7_75t_R _22141_ (.A1(_01617_),
    .A2(_13223_),
    .B1(_13880_),
    .B2(_00220_),
    .Y(_04717_));
 AO21x2_ASAP7_75t_R _22142_ (.A1(_13563_),
    .A2(_04715_),
    .B(_04717_),
    .Y(_04718_));
 BUFx2_ASAP7_75t_R output236 (.A(net236),
    .Y(instr_addr_o[27]));
 INVx2_ASAP7_75t_R _22144_ (.A(_04718_),
    .Y(_18226_));
 XOR2x2_ASAP7_75t_R _22145_ (.A(_01078_),
    .B(_02230_),
    .Y(_04719_));
 INVx4_ASAP7_75t_R _22146_ (.A(_04719_),
    .Y(net165));
 INVx1_ASAP7_75t_R _22147_ (.A(_01089_),
    .Y(_04720_));
 NAND2x1_ASAP7_75t_R _22148_ (.A(net345),
    .B(_01087_),
    .Y(_04721_));
 OA211x2_ASAP7_75t_R _22149_ (.A1(net345),
    .A2(_04720_),
    .B(_04721_),
    .C(net311),
    .Y(_04722_));
 INVx1_ASAP7_75t_R _22150_ (.A(_01088_),
    .Y(_04723_));
 NAND2x1_ASAP7_75t_R _22151_ (.A(net345),
    .B(_01086_),
    .Y(_04724_));
 OA211x2_ASAP7_75t_R _22152_ (.A1(net345),
    .A2(_04723_),
    .B(_04724_),
    .C(net355),
    .Y(_04725_));
 OR3x1_ASAP7_75t_R _22153_ (.A(net318),
    .B(_04722_),
    .C(_04725_),
    .Y(_04726_));
 INVx1_ASAP7_75t_R _22154_ (.A(_01080_),
    .Y(_04727_));
 INVx1_ASAP7_75t_R _22155_ (.A(_01081_),
    .Y(_04728_));
 NAND2x1_ASAP7_75t_R _22156_ (.A(net342),
    .B(_01684_),
    .Y(_04729_));
 OA21x2_ASAP7_75t_R _22157_ (.A1(net342),
    .A2(_04728_),
    .B(_04729_),
    .Y(_04730_));
 AO221x1_ASAP7_75t_R _22158_ (.A1(_04727_),
    .A2(_13190_),
    .B1(_04730_),
    .B2(net311),
    .C(_13598_),
    .Y(_04731_));
 AO21x1_ASAP7_75t_R _22159_ (.A1(_04726_),
    .A2(_04731_),
    .B(_13132_),
    .Y(_04732_));
 INVx1_ASAP7_75t_R _22160_ (.A(_01085_),
    .Y(_04733_));
 NAND2x1_ASAP7_75t_R _22161_ (.A(net345),
    .B(_01083_),
    .Y(_04734_));
 OA211x2_ASAP7_75t_R _22162_ (.A1(net345),
    .A2(_04733_),
    .B(_04734_),
    .C(net311),
    .Y(_04735_));
 INVx1_ASAP7_75t_R _22163_ (.A(_01084_),
    .Y(_04736_));
 NAND2x1_ASAP7_75t_R _22164_ (.A(net345),
    .B(_01082_),
    .Y(_04737_));
 OA211x2_ASAP7_75t_R _22165_ (.A1(net345),
    .A2(_04736_),
    .B(_04737_),
    .C(net355),
    .Y(_04738_));
 OR3x1_ASAP7_75t_R _22166_ (.A(_13598_),
    .B(_04735_),
    .C(_04738_),
    .Y(_04739_));
 INVx1_ASAP7_75t_R _22167_ (.A(_01093_),
    .Y(_04740_));
 NAND2x1_ASAP7_75t_R _22168_ (.A(net342),
    .B(_01091_),
    .Y(_04741_));
 OA211x2_ASAP7_75t_R _22169_ (.A1(net342),
    .A2(_04740_),
    .B(_04741_),
    .C(net311),
    .Y(_04742_));
 INVx1_ASAP7_75t_R _22170_ (.A(_01092_),
    .Y(_04743_));
 NAND2x1_ASAP7_75t_R _22171_ (.A(net342),
    .B(_01090_),
    .Y(_04744_));
 OA211x2_ASAP7_75t_R _22172_ (.A1(net342),
    .A2(_04743_),
    .B(_04744_),
    .C(net355),
    .Y(_04745_));
 OR3x1_ASAP7_75t_R _22173_ (.A(net318),
    .B(_04742_),
    .C(_04745_),
    .Y(_04746_));
 AO21x1_ASAP7_75t_R _22174_ (.A1(_04739_),
    .A2(_04746_),
    .B(net324),
    .Y(_04747_));
 AO21x2_ASAP7_75t_R _22175_ (.A1(_04732_),
    .A2(_04747_),
    .B(_13174_),
    .Y(_04748_));
 INVx1_ASAP7_75t_R _22176_ (.A(_01109_),
    .Y(_04749_));
 NAND2x1_ASAP7_75t_R _22177_ (.A(net342),
    .B(_01107_),
    .Y(_04750_));
 OA211x2_ASAP7_75t_R _22178_ (.A1(net342),
    .A2(_04749_),
    .B(_04750_),
    .C(net311),
    .Y(_04751_));
 INVx1_ASAP7_75t_R _22179_ (.A(_01108_),
    .Y(_04752_));
 NAND2x1_ASAP7_75t_R _22180_ (.A(net342),
    .B(_01106_),
    .Y(_04753_));
 OA211x2_ASAP7_75t_R _22181_ (.A1(net342),
    .A2(_04752_),
    .B(_04753_),
    .C(net355),
    .Y(_04754_));
 OR3x1_ASAP7_75t_R _22182_ (.A(net324),
    .B(_04751_),
    .C(_04754_),
    .Y(_04755_));
 INVx1_ASAP7_75t_R _22183_ (.A(_01105_),
    .Y(_04756_));
 NAND2x1_ASAP7_75t_R _22184_ (.A(net342),
    .B(_01103_),
    .Y(_04757_));
 OA211x2_ASAP7_75t_R _22185_ (.A1(net342),
    .A2(_04756_),
    .B(_04757_),
    .C(net311),
    .Y(_04758_));
 INVx1_ASAP7_75t_R _22186_ (.A(_01104_),
    .Y(_04759_));
 NAND2x1_ASAP7_75t_R _22187_ (.A(net342),
    .B(_01102_),
    .Y(_04760_));
 OA211x2_ASAP7_75t_R _22188_ (.A1(net342),
    .A2(_04759_),
    .B(_04760_),
    .C(net355),
    .Y(_04761_));
 OR3x1_ASAP7_75t_R _22189_ (.A(_13132_),
    .B(_04758_),
    .C(_04761_),
    .Y(_04762_));
 AND3x1_ASAP7_75t_R _22190_ (.A(_13598_),
    .B(_04755_),
    .C(_04762_),
    .Y(_04763_));
 INVx1_ASAP7_75t_R _22191_ (.A(_01097_),
    .Y(_04764_));
 NAND2x1_ASAP7_75t_R _22192_ (.A(net342),
    .B(_01095_),
    .Y(_04765_));
 OA211x2_ASAP7_75t_R _22193_ (.A1(net342),
    .A2(_04764_),
    .B(_04765_),
    .C(net311),
    .Y(_04766_));
 INVx1_ASAP7_75t_R _22194_ (.A(_01096_),
    .Y(_04767_));
 NAND2x1_ASAP7_75t_R _22195_ (.A(net342),
    .B(_01094_),
    .Y(_04768_));
 OA211x2_ASAP7_75t_R _22196_ (.A1(net342),
    .A2(_04767_),
    .B(_04768_),
    .C(net355),
    .Y(_04769_));
 OR3x1_ASAP7_75t_R _22197_ (.A(_13132_),
    .B(_04766_),
    .C(_04769_),
    .Y(_04770_));
 INVx1_ASAP7_75t_R _22198_ (.A(_01101_),
    .Y(_04771_));
 NAND2x1_ASAP7_75t_R _22199_ (.A(net342),
    .B(_01099_),
    .Y(_04772_));
 OA211x2_ASAP7_75t_R _22200_ (.A1(net342),
    .A2(_04771_),
    .B(_04772_),
    .C(net311),
    .Y(_04773_));
 INVx1_ASAP7_75t_R _22201_ (.A(_01100_),
    .Y(_04774_));
 NAND2x1_ASAP7_75t_R _22202_ (.A(net342),
    .B(_01098_),
    .Y(_04775_));
 OA211x2_ASAP7_75t_R _22203_ (.A1(net342),
    .A2(_04774_),
    .B(_04775_),
    .C(net355),
    .Y(_04776_));
 OR3x1_ASAP7_75t_R _22204_ (.A(net324),
    .B(_04773_),
    .C(_04776_),
    .Y(_04777_));
 AND3x1_ASAP7_75t_R _22205_ (.A(net318),
    .B(_04770_),
    .C(_04777_),
    .Y(_04778_));
 OR3x4_ASAP7_75t_R _22206_ (.A(net315),
    .B(_04763_),
    .C(_04778_),
    .Y(_04779_));
 NAND2x2_ASAP7_75t_R _22207_ (.A(_04748_),
    .B(_04779_),
    .Y(_04780_));
 OA21x2_ASAP7_75t_R _22208_ (.A1(_01743_),
    .A2(_15267_),
    .B(_16207_),
    .Y(_04781_));
 AO21x2_ASAP7_75t_R _22209_ (.A1(_13583_),
    .A2(_04780_),
    .B(_04781_),
    .Y(_04782_));
 BUFx2_ASAP7_75t_R output235 (.A(net235),
    .Y(instr_addr_o[26]));
 INVx1_ASAP7_75t_R _22211_ (.A(_04782_),
    .Y(_18232_));
 INVx2_ASAP7_75t_R _22212_ (.A(_00221_),
    .Y(\cs_registers_i.pc_id_i[25] ));
 NOR2x1_ASAP7_75t_R _22213_ (.A(_01616_),
    .B(_13223_),
    .Y(_04783_));
 AOI21x1_ASAP7_75t_R _22214_ (.A1(_00221_),
    .A2(_13553_),
    .B(_13561_),
    .Y(_04784_));
 NAND2x1_ASAP7_75t_R _22215_ (.A(net387),
    .B(_01099_),
    .Y(_04785_));
 OA211x2_ASAP7_75t_R _22216_ (.A1(net387),
    .A2(_04771_),
    .B(_04785_),
    .C(net307),
    .Y(_04786_));
 NAND2x1_ASAP7_75t_R _22217_ (.A(net388),
    .B(_01098_),
    .Y(_04787_));
 OA211x2_ASAP7_75t_R _22218_ (.A1(net388),
    .A2(_04774_),
    .B(_04787_),
    .C(net407),
    .Y(_04788_));
 OR3x1_ASAP7_75t_R _22219_ (.A(_13814_),
    .B(_04786_),
    .C(_04788_),
    .Y(_04789_));
 NAND2x1_ASAP7_75t_R _22220_ (.A(net387),
    .B(_01095_),
    .Y(_04790_));
 OA211x2_ASAP7_75t_R _22221_ (.A1(net387),
    .A2(_04764_),
    .B(_04790_),
    .C(net307),
    .Y(_04791_));
 NAND2x1_ASAP7_75t_R _22222_ (.A(net387),
    .B(_01094_),
    .Y(_04792_));
 OA211x2_ASAP7_75t_R _22223_ (.A1(net387),
    .A2(_04767_),
    .B(_04792_),
    .C(net407),
    .Y(_04793_));
 OR3x1_ASAP7_75t_R _22224_ (.A(net301),
    .B(_04791_),
    .C(_04793_),
    .Y(_04794_));
 AND3x1_ASAP7_75t_R _22225_ (.A(_13392_),
    .B(_04789_),
    .C(_04794_),
    .Y(_04795_));
 NAND2x1_ASAP7_75t_R _22226_ (.A(net388),
    .B(_01103_),
    .Y(_04796_));
 OA211x2_ASAP7_75t_R _22227_ (.A1(net388),
    .A2(_04756_),
    .B(_04796_),
    .C(_13424_),
    .Y(_04797_));
 NAND2x1_ASAP7_75t_R _22228_ (.A(net388),
    .B(_01102_),
    .Y(_04798_));
 OA211x2_ASAP7_75t_R _22229_ (.A1(net388),
    .A2(_04759_),
    .B(_04798_),
    .C(net407),
    .Y(_04799_));
 OR3x1_ASAP7_75t_R _22230_ (.A(_13397_),
    .B(_04797_),
    .C(_04799_),
    .Y(_04800_));
 NAND2x1_ASAP7_75t_R _22231_ (.A(net387),
    .B(_01107_),
    .Y(_04801_));
 OA211x2_ASAP7_75t_R _22232_ (.A1(net387),
    .A2(_04749_),
    .B(_04801_),
    .C(_13424_),
    .Y(_04802_));
 NAND2x1_ASAP7_75t_R _22233_ (.A(net387),
    .B(_01106_),
    .Y(_04803_));
 OA211x2_ASAP7_75t_R _22234_ (.A1(net387),
    .A2(_04752_),
    .B(_04803_),
    .C(net407),
    .Y(_04804_));
 OR3x1_ASAP7_75t_R _22235_ (.A(net370),
    .B(_04802_),
    .C(_04804_),
    .Y(_04805_));
 AND2x2_ASAP7_75t_R _22236_ (.A(_04800_),
    .B(_04805_),
    .Y(_04806_));
 NAND2x1_ASAP7_75t_R _22237_ (.A(net388),
    .B(_01083_),
    .Y(_04807_));
 OA211x2_ASAP7_75t_R _22238_ (.A1(net388),
    .A2(_04733_),
    .B(_04807_),
    .C(net307),
    .Y(_04808_));
 NAND2x1_ASAP7_75t_R _22239_ (.A(net388),
    .B(_01082_),
    .Y(_04809_));
 OA211x2_ASAP7_75t_R _22240_ (.A1(net388),
    .A2(_04736_),
    .B(_04809_),
    .C(net407),
    .Y(_04810_));
 OR3x1_ASAP7_75t_R _22241_ (.A(_13814_),
    .B(_04808_),
    .C(_04810_),
    .Y(_04811_));
 NAND2x1_ASAP7_75t_R _22242_ (.A(net387),
    .B(_01684_),
    .Y(_04812_));
 OA211x2_ASAP7_75t_R _22243_ (.A1(net387),
    .A2(_04728_),
    .B(_04812_),
    .C(net307),
    .Y(_04813_));
 AND3x1_ASAP7_75t_R _22244_ (.A(net407),
    .B(net303),
    .C(_04727_),
    .Y(_04814_));
 OA31x2_ASAP7_75t_R _22245_ (.A1(net301),
    .A2(_04813_),
    .A3(_04814_),
    .B1(net363),
    .Y(_04815_));
 AO32x1_ASAP7_75t_R _22246_ (.A1(_13392_),
    .A2(_04789_),
    .A3(_04794_),
    .B1(_04811_),
    .B2(_04815_),
    .Y(_04816_));
 NAND2x1_ASAP7_75t_R _22247_ (.A(net387),
    .B(_01091_),
    .Y(_04817_));
 OA211x2_ASAP7_75t_R _22248_ (.A1(net387),
    .A2(_04740_),
    .B(_04817_),
    .C(net307),
    .Y(_04818_));
 NAND2x1_ASAP7_75t_R _22249_ (.A(net387),
    .B(_01090_),
    .Y(_04819_));
 OA211x2_ASAP7_75t_R _22250_ (.A1(net387),
    .A2(_04743_),
    .B(_04819_),
    .C(net407),
    .Y(_04820_));
 OR3x1_ASAP7_75t_R _22251_ (.A(net369),
    .B(_04818_),
    .C(_04820_),
    .Y(_04821_));
 NAND2x1_ASAP7_75t_R _22252_ (.A(net388),
    .B(_01087_),
    .Y(_04822_));
 OA211x2_ASAP7_75t_R _22253_ (.A1(net388),
    .A2(_04720_),
    .B(_04822_),
    .C(net307),
    .Y(_04823_));
 NAND2x1_ASAP7_75t_R _22254_ (.A(net388),
    .B(_01086_),
    .Y(_04824_));
 OA211x2_ASAP7_75t_R _22255_ (.A1(net388),
    .A2(_04723_),
    .B(_04824_),
    .C(net407),
    .Y(_04825_));
 OR3x1_ASAP7_75t_R _22256_ (.A(_13397_),
    .B(_04823_),
    .C(_04825_),
    .Y(_04826_));
 AND4x1_ASAP7_75t_R _22257_ (.A(_04811_),
    .B(_04815_),
    .C(_04821_),
    .D(_04826_),
    .Y(_04827_));
 AO221x2_ASAP7_75t_R _22258_ (.A1(_04795_),
    .A2(_04806_),
    .B1(_04816_),
    .B2(net366),
    .C(_04827_),
    .Y(_04828_));
 OA22x2_ASAP7_75t_R _22259_ (.A1(_04783_),
    .A2(_04784_),
    .B1(_04828_),
    .B2(_13782_),
    .Y(_04829_));
 BUFx2_ASAP7_75t_R output234 (.A(net234),
    .Y(instr_addr_o[25]));
 INVx2_ASAP7_75t_R _22261_ (.A(_04829_),
    .Y(_18231_));
 AND2x2_ASAP7_75t_R _22262_ (.A(net332),
    .B(_01683_),
    .Y(_04830_));
 AO21x1_ASAP7_75t_R _22263_ (.A1(net313),
    .A2(_01113_),
    .B(_04830_),
    .Y(_04831_));
 OAI22x1_ASAP7_75t_R _22264_ (.A1(_01112_),
    .A2(_13586_),
    .B1(_04831_),
    .B2(net356),
    .Y(_04832_));
 INVx1_ASAP7_75t_R _22265_ (.A(_01121_),
    .Y(_04833_));
 NAND2x1_ASAP7_75t_R _22266_ (.A(net332),
    .B(_01119_),
    .Y(_04834_));
 OA211x2_ASAP7_75t_R _22267_ (.A1(net332),
    .A2(_04833_),
    .B(_04834_),
    .C(net308),
    .Y(_04835_));
 INVx1_ASAP7_75t_R _22268_ (.A(_01120_),
    .Y(_04836_));
 NAND2x1_ASAP7_75t_R _22269_ (.A(net332),
    .B(_01118_),
    .Y(_04837_));
 OA211x2_ASAP7_75t_R _22270_ (.A1(net332),
    .A2(_04836_),
    .B(_04837_),
    .C(net356),
    .Y(_04838_));
 OR3x1_ASAP7_75t_R _22271_ (.A(net318),
    .B(_04835_),
    .C(_04838_),
    .Y(_04839_));
 OA211x2_ASAP7_75t_R _22272_ (.A1(_13598_),
    .A2(_04832_),
    .B(_04839_),
    .C(net325),
    .Y(_04840_));
 INVx1_ASAP7_75t_R _22273_ (.A(_01122_),
    .Y(_04841_));
 NOR2x1_ASAP7_75t_R _22274_ (.A(net332),
    .B(_01124_),
    .Y(_04842_));
 AO21x1_ASAP7_75t_R _22275_ (.A1(net332),
    .A2(_04841_),
    .B(_04842_),
    .Y(_04843_));
 INVx1_ASAP7_75t_R _22276_ (.A(_01125_),
    .Y(_04844_));
 NAND2x1_ASAP7_75t_R _22277_ (.A(net332),
    .B(_01123_),
    .Y(_04845_));
 OA211x2_ASAP7_75t_R _22278_ (.A1(net332),
    .A2(_04844_),
    .B(_04845_),
    .C(net308),
    .Y(_04846_));
 AO21x1_ASAP7_75t_R _22279_ (.A1(net356),
    .A2(_04843_),
    .B(_04846_),
    .Y(_04847_));
 INVx1_ASAP7_75t_R _22280_ (.A(_01117_),
    .Y(_04848_));
 NAND2x1_ASAP7_75t_R _22281_ (.A(net332),
    .B(_01115_),
    .Y(_04849_));
 OA211x2_ASAP7_75t_R _22282_ (.A1(net332),
    .A2(_04848_),
    .B(_04849_),
    .C(net308),
    .Y(_04850_));
 INVx1_ASAP7_75t_R _22283_ (.A(_01116_),
    .Y(_04851_));
 NAND2x1_ASAP7_75t_R _22284_ (.A(net332),
    .B(_01114_),
    .Y(_04852_));
 OA211x2_ASAP7_75t_R _22285_ (.A1(net332),
    .A2(_04851_),
    .B(_04852_),
    .C(net356),
    .Y(_04853_));
 OR3x1_ASAP7_75t_R _22286_ (.A(_13598_),
    .B(_04850_),
    .C(_04853_),
    .Y(_04854_));
 OA211x2_ASAP7_75t_R _22287_ (.A1(net318),
    .A2(_04847_),
    .B(_04854_),
    .C(_13132_),
    .Y(_04855_));
 OR3x2_ASAP7_75t_R _22288_ (.A(_13174_),
    .B(_04840_),
    .C(_04855_),
    .Y(_04856_));
 INVx1_ASAP7_75t_R _22289_ (.A(_01129_),
    .Y(_04857_));
 NAND2x1_ASAP7_75t_R _22290_ (.A(net331),
    .B(_01127_),
    .Y(_04858_));
 OA211x2_ASAP7_75t_R _22291_ (.A1(net331),
    .A2(_04857_),
    .B(_04858_),
    .C(net308),
    .Y(_04859_));
 INVx1_ASAP7_75t_R _22292_ (.A(_01128_),
    .Y(_04860_));
 NAND2x1_ASAP7_75t_R _22293_ (.A(net331),
    .B(_01126_),
    .Y(_04861_));
 OA211x2_ASAP7_75t_R _22294_ (.A1(net331),
    .A2(_04860_),
    .B(_04861_),
    .C(net357),
    .Y(_04862_));
 OR3x1_ASAP7_75t_R _22295_ (.A(_13132_),
    .B(_04859_),
    .C(_04862_),
    .Y(_04863_));
 INVx1_ASAP7_75t_R _22296_ (.A(_01133_),
    .Y(_04864_));
 NAND2x1_ASAP7_75t_R _22297_ (.A(net331),
    .B(_01131_),
    .Y(_04865_));
 OA211x2_ASAP7_75t_R _22298_ (.A1(net331),
    .A2(_04864_),
    .B(_04865_),
    .C(net308),
    .Y(_04866_));
 INVx1_ASAP7_75t_R _22299_ (.A(_01132_),
    .Y(_04867_));
 NAND2x1_ASAP7_75t_R _22300_ (.A(net331),
    .B(_01130_),
    .Y(_04868_));
 OA211x2_ASAP7_75t_R _22301_ (.A1(net331),
    .A2(_04867_),
    .B(_04868_),
    .C(net356),
    .Y(_04869_));
 OR3x1_ASAP7_75t_R _22302_ (.A(net325),
    .B(_04866_),
    .C(_04869_),
    .Y(_04870_));
 AND3x1_ASAP7_75t_R _22303_ (.A(net318),
    .B(_04863_),
    .C(_04870_),
    .Y(_04871_));
 INVx1_ASAP7_75t_R _22304_ (.A(_01137_),
    .Y(_04872_));
 NAND2x1_ASAP7_75t_R _22305_ (.A(net331),
    .B(_01135_),
    .Y(_04873_));
 OA211x2_ASAP7_75t_R _22306_ (.A1(net331),
    .A2(_04872_),
    .B(_04873_),
    .C(_13145_),
    .Y(_04874_));
 INVx1_ASAP7_75t_R _22307_ (.A(_01136_),
    .Y(_04875_));
 NAND2x1_ASAP7_75t_R _22308_ (.A(net331),
    .B(_01134_),
    .Y(_04876_));
 OA211x2_ASAP7_75t_R _22309_ (.A1(net331),
    .A2(_04875_),
    .B(_04876_),
    .C(net358),
    .Y(_04877_));
 OR3x1_ASAP7_75t_R _22310_ (.A(_13132_),
    .B(_04874_),
    .C(_04877_),
    .Y(_04878_));
 INVx1_ASAP7_75t_R _22311_ (.A(_01141_),
    .Y(_04879_));
 NAND2x1_ASAP7_75t_R _22312_ (.A(net331),
    .B(_01139_),
    .Y(_04880_));
 OA211x2_ASAP7_75t_R _22313_ (.A1(net331),
    .A2(_04879_),
    .B(_04880_),
    .C(_13145_),
    .Y(_04881_));
 INVx1_ASAP7_75t_R _22314_ (.A(_01140_),
    .Y(_04882_));
 NAND2x1_ASAP7_75t_R _22315_ (.A(net331),
    .B(_01138_),
    .Y(_04883_));
 OA211x2_ASAP7_75t_R _22316_ (.A1(net331),
    .A2(_04882_),
    .B(_04883_),
    .C(net358),
    .Y(_04884_));
 OR3x1_ASAP7_75t_R _22317_ (.A(net325),
    .B(_04881_),
    .C(_04884_),
    .Y(_04885_));
 AND3x1_ASAP7_75t_R _22318_ (.A(_13598_),
    .B(_04878_),
    .C(_04885_),
    .Y(_04886_));
 OR3x4_ASAP7_75t_R _22319_ (.A(net315),
    .B(_04871_),
    .C(_04886_),
    .Y(_04887_));
 NAND2x2_ASAP7_75t_R _22320_ (.A(_04856_),
    .B(_04887_),
    .Y(_04888_));
 OA21x2_ASAP7_75t_R _22321_ (.A1(_00283_),
    .A2(_15267_),
    .B(_16207_),
    .Y(_04889_));
 AOI21x1_ASAP7_75t_R _22322_ (.A1(_13583_),
    .A2(_04888_),
    .B(_04889_),
    .Y(_18236_));
 AND2x2_ASAP7_75t_R _22323_ (.A(net391),
    .B(_01683_),
    .Y(_04890_));
 AO21x1_ASAP7_75t_R _22324_ (.A1(net302),
    .A2(_01113_),
    .B(_04890_),
    .Y(_04891_));
 OAI22x1_ASAP7_75t_R _22325_ (.A1(_01112_),
    .A2(_13471_),
    .B1(_04891_),
    .B2(net409),
    .Y(_04892_));
 NAND2x1_ASAP7_75t_R _22326_ (.A(net390),
    .B(_01127_),
    .Y(_04893_));
 OA211x2_ASAP7_75t_R _22327_ (.A1(net390),
    .A2(_04857_),
    .B(_04893_),
    .C(_13424_),
    .Y(_04894_));
 NAND2x1_ASAP7_75t_R _22328_ (.A(net390),
    .B(_01126_),
    .Y(_04895_));
 OA211x2_ASAP7_75t_R _22329_ (.A1(net390),
    .A2(_04860_),
    .B(_04895_),
    .C(net408),
    .Y(_04896_));
 OR3x1_ASAP7_75t_R _22330_ (.A(net362),
    .B(_04894_),
    .C(_04896_),
    .Y(_04897_));
 OA211x2_ASAP7_75t_R _22331_ (.A1(_13392_),
    .A2(_04892_),
    .B(_04897_),
    .C(net370),
    .Y(_04898_));
 NAND2x1_ASAP7_75t_R _22332_ (.A(net391),
    .B(_01115_),
    .Y(_04899_));
 OA211x2_ASAP7_75t_R _22333_ (.A1(net391),
    .A2(_04848_),
    .B(_04899_),
    .C(net306),
    .Y(_04900_));
 NAND2x1_ASAP7_75t_R _22334_ (.A(net391),
    .B(_01114_),
    .Y(_04901_));
 OA211x2_ASAP7_75t_R _22335_ (.A1(net391),
    .A2(_04851_),
    .B(_04901_),
    .C(net409),
    .Y(_04902_));
 OR3x1_ASAP7_75t_R _22336_ (.A(_13392_),
    .B(_04900_),
    .C(_04902_),
    .Y(_04903_));
 NAND2x1_ASAP7_75t_R _22337_ (.A(net390),
    .B(_01131_),
    .Y(_04904_));
 OA211x2_ASAP7_75t_R _22338_ (.A1(net390),
    .A2(_04864_),
    .B(_04904_),
    .C(_13424_),
    .Y(_04905_));
 NAND2x1_ASAP7_75t_R _22339_ (.A(net390),
    .B(_01130_),
    .Y(_04906_));
 OA211x2_ASAP7_75t_R _22340_ (.A1(net390),
    .A2(_04867_),
    .B(_04906_),
    .C(net408),
    .Y(_04907_));
 OR3x1_ASAP7_75t_R _22341_ (.A(net362),
    .B(_04905_),
    .C(_04907_),
    .Y(_04908_));
 AND3x1_ASAP7_75t_R _22342_ (.A(_13397_),
    .B(_04903_),
    .C(_04908_),
    .Y(_04909_));
 OR3x4_ASAP7_75t_R _22343_ (.A(_13484_),
    .B(_04898_),
    .C(_04909_),
    .Y(_04910_));
 NAND2x1_ASAP7_75t_R _22344_ (.A(net390),
    .B(_01135_),
    .Y(_04911_));
 OA211x2_ASAP7_75t_R _22345_ (.A1(net390),
    .A2(_04872_),
    .B(_04911_),
    .C(_13424_),
    .Y(_04912_));
 NAND2x1_ASAP7_75t_R _22346_ (.A(net390),
    .B(_01134_),
    .Y(_04913_));
 OA211x2_ASAP7_75t_R _22347_ (.A1(net390),
    .A2(_04875_),
    .B(_04913_),
    .C(net408),
    .Y(_04914_));
 OR3x1_ASAP7_75t_R _22348_ (.A(_13397_),
    .B(_04912_),
    .C(_04914_),
    .Y(_04915_));
 NAND2x1_ASAP7_75t_R _22349_ (.A(net390),
    .B(_01139_),
    .Y(_04916_));
 OA211x2_ASAP7_75t_R _22350_ (.A1(net390),
    .A2(_04879_),
    .B(_04916_),
    .C(_13424_),
    .Y(_04917_));
 NAND2x1_ASAP7_75t_R _22351_ (.A(net390),
    .B(_01138_),
    .Y(_04918_));
 OA211x2_ASAP7_75t_R _22352_ (.A1(net390),
    .A2(_04882_),
    .B(_04918_),
    .C(net408),
    .Y(_04919_));
 OR3x1_ASAP7_75t_R _22353_ (.A(net372),
    .B(_04917_),
    .C(_04919_),
    .Y(_04920_));
 AND3x1_ASAP7_75t_R _22354_ (.A(_13392_),
    .B(_04915_),
    .C(_04920_),
    .Y(_04921_));
 NAND2x1_ASAP7_75t_R _22355_ (.A(net409),
    .B(_01120_),
    .Y(_04922_));
 OA211x2_ASAP7_75t_R _22356_ (.A1(net409),
    .A2(_04833_),
    .B(_04922_),
    .C(net370),
    .Y(_04923_));
 NAND2x1_ASAP7_75t_R _22357_ (.A(net409),
    .B(_01124_),
    .Y(_04924_));
 OA211x2_ASAP7_75t_R _22358_ (.A1(net409),
    .A2(_04844_),
    .B(_04924_),
    .C(_13397_),
    .Y(_04925_));
 OR3x1_ASAP7_75t_R _22359_ (.A(net391),
    .B(_04923_),
    .C(_04925_),
    .Y(_04926_));
 INVx1_ASAP7_75t_R _22360_ (.A(_01123_),
    .Y(_04927_));
 NAND2x1_ASAP7_75t_R _22361_ (.A(net370),
    .B(_01119_),
    .Y(_04928_));
 OA211x2_ASAP7_75t_R _22362_ (.A1(net370),
    .A2(_04927_),
    .B(_04928_),
    .C(net306),
    .Y(_04929_));
 NAND2x1_ASAP7_75t_R _22363_ (.A(net370),
    .B(_01118_),
    .Y(_04930_));
 OA211x2_ASAP7_75t_R _22364_ (.A1(net370),
    .A2(_04841_),
    .B(_04930_),
    .C(net409),
    .Y(_04931_));
 OR3x1_ASAP7_75t_R _22365_ (.A(net302),
    .B(_04929_),
    .C(_04931_),
    .Y(_04932_));
 AND3x1_ASAP7_75t_R _22366_ (.A(net362),
    .B(_04926_),
    .C(_04932_),
    .Y(_04933_));
 OR3x4_ASAP7_75t_R _22367_ (.A(net365),
    .B(_04921_),
    .C(_04933_),
    .Y(_04934_));
 NAND2x2_ASAP7_75t_R _22368_ (.A(_04910_),
    .B(_04934_),
    .Y(_04935_));
 OA22x2_ASAP7_75t_R _22369_ (.A1(_01615_),
    .A2(_13223_),
    .B1(_13880_),
    .B2(_00223_),
    .Y(_04936_));
 OAI21x1_ASAP7_75t_R _22370_ (.A1(_13782_),
    .A2(_04935_),
    .B(_04936_),
    .Y(_18235_));
 INVx1_ASAP7_75t_R _22371_ (.A(_18235_),
    .Y(_18237_));
 XNOR2x2_ASAP7_75t_R _22372_ (.A(_01145_),
    .B(_01143_),
    .Y(_04937_));
 INVx2_ASAP7_75t_R _22373_ (.A(_04937_),
    .Y(net167));
 AND2x2_ASAP7_75t_R _22374_ (.A(net334),
    .B(_01682_),
    .Y(_04938_));
 AO21x1_ASAP7_75t_R _22375_ (.A1(net313),
    .A2(_01147_),
    .B(_04938_),
    .Y(_04939_));
 OAI22x1_ASAP7_75t_R _22376_ (.A1(_01146_),
    .A2(_13586_),
    .B1(_04939_),
    .B2(net357),
    .Y(_04940_));
 INVx1_ASAP7_75t_R _22377_ (.A(_01155_),
    .Y(_04941_));
 NAND2x1_ASAP7_75t_R _22378_ (.A(net334),
    .B(_01153_),
    .Y(_04942_));
 OA211x2_ASAP7_75t_R _22379_ (.A1(net334),
    .A2(_04941_),
    .B(_04942_),
    .C(net308),
    .Y(_04943_));
 INVx1_ASAP7_75t_R _22380_ (.A(_01154_),
    .Y(_04944_));
 NAND2x1_ASAP7_75t_R _22381_ (.A(net334),
    .B(_01152_),
    .Y(_04945_));
 OA211x2_ASAP7_75t_R _22382_ (.A1(net334),
    .A2(_04944_),
    .B(_04945_),
    .C(net357),
    .Y(_04946_));
 OR3x1_ASAP7_75t_R _22383_ (.A(net319),
    .B(_04943_),
    .C(_04946_),
    .Y(_04947_));
 OA211x2_ASAP7_75t_R _22384_ (.A1(_13598_),
    .A2(_04940_),
    .B(_04947_),
    .C(net325),
    .Y(_04948_));
 INVx1_ASAP7_75t_R _22385_ (.A(_01151_),
    .Y(_04949_));
 NAND2x1_ASAP7_75t_R _22386_ (.A(net333),
    .B(_01149_),
    .Y(_04950_));
 OA211x2_ASAP7_75t_R _22387_ (.A1(net333),
    .A2(_04949_),
    .B(_04950_),
    .C(net308),
    .Y(_04951_));
 INVx1_ASAP7_75t_R _22388_ (.A(_01150_),
    .Y(_04952_));
 NAND2x1_ASAP7_75t_R _22389_ (.A(net333),
    .B(_01148_),
    .Y(_04953_));
 OA211x2_ASAP7_75t_R _22390_ (.A1(net333),
    .A2(_04952_),
    .B(_04953_),
    .C(net358),
    .Y(_04954_));
 OR3x1_ASAP7_75t_R _22391_ (.A(_13598_),
    .B(_04951_),
    .C(_04954_),
    .Y(_04955_));
 INVx1_ASAP7_75t_R _22392_ (.A(_01159_),
    .Y(_04956_));
 NAND2x1_ASAP7_75t_R _22393_ (.A(net333),
    .B(_01157_),
    .Y(_04957_));
 OA211x2_ASAP7_75t_R _22394_ (.A1(net333),
    .A2(_04956_),
    .B(_04957_),
    .C(net308),
    .Y(_04958_));
 INVx1_ASAP7_75t_R _22395_ (.A(_01158_),
    .Y(_04959_));
 NAND2x1_ASAP7_75t_R _22396_ (.A(net333),
    .B(_01156_),
    .Y(_04960_));
 OA211x2_ASAP7_75t_R _22397_ (.A1(net333),
    .A2(_04959_),
    .B(_04960_),
    .C(net357),
    .Y(_04961_));
 OR3x1_ASAP7_75t_R _22398_ (.A(net318),
    .B(_04958_),
    .C(_04961_),
    .Y(_04962_));
 AND3x1_ASAP7_75t_R _22399_ (.A(_13132_),
    .B(_04955_),
    .C(_04962_),
    .Y(_04963_));
 OR3x2_ASAP7_75t_R _22400_ (.A(_13174_),
    .B(_04948_),
    .C(_04963_),
    .Y(_04964_));
 INVx1_ASAP7_75t_R _22401_ (.A(_01167_),
    .Y(_04965_));
 NAND2x1_ASAP7_75t_R _22402_ (.A(net333),
    .B(_01165_),
    .Y(_04966_));
 OA211x2_ASAP7_75t_R _22403_ (.A1(net333),
    .A2(_04965_),
    .B(_04966_),
    .C(_13145_),
    .Y(_04967_));
 INVx1_ASAP7_75t_R _22404_ (.A(_01166_),
    .Y(_04968_));
 NAND2x1_ASAP7_75t_R _22405_ (.A(net333),
    .B(_01164_),
    .Y(_04969_));
 OA211x2_ASAP7_75t_R _22406_ (.A1(net333),
    .A2(_04968_),
    .B(_04969_),
    .C(net358),
    .Y(_04970_));
 OR3x1_ASAP7_75t_R _22407_ (.A(_13598_),
    .B(_04967_),
    .C(_04970_),
    .Y(_04971_));
 INVx1_ASAP7_75t_R _22408_ (.A(_01175_),
    .Y(_04972_));
 NAND2x1_ASAP7_75t_R _22409_ (.A(net333),
    .B(_01173_),
    .Y(_04973_));
 OA211x2_ASAP7_75t_R _22410_ (.A1(net333),
    .A2(_04972_),
    .B(_04973_),
    .C(_13145_),
    .Y(_04974_));
 INVx1_ASAP7_75t_R _22411_ (.A(_01174_),
    .Y(_04975_));
 NAND2x1_ASAP7_75t_R _22412_ (.A(net333),
    .B(_01172_),
    .Y(_04976_));
 OA211x2_ASAP7_75t_R _22413_ (.A1(net333),
    .A2(_04975_),
    .B(_04976_),
    .C(net358),
    .Y(_04977_));
 OR3x1_ASAP7_75t_R _22414_ (.A(net318),
    .B(_04974_),
    .C(_04977_),
    .Y(_04978_));
 AND3x1_ASAP7_75t_R _22415_ (.A(_13132_),
    .B(_04971_),
    .C(_04978_),
    .Y(_04979_));
 INVx1_ASAP7_75t_R _22416_ (.A(_01168_),
    .Y(_04980_));
 NOR2x1_ASAP7_75t_R _22417_ (.A(net333),
    .B(_01170_),
    .Y(_04981_));
 AO21x1_ASAP7_75t_R _22418_ (.A1(net333),
    .A2(_04980_),
    .B(_04981_),
    .Y(_04982_));
 INVx1_ASAP7_75t_R _22419_ (.A(_01171_),
    .Y(_04983_));
 NAND2x1_ASAP7_75t_R _22420_ (.A(net333),
    .B(_01169_),
    .Y(_04984_));
 OA211x2_ASAP7_75t_R _22421_ (.A1(net333),
    .A2(_04983_),
    .B(_04984_),
    .C(_13145_),
    .Y(_04985_));
 AO21x1_ASAP7_75t_R _22422_ (.A1(net358),
    .A2(_04982_),
    .B(_04985_),
    .Y(_04986_));
 INVx1_ASAP7_75t_R _22423_ (.A(_01163_),
    .Y(_04987_));
 NAND2x1_ASAP7_75t_R _22424_ (.A(net333),
    .B(_01161_),
    .Y(_04988_));
 OA211x2_ASAP7_75t_R _22425_ (.A1(net333),
    .A2(_04987_),
    .B(_04988_),
    .C(_13145_),
    .Y(_04989_));
 INVx1_ASAP7_75t_R _22426_ (.A(_01162_),
    .Y(_04990_));
 NAND2x1_ASAP7_75t_R _22427_ (.A(net333),
    .B(_01160_),
    .Y(_04991_));
 OA211x2_ASAP7_75t_R _22428_ (.A1(net333),
    .A2(_04990_),
    .B(_04991_),
    .C(net358),
    .Y(_04992_));
 OR3x1_ASAP7_75t_R _22429_ (.A(_13598_),
    .B(_04989_),
    .C(_04992_),
    .Y(_04993_));
 OA211x2_ASAP7_75t_R _22430_ (.A1(net318),
    .A2(_04986_),
    .B(_04993_),
    .C(net325),
    .Y(_04994_));
 OR3x4_ASAP7_75t_R _22431_ (.A(net315),
    .B(_04979_),
    .C(_04994_),
    .Y(_04995_));
 NAND2x2_ASAP7_75t_R _22432_ (.A(_04964_),
    .B(_04995_),
    .Y(_04996_));
 OA21x2_ASAP7_75t_R _22433_ (.A1(_01742_),
    .A2(_15267_),
    .B(_16207_),
    .Y(_04997_));
 AO21x2_ASAP7_75t_R _22434_ (.A1(_13583_),
    .A2(_04996_),
    .B(_04997_),
    .Y(_04998_));
 BUFx2_ASAP7_75t_R output233 (.A(net233),
    .Y(instr_addr_o[24]));
 INVx1_ASAP7_75t_R _22436_ (.A(_04998_),
    .Y(_18241_));
 INVx3_ASAP7_75t_R _22437_ (.A(_00224_),
    .Y(\cs_registers_i.pc_id_i[27] ));
 INVx1_ASAP7_75t_R _22438_ (.A(_01614_),
    .Y(_04999_));
 NAND2x1_ASAP7_75t_R _22439_ (.A(net394),
    .B(_01153_),
    .Y(_05000_));
 OA211x2_ASAP7_75t_R _22440_ (.A1(net394),
    .A2(_04941_),
    .B(_05000_),
    .C(net306),
    .Y(_05001_));
 NAND2x1_ASAP7_75t_R _22441_ (.A(net394),
    .B(_01152_),
    .Y(_05002_));
 OA211x2_ASAP7_75t_R _22442_ (.A1(net394),
    .A2(_04944_),
    .B(_05002_),
    .C(net410),
    .Y(_05003_));
 INVx1_ASAP7_75t_R _22443_ (.A(_01147_),
    .Y(_05004_));
 NAND2x1_ASAP7_75t_R _22444_ (.A(net394),
    .B(_01682_),
    .Y(_05005_));
 OA211x2_ASAP7_75t_R _22445_ (.A1(net394),
    .A2(_05004_),
    .B(_05005_),
    .C(net306),
    .Y(_05006_));
 NOR2x1_ASAP7_75t_R _22446_ (.A(_01146_),
    .B(_13471_),
    .Y(_05007_));
 OA33x2_ASAP7_75t_R _22447_ (.A1(_14743_),
    .A2(_05001_),
    .A3(_05003_),
    .B1(_05006_),
    .B2(_05007_),
    .B3(_13828_),
    .Y(_05008_));
 NAND2x1_ASAP7_75t_R _22448_ (.A(net393),
    .B(_01149_),
    .Y(_05009_));
 OA211x2_ASAP7_75t_R _22449_ (.A1(net393),
    .A2(_04949_),
    .B(_05009_),
    .C(net306),
    .Y(_05010_));
 NAND2x1_ASAP7_75t_R _22450_ (.A(net393),
    .B(_01148_),
    .Y(_05011_));
 OA211x2_ASAP7_75t_R _22451_ (.A1(net393),
    .A2(_04952_),
    .B(_05011_),
    .C(net408),
    .Y(_05012_));
 OR3x1_ASAP7_75t_R _22452_ (.A(_13484_),
    .B(_05010_),
    .C(_05012_),
    .Y(_05013_));
 NAND2x1_ASAP7_75t_R _22453_ (.A(net393),
    .B(_01157_),
    .Y(_05014_));
 OA211x2_ASAP7_75t_R _22454_ (.A1(net393),
    .A2(_04956_),
    .B(_05014_),
    .C(net306),
    .Y(_05015_));
 NAND2x1_ASAP7_75t_R _22455_ (.A(net393),
    .B(_01156_),
    .Y(_05016_));
 OA211x2_ASAP7_75t_R _22456_ (.A1(net393),
    .A2(_04959_),
    .B(_05016_),
    .C(net408),
    .Y(_05017_));
 OR3x1_ASAP7_75t_R _22457_ (.A(net365),
    .B(_05015_),
    .C(_05017_),
    .Y(_05018_));
 AO21x1_ASAP7_75t_R _22458_ (.A1(_05013_),
    .A2(_05018_),
    .B(net372),
    .Y(_05019_));
 AO21x1_ASAP7_75t_R _22459_ (.A1(_05008_),
    .A2(_05019_),
    .B(_13392_),
    .Y(_05020_));
 NAND2x1_ASAP7_75t_R _22460_ (.A(_13424_),
    .B(_01169_),
    .Y(_05021_));
 OA211x2_ASAP7_75t_R _22461_ (.A1(_13424_),
    .A2(_04980_),
    .B(_05021_),
    .C(net372),
    .Y(_05022_));
 AND2x2_ASAP7_75t_R _22462_ (.A(net408),
    .B(_01172_),
    .Y(_05023_));
 AO21x1_ASAP7_75t_R _22463_ (.A1(_13424_),
    .A2(_01173_),
    .B(_05023_),
    .Y(_05024_));
 OAI21x1_ASAP7_75t_R _22464_ (.A1(net372),
    .A2(_05024_),
    .B(net394),
    .Y(_05025_));
 NAND2x1_ASAP7_75t_R _22465_ (.A(net408),
    .B(_01174_),
    .Y(_05026_));
 OA211x2_ASAP7_75t_R _22466_ (.A1(net408),
    .A2(_04972_),
    .B(_05026_),
    .C(_13397_),
    .Y(_05027_));
 NAND2x1_ASAP7_75t_R _22467_ (.A(net408),
    .B(_01170_),
    .Y(_05028_));
 OA211x2_ASAP7_75t_R _22468_ (.A1(net408),
    .A2(_04983_),
    .B(_05028_),
    .C(net372),
    .Y(_05029_));
 OR3x1_ASAP7_75t_R _22469_ (.A(net394),
    .B(_05027_),
    .C(_05029_),
    .Y(_05030_));
 OA211x2_ASAP7_75t_R _22470_ (.A1(_05022_),
    .A2(_05025_),
    .B(_05030_),
    .C(_13484_),
    .Y(_05031_));
 NAND2x1_ASAP7_75t_R _22471_ (.A(net393),
    .B(_01164_),
    .Y(_05032_));
 OA211x2_ASAP7_75t_R _22472_ (.A1(net393),
    .A2(_04968_),
    .B(_05032_),
    .C(_13397_),
    .Y(_05033_));
 NAND2x1_ASAP7_75t_R _22473_ (.A(net393),
    .B(_01160_),
    .Y(_05034_));
 OA211x2_ASAP7_75t_R _22474_ (.A1(net393),
    .A2(_04990_),
    .B(_05034_),
    .C(net372),
    .Y(_05035_));
 OR3x1_ASAP7_75t_R _22475_ (.A(_13424_),
    .B(_05033_),
    .C(_05035_),
    .Y(_05036_));
 NAND2x1_ASAP7_75t_R _22476_ (.A(net393),
    .B(_01165_),
    .Y(_05037_));
 OA211x2_ASAP7_75t_R _22477_ (.A1(net393),
    .A2(_04965_),
    .B(_05037_),
    .C(_13397_),
    .Y(_05038_));
 NAND2x1_ASAP7_75t_R _22478_ (.A(net393),
    .B(_01161_),
    .Y(_05039_));
 OA211x2_ASAP7_75t_R _22479_ (.A1(net393),
    .A2(_04987_),
    .B(_05039_),
    .C(net372),
    .Y(_05040_));
 OR3x1_ASAP7_75t_R _22480_ (.A(net408),
    .B(_05038_),
    .C(_05040_),
    .Y(_05041_));
 AND3x1_ASAP7_75t_R _22481_ (.A(net365),
    .B(_05036_),
    .C(_05041_),
    .Y(_05042_));
 OR3x4_ASAP7_75t_R _22482_ (.A(net364),
    .B(_05031_),
    .C(_05042_),
    .Y(_05043_));
 AND2x4_ASAP7_75t_R _22483_ (.A(_05020_),
    .B(_05043_),
    .Y(_05044_));
 AO222x2_ASAP7_75t_R _22484_ (.A1(_04999_),
    .A2(_13270_),
    .B1(_13563_),
    .B2(_05044_),
    .C1(_14503_),
    .C2(\cs_registers_i.pc_id_i[27] ),
    .Y(_05045_));
 BUFx2_ASAP7_75t_R output232 (.A(net232),
    .Y(instr_addr_o[23]));
 INVx1_ASAP7_75t_R _22486_ (.A(_05045_),
    .Y(_18242_));
 BUFx2_ASAP7_75t_R output231 (.A(net231),
    .Y(instr_addr_o[22]));
 AND2x2_ASAP7_75t_R _22488_ (.A(net351),
    .B(_01681_),
    .Y(_05047_));
 AO21x1_ASAP7_75t_R _22489_ (.A1(_13127_),
    .A2(_01179_),
    .B(_05047_),
    .Y(_05048_));
 OAI22x1_ASAP7_75t_R _22490_ (.A1(_01178_),
    .A2(_13586_),
    .B1(_05048_),
    .B2(net360),
    .Y(_05049_));
 INVx1_ASAP7_75t_R _22491_ (.A(_01187_),
    .Y(_05050_));
 NAND2x1_ASAP7_75t_R _22492_ (.A(net351),
    .B(_01185_),
    .Y(_05051_));
 OA211x2_ASAP7_75t_R _22493_ (.A1(net351),
    .A2(_05050_),
    .B(_05051_),
    .C(net309),
    .Y(_05052_));
 INVx1_ASAP7_75t_R _22494_ (.A(_01186_),
    .Y(_05053_));
 NAND2x1_ASAP7_75t_R _22495_ (.A(net351),
    .B(_01184_),
    .Y(_05054_));
 OA211x2_ASAP7_75t_R _22496_ (.A1(net351),
    .A2(_05053_),
    .B(_05054_),
    .C(net360),
    .Y(_05055_));
 OR3x1_ASAP7_75t_R _22497_ (.A(net320),
    .B(_05052_),
    .C(_05055_),
    .Y(_05056_));
 OA21x2_ASAP7_75t_R _22498_ (.A1(_13598_),
    .A2(_05049_),
    .B(_05056_),
    .Y(_05057_));
 INVx1_ASAP7_75t_R _22499_ (.A(_01183_),
    .Y(_05058_));
 NAND2x1_ASAP7_75t_R _22500_ (.A(net353),
    .B(_01181_),
    .Y(_05059_));
 OA211x2_ASAP7_75t_R _22501_ (.A1(net353),
    .A2(_05058_),
    .B(_05059_),
    .C(net309),
    .Y(_05060_));
 INVx1_ASAP7_75t_R _22502_ (.A(_01182_),
    .Y(_05061_));
 NAND2x1_ASAP7_75t_R _22503_ (.A(net353),
    .B(_01180_),
    .Y(_05062_));
 OA211x2_ASAP7_75t_R _22504_ (.A1(net353),
    .A2(_05061_),
    .B(_05062_),
    .C(net361),
    .Y(_05063_));
 OR3x1_ASAP7_75t_R _22505_ (.A(_13598_),
    .B(_05060_),
    .C(_05063_),
    .Y(_05064_));
 INVx1_ASAP7_75t_R _22506_ (.A(_01191_),
    .Y(_05065_));
 NAND2x1_ASAP7_75t_R _22507_ (.A(net353),
    .B(_01189_),
    .Y(_05066_));
 OA211x2_ASAP7_75t_R _22508_ (.A1(net353),
    .A2(_05065_),
    .B(_05066_),
    .C(net309),
    .Y(_05067_));
 INVx1_ASAP7_75t_R _22509_ (.A(_01190_),
    .Y(_05068_));
 NAND2x1_ASAP7_75t_R _22510_ (.A(net353),
    .B(_01188_),
    .Y(_05069_));
 OA211x2_ASAP7_75t_R _22511_ (.A1(net353),
    .A2(_05068_),
    .B(_05069_),
    .C(net361),
    .Y(_05070_));
 OR3x1_ASAP7_75t_R _22512_ (.A(_00245_),
    .B(_05067_),
    .C(_05070_),
    .Y(_05071_));
 AND3x1_ASAP7_75t_R _22513_ (.A(_13132_),
    .B(_05064_),
    .C(_05071_),
    .Y(_05072_));
 AO21x1_ASAP7_75t_R _22514_ (.A1(_01744_),
    .A2(_05057_),
    .B(_05072_),
    .Y(_05073_));
 INVx1_ASAP7_75t_R _22515_ (.A(_01199_),
    .Y(_05074_));
 NAND2x1_ASAP7_75t_R _22516_ (.A(net352),
    .B(_01197_),
    .Y(_05075_));
 OA211x2_ASAP7_75t_R _22517_ (.A1(net352),
    .A2(_05074_),
    .B(_05075_),
    .C(net309),
    .Y(_05076_));
 INVx1_ASAP7_75t_R _22518_ (.A(_01198_),
    .Y(_05077_));
 NAND2x1_ASAP7_75t_R _22519_ (.A(net352),
    .B(_01196_),
    .Y(_05078_));
 OA211x2_ASAP7_75t_R _22520_ (.A1(net352),
    .A2(_05077_),
    .B(_05078_),
    .C(net361),
    .Y(_05079_));
 OR3x1_ASAP7_75t_R _22521_ (.A(_13598_),
    .B(_05076_),
    .C(_05079_),
    .Y(_05080_));
 INVx1_ASAP7_75t_R _22522_ (.A(_01207_),
    .Y(_05081_));
 NAND2x1_ASAP7_75t_R _22523_ (.A(net351),
    .B(_01205_),
    .Y(_05082_));
 OA211x2_ASAP7_75t_R _22524_ (.A1(net352),
    .A2(_05081_),
    .B(_05082_),
    .C(net309),
    .Y(_05083_));
 INVx1_ASAP7_75t_R _22525_ (.A(_01206_),
    .Y(_05084_));
 NAND2x1_ASAP7_75t_R _22526_ (.A(net352),
    .B(_01204_),
    .Y(_05085_));
 OA211x2_ASAP7_75t_R _22527_ (.A1(net352),
    .A2(_05084_),
    .B(_05085_),
    .C(net361),
    .Y(_05086_));
 OR3x1_ASAP7_75t_R _22528_ (.A(_00245_),
    .B(_05083_),
    .C(_05086_),
    .Y(_05087_));
 AND3x1_ASAP7_75t_R _22529_ (.A(_13132_),
    .B(_05080_),
    .C(_05087_),
    .Y(_05088_));
 INVx1_ASAP7_75t_R _22530_ (.A(_01195_),
    .Y(_05089_));
 NAND2x1_ASAP7_75t_R _22531_ (.A(net351),
    .B(_01193_),
    .Y(_05090_));
 OA211x2_ASAP7_75t_R _22532_ (.A1(net351),
    .A2(_05089_),
    .B(_05090_),
    .C(net309),
    .Y(_05091_));
 INVx1_ASAP7_75t_R _22533_ (.A(_01194_),
    .Y(_05092_));
 NAND2x1_ASAP7_75t_R _22534_ (.A(net351),
    .B(_01192_),
    .Y(_05093_));
 OA211x2_ASAP7_75t_R _22535_ (.A1(net351),
    .A2(_05092_),
    .B(_05093_),
    .C(net360),
    .Y(_05094_));
 OR3x1_ASAP7_75t_R _22536_ (.A(_13598_),
    .B(_05091_),
    .C(_05094_),
    .Y(_05095_));
 INVx1_ASAP7_75t_R _22537_ (.A(_01203_),
    .Y(_05096_));
 NAND2x1_ASAP7_75t_R _22538_ (.A(net351),
    .B(_01201_),
    .Y(_05097_));
 OA211x2_ASAP7_75t_R _22539_ (.A1(net351),
    .A2(_05096_),
    .B(_05097_),
    .C(net309),
    .Y(_05098_));
 INVx1_ASAP7_75t_R _22540_ (.A(_01202_),
    .Y(_05099_));
 NAND2x1_ASAP7_75t_R _22541_ (.A(net351),
    .B(_01200_),
    .Y(_05100_));
 OA211x2_ASAP7_75t_R _22542_ (.A1(net351),
    .A2(_05099_),
    .B(_05100_),
    .C(net360),
    .Y(_05101_));
 OR3x1_ASAP7_75t_R _22543_ (.A(_00245_),
    .B(_05098_),
    .C(_05101_),
    .Y(_05102_));
 AND3x1_ASAP7_75t_R _22544_ (.A(_01744_),
    .B(_05095_),
    .C(_05102_),
    .Y(_05103_));
 OR3x1_ASAP7_75t_R _22545_ (.A(net316),
    .B(_05088_),
    .C(_05103_),
    .Y(_05104_));
 OAI21x1_ASAP7_75t_R _22546_ (.A1(_13174_),
    .A2(_05073_),
    .B(_05104_),
    .Y(_05105_));
 OA21x2_ASAP7_75t_R _22547_ (.A1(_01741_),
    .A2(_15267_),
    .B(_16207_),
    .Y(_05106_));
 AO21x2_ASAP7_75t_R _22548_ (.A1(_13583_),
    .A2(_05105_),
    .B(_05106_),
    .Y(_05107_));
 BUFx2_ASAP7_75t_R output230 (.A(net230),
    .Y(instr_addr_o[21]));
 INVx1_ASAP7_75t_R _22550_ (.A(_05107_),
    .Y(_18247_));
 AND2x2_ASAP7_75t_R _22551_ (.A(_00226_),
    .B(_13553_),
    .Y(_05108_));
 NAND2x1_ASAP7_75t_R _22552_ (.A(net379),
    .B(_01181_),
    .Y(_05109_));
 OA211x2_ASAP7_75t_R _22553_ (.A1(net379),
    .A2(_05058_),
    .B(_05109_),
    .C(net304),
    .Y(_05110_));
 NAND2x1_ASAP7_75t_R _22554_ (.A(net403),
    .B(_01180_),
    .Y(_05111_));
 OA211x2_ASAP7_75t_R _22555_ (.A1(net403),
    .A2(_05061_),
    .B(_05111_),
    .C(_00290_),
    .Y(_05112_));
 OR3x1_ASAP7_75t_R _22556_ (.A(_13484_),
    .B(_05110_),
    .C(_05112_),
    .Y(_05113_));
 NAND2x1_ASAP7_75t_R _22557_ (.A(net403),
    .B(_01189_),
    .Y(_05114_));
 OA211x2_ASAP7_75t_R _22558_ (.A1(net403),
    .A2(_05065_),
    .B(_05114_),
    .C(net304),
    .Y(_05115_));
 NAND2x1_ASAP7_75t_R _22559_ (.A(net403),
    .B(_01188_),
    .Y(_05116_));
 OA211x2_ASAP7_75t_R _22560_ (.A1(net403),
    .A2(_05068_),
    .B(_05116_),
    .C(_00290_),
    .Y(_05117_));
 OR3x1_ASAP7_75t_R _22561_ (.A(_00287_),
    .B(_05115_),
    .C(_05117_),
    .Y(_05118_));
 AO21x1_ASAP7_75t_R _22562_ (.A1(_05113_),
    .A2(_05118_),
    .B(net374),
    .Y(_05119_));
 AND2x2_ASAP7_75t_R _22563_ (.A(_00289_),
    .B(_01681_),
    .Y(_05120_));
 AO21x1_ASAP7_75t_R _22564_ (.A1(_13433_),
    .A2(_01179_),
    .B(_05120_),
    .Y(_05121_));
 OAI22x1_ASAP7_75t_R _22565_ (.A1(_01178_),
    .A2(_13471_),
    .B1(_05121_),
    .B2(_00290_),
    .Y(_05122_));
 NAND2x1_ASAP7_75t_R _22566_ (.A(net402),
    .B(_01185_),
    .Y(_05123_));
 OA211x2_ASAP7_75t_R _22567_ (.A1(net402),
    .A2(_05050_),
    .B(_05123_),
    .C(net305),
    .Y(_05124_));
 NAND2x1_ASAP7_75t_R _22568_ (.A(net402),
    .B(_01184_),
    .Y(_05125_));
 OA211x2_ASAP7_75t_R _22569_ (.A1(net402),
    .A2(_05053_),
    .B(_05125_),
    .C(_00290_),
    .Y(_05126_));
 OR3x1_ASAP7_75t_R _22570_ (.A(_14743_),
    .B(_05124_),
    .C(_05126_),
    .Y(_05127_));
 OA211x2_ASAP7_75t_R _22571_ (.A1(net300),
    .A2(_05122_),
    .B(_05127_),
    .C(_00286_),
    .Y(_05128_));
 NAND2x1_ASAP7_75t_R _22572_ (.A(net402),
    .B(_01201_),
    .Y(_05129_));
 OA211x2_ASAP7_75t_R _22573_ (.A1(net402),
    .A2(_05096_),
    .B(_05129_),
    .C(net305),
    .Y(_05130_));
 NAND2x1_ASAP7_75t_R _22574_ (.A(net402),
    .B(_01200_),
    .Y(_05131_));
 OA211x2_ASAP7_75t_R _22575_ (.A1(net402),
    .A2(_05099_),
    .B(_05131_),
    .C(_00290_),
    .Y(_05132_));
 OR3x1_ASAP7_75t_R _22576_ (.A(_13397_),
    .B(_05130_),
    .C(_05132_),
    .Y(_05133_));
 NAND2x1_ASAP7_75t_R _22577_ (.A(net402),
    .B(_01205_),
    .Y(_05134_));
 OA211x2_ASAP7_75t_R _22578_ (.A1(net402),
    .A2(_05081_),
    .B(_05134_),
    .C(net305),
    .Y(_05135_));
 NAND2x1_ASAP7_75t_R _22579_ (.A(net402),
    .B(_01204_),
    .Y(_05136_));
 OA211x2_ASAP7_75t_R _22580_ (.A1(net402),
    .A2(_05084_),
    .B(_05136_),
    .C(_00290_),
    .Y(_05137_));
 OR3x1_ASAP7_75t_R _22581_ (.A(net374),
    .B(_05135_),
    .C(_05137_),
    .Y(_05138_));
 AO21x1_ASAP7_75t_R _22582_ (.A1(_05133_),
    .A2(_05138_),
    .B(_00287_),
    .Y(_05139_));
 NAND2x1_ASAP7_75t_R _22583_ (.A(net403),
    .B(_01197_),
    .Y(_05140_));
 OA211x2_ASAP7_75t_R _22584_ (.A1(net403),
    .A2(_05074_),
    .B(_05140_),
    .C(net305),
    .Y(_05141_));
 NAND2x1_ASAP7_75t_R _22585_ (.A(net403),
    .B(_01196_),
    .Y(_05142_));
 OA211x2_ASAP7_75t_R _22586_ (.A1(net403),
    .A2(_05077_),
    .B(_05142_),
    .C(_00290_),
    .Y(_05143_));
 OR3x1_ASAP7_75t_R _22587_ (.A(net298),
    .B(_05141_),
    .C(_05143_),
    .Y(_05144_));
 NAND2x1_ASAP7_75t_R _22588_ (.A(net402),
    .B(_01193_),
    .Y(_05145_));
 OA211x2_ASAP7_75t_R _22589_ (.A1(net402),
    .A2(_05089_),
    .B(_05145_),
    .C(net307),
    .Y(_05146_));
 NAND2x1_ASAP7_75t_R _22590_ (.A(_00289_),
    .B(_01192_),
    .Y(_05147_));
 OA211x2_ASAP7_75t_R _22591_ (.A1(_00289_),
    .A2(_05092_),
    .B(_05147_),
    .C(_00290_),
    .Y(_05148_));
 OR3x1_ASAP7_75t_R _22592_ (.A(net300),
    .B(_05146_),
    .C(_05148_),
    .Y(_05149_));
 AND3x1_ASAP7_75t_R _22593_ (.A(_13392_),
    .B(_05144_),
    .C(_05149_),
    .Y(_05150_));
 AOI221x1_ASAP7_75t_R _22594_ (.A1(_05119_),
    .A2(_05128_),
    .B1(_05139_),
    .B2(_05150_),
    .C(_13553_),
    .Y(_05151_));
 OR3x1_ASAP7_75t_R _22595_ (.A(_13561_),
    .B(_05108_),
    .C(_05151_),
    .Y(_05152_));
 AO21x1_ASAP7_75t_R _22596_ (.A1(_13219_),
    .A2(_13222_),
    .B(_01613_),
    .Y(_05153_));
 NAND2x2_ASAP7_75t_R _22597_ (.A(_05152_),
    .B(_05153_),
    .Y(_18248_));
 INVx4_ASAP7_75t_R _22598_ (.A(_18248_),
    .Y(_18246_));
 XNOR2x2_ASAP7_75t_R _22599_ (.A(_01211_),
    .B(_01209_),
    .Y(_05154_));
 INVx3_ASAP7_75t_R _22600_ (.A(_05154_),
    .Y(net169));
 AND2x2_ASAP7_75t_R _22601_ (.A(net338),
    .B(_01680_),
    .Y(_05155_));
 AO21x1_ASAP7_75t_R _22602_ (.A1(net313),
    .A2(_01213_),
    .B(_05155_),
    .Y(_05156_));
 OAI22x1_ASAP7_75t_R _22603_ (.A1(_01212_),
    .A2(_13586_),
    .B1(_05156_),
    .B2(net358),
    .Y(_05157_));
 INVx1_ASAP7_75t_R _22604_ (.A(_01221_),
    .Y(_05158_));
 NAND2x1_ASAP7_75t_R _22605_ (.A(net338),
    .B(_01219_),
    .Y(_05159_));
 OA211x2_ASAP7_75t_R _22606_ (.A1(net338),
    .A2(_05158_),
    .B(_05159_),
    .C(net308),
    .Y(_05160_));
 INVx1_ASAP7_75t_R _22607_ (.A(_01220_),
    .Y(_05161_));
 NAND2x1_ASAP7_75t_R _22608_ (.A(net338),
    .B(_01218_),
    .Y(_05162_));
 OA211x2_ASAP7_75t_R _22609_ (.A1(net338),
    .A2(_05161_),
    .B(_05162_),
    .C(net359),
    .Y(_05163_));
 OR3x1_ASAP7_75t_R _22610_ (.A(net319),
    .B(_05160_),
    .C(_05163_),
    .Y(_05164_));
 OA211x2_ASAP7_75t_R _22611_ (.A1(_13598_),
    .A2(_05157_),
    .B(_05164_),
    .C(net325),
    .Y(_05165_));
 INVx1_ASAP7_75t_R _22612_ (.A(_01217_),
    .Y(_05166_));
 NAND2x1_ASAP7_75t_R _22613_ (.A(net338),
    .B(_01215_),
    .Y(_05167_));
 OA211x2_ASAP7_75t_R _22614_ (.A1(net338),
    .A2(_05166_),
    .B(_05167_),
    .C(net308),
    .Y(_05168_));
 INVx1_ASAP7_75t_R _22615_ (.A(_01216_),
    .Y(_05169_));
 NAND2x1_ASAP7_75t_R _22616_ (.A(net338),
    .B(_01214_),
    .Y(_05170_));
 OA211x2_ASAP7_75t_R _22617_ (.A1(net338),
    .A2(_05169_),
    .B(_05170_),
    .C(net358),
    .Y(_05171_));
 OR3x1_ASAP7_75t_R _22618_ (.A(_13598_),
    .B(_05168_),
    .C(_05171_),
    .Y(_05172_));
 INVx1_ASAP7_75t_R _22619_ (.A(_01225_),
    .Y(_05173_));
 NAND2x1_ASAP7_75t_R _22620_ (.A(net338),
    .B(_01223_),
    .Y(_05174_));
 OA211x2_ASAP7_75t_R _22621_ (.A1(net338),
    .A2(_05173_),
    .B(_05174_),
    .C(net308),
    .Y(_05175_));
 INVx1_ASAP7_75t_R _22622_ (.A(_01224_),
    .Y(_05176_));
 NAND2x1_ASAP7_75t_R _22623_ (.A(net338),
    .B(_01222_),
    .Y(_05177_));
 OA211x2_ASAP7_75t_R _22624_ (.A1(net338),
    .A2(_05176_),
    .B(_05177_),
    .C(net359),
    .Y(_05178_));
 OR3x1_ASAP7_75t_R _22625_ (.A(net319),
    .B(_05175_),
    .C(_05178_),
    .Y(_05179_));
 AND3x1_ASAP7_75t_R _22626_ (.A(_13132_),
    .B(_05172_),
    .C(_05179_),
    .Y(_05180_));
 OR3x2_ASAP7_75t_R _22627_ (.A(_13174_),
    .B(_05165_),
    .C(_05180_),
    .Y(_05181_));
 INVx1_ASAP7_75t_R _22628_ (.A(_01233_),
    .Y(_05182_));
 NAND2x1_ASAP7_75t_R _22629_ (.A(net337),
    .B(_01231_),
    .Y(_05183_));
 OA211x2_ASAP7_75t_R _22630_ (.A1(net337),
    .A2(_05182_),
    .B(_05183_),
    .C(net308),
    .Y(_05184_));
 INVx1_ASAP7_75t_R _22631_ (.A(_01232_),
    .Y(_05185_));
 NAND2x1_ASAP7_75t_R _22632_ (.A(net337),
    .B(_01230_),
    .Y(_05186_));
 OA211x2_ASAP7_75t_R _22633_ (.A1(net337),
    .A2(_05185_),
    .B(_05186_),
    .C(net358),
    .Y(_05187_));
 OR3x1_ASAP7_75t_R _22634_ (.A(net325),
    .B(_05184_),
    .C(_05187_),
    .Y(_05188_));
 INVx1_ASAP7_75t_R _22635_ (.A(_01229_),
    .Y(_05189_));
 NAND2x1_ASAP7_75t_R _22636_ (.A(net337),
    .B(_01227_),
    .Y(_05190_));
 OA211x2_ASAP7_75t_R _22637_ (.A1(net337),
    .A2(_05189_),
    .B(_05190_),
    .C(net308),
    .Y(_05191_));
 INVx1_ASAP7_75t_R _22638_ (.A(_01228_),
    .Y(_05192_));
 NAND2x1_ASAP7_75t_R _22639_ (.A(net338),
    .B(_01226_),
    .Y(_05193_));
 OA211x2_ASAP7_75t_R _22640_ (.A1(net338),
    .A2(_05192_),
    .B(_05193_),
    .C(net358),
    .Y(_05194_));
 OR3x1_ASAP7_75t_R _22641_ (.A(_13132_),
    .B(_05191_),
    .C(_05194_),
    .Y(_05195_));
 AND3x1_ASAP7_75t_R _22642_ (.A(net319),
    .B(_05188_),
    .C(_05195_),
    .Y(_05196_));
 INVx1_ASAP7_75t_R _22643_ (.A(_01236_),
    .Y(_05197_));
 NAND2x1_ASAP7_75t_R _22644_ (.A(net338),
    .B(_01234_),
    .Y(_05198_));
 OA211x2_ASAP7_75t_R _22645_ (.A1(net338),
    .A2(_05197_),
    .B(_05198_),
    .C(net359),
    .Y(_05199_));
 INVx1_ASAP7_75t_R _22646_ (.A(_01237_),
    .Y(_05200_));
 NAND2x1_ASAP7_75t_R _22647_ (.A(net338),
    .B(_01235_),
    .Y(_05201_));
 OA211x2_ASAP7_75t_R _22648_ (.A1(net338),
    .A2(_05200_),
    .B(_05201_),
    .C(net308),
    .Y(_05202_));
 OR3x1_ASAP7_75t_R _22649_ (.A(_13132_),
    .B(_05199_),
    .C(_05202_),
    .Y(_05203_));
 INVx1_ASAP7_75t_R _22650_ (.A(_01241_),
    .Y(_05204_));
 NAND2x1_ASAP7_75t_R _22651_ (.A(net338),
    .B(_01239_),
    .Y(_05205_));
 OA211x2_ASAP7_75t_R _22652_ (.A1(net338),
    .A2(_05204_),
    .B(_05205_),
    .C(net308),
    .Y(_05206_));
 INVx1_ASAP7_75t_R _22653_ (.A(_01238_),
    .Y(_05207_));
 NAND2x1_ASAP7_75t_R _22654_ (.A(net313),
    .B(_01240_),
    .Y(_05208_));
 OA211x2_ASAP7_75t_R _22655_ (.A1(net313),
    .A2(_05207_),
    .B(_05208_),
    .C(net359),
    .Y(_05209_));
 OR3x1_ASAP7_75t_R _22656_ (.A(net325),
    .B(_05206_),
    .C(_05209_),
    .Y(_05210_));
 AND3x1_ASAP7_75t_R _22657_ (.A(_13598_),
    .B(_05203_),
    .C(_05210_),
    .Y(_05211_));
 OR3x1_ASAP7_75t_R _22658_ (.A(net315),
    .B(_05196_),
    .C(_05211_),
    .Y(_05212_));
 NAND2x2_ASAP7_75t_R _22659_ (.A(_05181_),
    .B(_05212_),
    .Y(_05213_));
 OA21x2_ASAP7_75t_R _22660_ (.A1(_01740_),
    .A2(_15267_),
    .B(_16207_),
    .Y(_05214_));
 AO21x2_ASAP7_75t_R _22661_ (.A1(_13583_),
    .A2(_05213_),
    .B(_05214_),
    .Y(_05215_));
 BUFx2_ASAP7_75t_R output229 (.A(net229),
    .Y(instr_addr_o[20]));
 INVx1_ASAP7_75t_R _22663_ (.A(_05215_),
    .Y(_18252_));
 INVx1_ASAP7_75t_R _22664_ (.A(_00227_),
    .Y(\cs_registers_i.pc_id_i[29] ));
 INVx1_ASAP7_75t_R _22665_ (.A(_01239_),
    .Y(_05216_));
 NAND2x1_ASAP7_75t_R _22666_ (.A(net371),
    .B(_01235_),
    .Y(_05217_));
 OA211x2_ASAP7_75t_R _22667_ (.A1(net371),
    .A2(_05216_),
    .B(_05217_),
    .C(net306),
    .Y(_05218_));
 NAND2x1_ASAP7_75t_R _22668_ (.A(net371),
    .B(_01234_),
    .Y(_05219_));
 OA211x2_ASAP7_75t_R _22669_ (.A1(net371),
    .A2(_05207_),
    .B(_05219_),
    .C(net410),
    .Y(_05220_));
 OR3x1_ASAP7_75t_R _22670_ (.A(net302),
    .B(_05218_),
    .C(_05220_),
    .Y(_05221_));
 NAND2x1_ASAP7_75t_R _22671_ (.A(net410),
    .B(_01236_),
    .Y(_05222_));
 OA211x2_ASAP7_75t_R _22672_ (.A1(net410),
    .A2(_05200_),
    .B(_05222_),
    .C(net371),
    .Y(_05223_));
 NAND2x1_ASAP7_75t_R _22673_ (.A(net410),
    .B(_01240_),
    .Y(_05224_));
 OA211x2_ASAP7_75t_R _22674_ (.A1(net410),
    .A2(_05204_),
    .B(_05224_),
    .C(_13397_),
    .Y(_05225_));
 OR3x1_ASAP7_75t_R _22675_ (.A(net398),
    .B(_05223_),
    .C(_05225_),
    .Y(_05226_));
 AND3x1_ASAP7_75t_R _22676_ (.A(_13392_),
    .B(_05221_),
    .C(_05226_),
    .Y(_05227_));
 NAND2x1_ASAP7_75t_R _22677_ (.A(net398),
    .B(_01222_),
    .Y(_05228_));
 OA211x2_ASAP7_75t_R _22678_ (.A1(net398),
    .A2(_05176_),
    .B(_05228_),
    .C(_13397_),
    .Y(_05229_));
 NAND2x1_ASAP7_75t_R _22679_ (.A(net398),
    .B(_01218_),
    .Y(_05230_));
 OA211x2_ASAP7_75t_R _22680_ (.A1(net398),
    .A2(_05161_),
    .B(_05230_),
    .C(net371),
    .Y(_05231_));
 OR3x1_ASAP7_75t_R _22681_ (.A(net306),
    .B(_05229_),
    .C(_05231_),
    .Y(_05232_));
 NAND2x1_ASAP7_75t_R _22682_ (.A(net399),
    .B(_01223_),
    .Y(_05233_));
 OA211x2_ASAP7_75t_R _22683_ (.A1(net399),
    .A2(_05173_),
    .B(_05233_),
    .C(_13397_),
    .Y(_05234_));
 NAND2x1_ASAP7_75t_R _22684_ (.A(net399),
    .B(_01219_),
    .Y(_05235_));
 OA211x2_ASAP7_75t_R _22685_ (.A1(net399),
    .A2(_05158_),
    .B(_05235_),
    .C(net371),
    .Y(_05236_));
 OR3x1_ASAP7_75t_R _22686_ (.A(net410),
    .B(_05234_),
    .C(_05236_),
    .Y(_05237_));
 AND3x1_ASAP7_75t_R _22687_ (.A(net364),
    .B(_05232_),
    .C(_05237_),
    .Y(_05238_));
 OR3x2_ASAP7_75t_R _22688_ (.A(net367),
    .B(_05227_),
    .C(_05238_),
    .Y(_05239_));
 NAND2x1_ASAP7_75t_R _22689_ (.A(net399),
    .B(_01215_),
    .Y(_05240_));
 OA211x2_ASAP7_75t_R _22690_ (.A1(net399),
    .A2(_05166_),
    .B(_05240_),
    .C(net306),
    .Y(_05241_));
 NAND2x1_ASAP7_75t_R _22691_ (.A(net399),
    .B(_01214_),
    .Y(_05242_));
 OA211x2_ASAP7_75t_R _22692_ (.A1(net399),
    .A2(_05169_),
    .B(_05242_),
    .C(net410),
    .Y(_05243_));
 INVx1_ASAP7_75t_R _22693_ (.A(_01213_),
    .Y(_05244_));
 NAND2x1_ASAP7_75t_R _22694_ (.A(net399),
    .B(_01680_),
    .Y(_05245_));
 OA211x2_ASAP7_75t_R _22695_ (.A1(net399),
    .A2(_05244_),
    .B(_05245_),
    .C(net306),
    .Y(_05246_));
 NOR2x1_ASAP7_75t_R _22696_ (.A(_01212_),
    .B(_13471_),
    .Y(_05247_));
 OA33x2_ASAP7_75t_R _22697_ (.A1(_13814_),
    .A2(_05241_),
    .A3(_05243_),
    .B1(_05246_),
    .B2(_05247_),
    .B3(_13828_),
    .Y(_05248_));
 NAND2x1_ASAP7_75t_R _22698_ (.A(net397),
    .B(_01227_),
    .Y(_05249_));
 OA211x2_ASAP7_75t_R _22699_ (.A1(net397),
    .A2(_05189_),
    .B(_05249_),
    .C(net306),
    .Y(_05250_));
 NAND2x1_ASAP7_75t_R _22700_ (.A(net397),
    .B(_01226_),
    .Y(_05251_));
 OA211x2_ASAP7_75t_R _22701_ (.A1(net397),
    .A2(_05192_),
    .B(_05251_),
    .C(net410),
    .Y(_05252_));
 OR3x1_ASAP7_75t_R _22702_ (.A(_13397_),
    .B(_05250_),
    .C(_05252_),
    .Y(_05253_));
 NAND2x1_ASAP7_75t_R _22703_ (.A(net397),
    .B(_01231_),
    .Y(_05254_));
 OA211x2_ASAP7_75t_R _22704_ (.A1(net397),
    .A2(_05182_),
    .B(_05254_),
    .C(net306),
    .Y(_05255_));
 NAND2x1_ASAP7_75t_R _22705_ (.A(net397),
    .B(_01230_),
    .Y(_05256_));
 OA211x2_ASAP7_75t_R _22706_ (.A1(net397),
    .A2(_05185_),
    .B(_05256_),
    .C(net410),
    .Y(_05257_));
 OR3x1_ASAP7_75t_R _22707_ (.A(net371),
    .B(_05255_),
    .C(_05257_),
    .Y(_05258_));
 AO21x1_ASAP7_75t_R _22708_ (.A1(_05253_),
    .A2(_05258_),
    .B(_04690_),
    .Y(_05259_));
 OA21x2_ASAP7_75t_R _22709_ (.A1(_13392_),
    .A2(_05248_),
    .B(_05259_),
    .Y(_05260_));
 NAND2x2_ASAP7_75t_R _22710_ (.A(_05239_),
    .B(_05260_),
    .Y(_05261_));
 OA22x2_ASAP7_75t_R _22711_ (.A1(_01612_),
    .A2(_13223_),
    .B1(_13880_),
    .B2(_00227_),
    .Y(_05262_));
 OAI21x1_ASAP7_75t_R _22712_ (.A1(_13782_),
    .A2(_05261_),
    .B(_05262_),
    .Y(_18253_));
 INVx2_ASAP7_75t_R _22713_ (.A(_18253_),
    .Y(_18251_));
 INVx1_ASAP7_75t_R _22714_ (.A(_01253_),
    .Y(_05263_));
 NAND2x1_ASAP7_75t_R _22715_ (.A(net346),
    .B(_01251_),
    .Y(_05264_));
 OA211x2_ASAP7_75t_R _22716_ (.A1(net346),
    .A2(_05263_),
    .B(_05264_),
    .C(net309),
    .Y(_05265_));
 INVx1_ASAP7_75t_R _22717_ (.A(_01252_),
    .Y(_05266_));
 NAND2x1_ASAP7_75t_R _22718_ (.A(net346),
    .B(_01250_),
    .Y(_05267_));
 OA211x2_ASAP7_75t_R _22719_ (.A1(net346),
    .A2(_05266_),
    .B(_05267_),
    .C(net356),
    .Y(_05268_));
 OR3x1_ASAP7_75t_R _22720_ (.A(net317),
    .B(_05265_),
    .C(_05268_),
    .Y(_05269_));
 INVx1_ASAP7_75t_R _22721_ (.A(_01244_),
    .Y(_05270_));
 INVx1_ASAP7_75t_R _22722_ (.A(_01245_),
    .Y(_05271_));
 NAND2x1_ASAP7_75t_R _22723_ (.A(net346),
    .B(_01679_),
    .Y(_05272_));
 OA21x2_ASAP7_75t_R _22724_ (.A1(net346),
    .A2(_05271_),
    .B(_05272_),
    .Y(_05273_));
 AO221x1_ASAP7_75t_R _22725_ (.A1(_05270_),
    .A2(_13190_),
    .B1(_05273_),
    .B2(net309),
    .C(_13598_),
    .Y(_05274_));
 AO21x1_ASAP7_75t_R _22726_ (.A1(_05269_),
    .A2(_05274_),
    .B(_13132_),
    .Y(_05275_));
 INVx1_ASAP7_75t_R _22727_ (.A(_01249_),
    .Y(_05276_));
 NAND2x1_ASAP7_75t_R _22728_ (.A(net346),
    .B(_01247_),
    .Y(_05277_));
 OA211x2_ASAP7_75t_R _22729_ (.A1(net346),
    .A2(_05276_),
    .B(_05277_),
    .C(net309),
    .Y(_05278_));
 INVx1_ASAP7_75t_R _22730_ (.A(_01248_),
    .Y(_05279_));
 NAND2x1_ASAP7_75t_R _22731_ (.A(net346),
    .B(_01246_),
    .Y(_05280_));
 OA211x2_ASAP7_75t_R _22732_ (.A1(net346),
    .A2(_05279_),
    .B(_05280_),
    .C(net355),
    .Y(_05281_));
 OR3x1_ASAP7_75t_R _22733_ (.A(_13598_),
    .B(_05278_),
    .C(_05281_),
    .Y(_05282_));
 INVx1_ASAP7_75t_R _22734_ (.A(_01257_),
    .Y(_05283_));
 NAND2x1_ASAP7_75t_R _22735_ (.A(net346),
    .B(_01255_),
    .Y(_05284_));
 OA211x2_ASAP7_75t_R _22736_ (.A1(net346),
    .A2(_05283_),
    .B(_05284_),
    .C(net310),
    .Y(_05285_));
 INVx1_ASAP7_75t_R _22737_ (.A(_01256_),
    .Y(_05286_));
 NAND2x1_ASAP7_75t_R _22738_ (.A(net346),
    .B(_01254_),
    .Y(_05287_));
 OA211x2_ASAP7_75t_R _22739_ (.A1(net346),
    .A2(_05286_),
    .B(_05287_),
    .C(net356),
    .Y(_05288_));
 OR3x1_ASAP7_75t_R _22740_ (.A(net317),
    .B(_05285_),
    .C(_05288_),
    .Y(_05289_));
 AO21x1_ASAP7_75t_R _22741_ (.A1(_05282_),
    .A2(_05289_),
    .B(net324),
    .Y(_05290_));
 AO21x2_ASAP7_75t_R _22742_ (.A1(_05275_),
    .A2(_05290_),
    .B(_13174_),
    .Y(_05291_));
 INVx1_ASAP7_75t_R _22743_ (.A(_01265_),
    .Y(_05292_));
 NAND2x1_ASAP7_75t_R _22744_ (.A(net345),
    .B(_01263_),
    .Y(_05293_));
 OA211x2_ASAP7_75t_R _22745_ (.A1(net345),
    .A2(_05292_),
    .B(_05293_),
    .C(net310),
    .Y(_05294_));
 INVx1_ASAP7_75t_R _22746_ (.A(_01264_),
    .Y(_05295_));
 NAND2x1_ASAP7_75t_R _22747_ (.A(net345),
    .B(_01262_),
    .Y(_05296_));
 OA211x2_ASAP7_75t_R _22748_ (.A1(net345),
    .A2(_05295_),
    .B(_05296_),
    .C(net355),
    .Y(_05297_));
 OR3x1_ASAP7_75t_R _22749_ (.A(net324),
    .B(_05294_),
    .C(_05297_),
    .Y(_05298_));
 INVx1_ASAP7_75t_R _22750_ (.A(_01261_),
    .Y(_05299_));
 NAND2x1_ASAP7_75t_R _22751_ (.A(net345),
    .B(_01259_),
    .Y(_05300_));
 OA211x2_ASAP7_75t_R _22752_ (.A1(net345),
    .A2(_05299_),
    .B(_05300_),
    .C(net310),
    .Y(_05301_));
 INVx1_ASAP7_75t_R _22753_ (.A(_01260_),
    .Y(_05302_));
 NAND2x1_ASAP7_75t_R _22754_ (.A(net345),
    .B(_01258_),
    .Y(_05303_));
 OA211x2_ASAP7_75t_R _22755_ (.A1(net345),
    .A2(_05302_),
    .B(_05303_),
    .C(net355),
    .Y(_05304_));
 OR3x1_ASAP7_75t_R _22756_ (.A(_13132_),
    .B(_05301_),
    .C(_05304_),
    .Y(_05305_));
 AND3x1_ASAP7_75t_R _22757_ (.A(net317),
    .B(_05298_),
    .C(_05305_),
    .Y(_05306_));
 INVx1_ASAP7_75t_R _22758_ (.A(_01269_),
    .Y(_05307_));
 NAND2x1_ASAP7_75t_R _22759_ (.A(net345),
    .B(_01267_),
    .Y(_05308_));
 OA211x2_ASAP7_75t_R _22760_ (.A1(net345),
    .A2(_05307_),
    .B(_05308_),
    .C(net310),
    .Y(_05309_));
 INVx1_ASAP7_75t_R _22761_ (.A(_01268_),
    .Y(_05310_));
 NAND2x1_ASAP7_75t_R _22762_ (.A(net345),
    .B(_01266_),
    .Y(_05311_));
 OA211x2_ASAP7_75t_R _22763_ (.A1(net344),
    .A2(_05310_),
    .B(_05311_),
    .C(net355),
    .Y(_05312_));
 OR3x1_ASAP7_75t_R _22764_ (.A(_13132_),
    .B(_05309_),
    .C(_05312_),
    .Y(_05313_));
 INVx1_ASAP7_75t_R _22765_ (.A(_01273_),
    .Y(_05314_));
 NAND2x1_ASAP7_75t_R _22766_ (.A(net344),
    .B(_01271_),
    .Y(_05315_));
 OA211x2_ASAP7_75t_R _22767_ (.A1(net344),
    .A2(_05314_),
    .B(_05315_),
    .C(net310),
    .Y(_05316_));
 INVx1_ASAP7_75t_R _22768_ (.A(_01272_),
    .Y(_05317_));
 NAND2x1_ASAP7_75t_R _22769_ (.A(net344),
    .B(_01270_),
    .Y(_05318_));
 OA211x2_ASAP7_75t_R _22770_ (.A1(net344),
    .A2(_05317_),
    .B(_05318_),
    .C(net355),
    .Y(_05319_));
 OR3x1_ASAP7_75t_R _22771_ (.A(net325),
    .B(_05316_),
    .C(_05319_),
    .Y(_05320_));
 AND3x1_ASAP7_75t_R _22772_ (.A(_13598_),
    .B(_05313_),
    .C(_05320_),
    .Y(_05321_));
 OR3x4_ASAP7_75t_R _22773_ (.A(net314),
    .B(_05306_),
    .C(_05321_),
    .Y(_05322_));
 NAND2x2_ASAP7_75t_R _22774_ (.A(_05291_),
    .B(_05322_),
    .Y(_05323_));
 OA21x2_ASAP7_75t_R _22775_ (.A1(_01739_),
    .A2(_15267_),
    .B(_16207_),
    .Y(_05324_));
 AO21x2_ASAP7_75t_R _22776_ (.A1(_13583_),
    .A2(_05323_),
    .B(_05324_),
    .Y(_05325_));
 BUFx2_ASAP7_75t_R output228 (.A(net228),
    .Y(instr_addr_o[19]));
 INVx1_ASAP7_75t_R _22778_ (.A(_05325_),
    .Y(_18257_));
 INVx1_ASAP7_75t_R _22779_ (.A(_01611_),
    .Y(_05326_));
 NAND2x1_ASAP7_75t_R _22780_ (.A(net389),
    .B(_01262_),
    .Y(_05327_));
 OA211x2_ASAP7_75t_R _22781_ (.A1(net389),
    .A2(_05295_),
    .B(_05327_),
    .C(net407),
    .Y(_05328_));
 NAND2x1_ASAP7_75t_R _22782_ (.A(net389),
    .B(_01263_),
    .Y(_05329_));
 OA211x2_ASAP7_75t_R _22783_ (.A1(net389),
    .A2(_05292_),
    .B(_05329_),
    .C(net307),
    .Y(_05330_));
 OR3x1_ASAP7_75t_R _22784_ (.A(_13814_),
    .B(_05328_),
    .C(_05330_),
    .Y(_05331_));
 NAND2x1_ASAP7_75t_R _22785_ (.A(net389),
    .B(_01258_),
    .Y(_05332_));
 OA211x2_ASAP7_75t_R _22786_ (.A1(net389),
    .A2(_05302_),
    .B(_05332_),
    .C(net407),
    .Y(_05333_));
 NAND2x1_ASAP7_75t_R _22787_ (.A(net392),
    .B(_01259_),
    .Y(_05334_));
 OA211x2_ASAP7_75t_R _22788_ (.A1(net392),
    .A2(_05299_),
    .B(_05334_),
    .C(net307),
    .Y(_05335_));
 OR3x1_ASAP7_75t_R _22789_ (.A(net300),
    .B(_05333_),
    .C(_05335_),
    .Y(_05336_));
 NAND2x1_ASAP7_75t_R _22790_ (.A(net392),
    .B(_01247_),
    .Y(_05337_));
 OA211x2_ASAP7_75t_R _22791_ (.A1(net392),
    .A2(_05276_),
    .B(_05337_),
    .C(net307),
    .Y(_05338_));
 NAND2x1_ASAP7_75t_R _22792_ (.A(net392),
    .B(_01246_),
    .Y(_05339_));
 OA211x2_ASAP7_75t_R _22793_ (.A1(net392),
    .A2(_05279_),
    .B(_05339_),
    .C(net407),
    .Y(_05340_));
 OR3x1_ASAP7_75t_R _22794_ (.A(_13814_),
    .B(_05338_),
    .C(_05340_),
    .Y(_05341_));
 NAND2x1_ASAP7_75t_R _22795_ (.A(net392),
    .B(_01679_),
    .Y(_05342_));
 OA211x2_ASAP7_75t_R _22796_ (.A1(net392),
    .A2(_05271_),
    .B(_05342_),
    .C(net306),
    .Y(_05343_));
 AND3x1_ASAP7_75t_R _22797_ (.A(net407),
    .B(net302),
    .C(_05270_),
    .Y(_05344_));
 OA31x2_ASAP7_75t_R _22798_ (.A1(net300),
    .A2(_05343_),
    .A3(_05344_),
    .B1(net362),
    .Y(_05345_));
 AO32x1_ASAP7_75t_R _22799_ (.A1(_13392_),
    .A2(_05331_),
    .A3(_05336_),
    .B1(_05341_),
    .B2(_05345_),
    .Y(_05346_));
 NAND2x1_ASAP7_75t_R _22800_ (.A(net389),
    .B(_01267_),
    .Y(_05347_));
 OA211x2_ASAP7_75t_R _22801_ (.A1(net389),
    .A2(_05307_),
    .B(_05347_),
    .C(net307),
    .Y(_05348_));
 NAND2x1_ASAP7_75t_R _22802_ (.A(net389),
    .B(_01266_),
    .Y(_05349_));
 OA211x2_ASAP7_75t_R _22803_ (.A1(net389),
    .A2(_05310_),
    .B(_05349_),
    .C(net407),
    .Y(_05350_));
 OR3x1_ASAP7_75t_R _22804_ (.A(_13397_),
    .B(_05348_),
    .C(_05350_),
    .Y(_05351_));
 NAND2x1_ASAP7_75t_R _22805_ (.A(net389),
    .B(_01271_),
    .Y(_05352_));
 OA211x2_ASAP7_75t_R _22806_ (.A1(net389),
    .A2(_05314_),
    .B(_05352_),
    .C(net307),
    .Y(_05353_));
 NAND2x1_ASAP7_75t_R _22807_ (.A(net389),
    .B(_01270_),
    .Y(_05354_));
 OA211x2_ASAP7_75t_R _22808_ (.A1(net389),
    .A2(_05317_),
    .B(_05354_),
    .C(net407),
    .Y(_05355_));
 OR3x1_ASAP7_75t_R _22809_ (.A(net370),
    .B(_05353_),
    .C(_05355_),
    .Y(_05356_));
 AND5x1_ASAP7_75t_R _22810_ (.A(_13392_),
    .B(_05331_),
    .C(_05336_),
    .D(_05351_),
    .E(_05356_),
    .Y(_05357_));
 NAND2x1_ASAP7_75t_R _22811_ (.A(net392),
    .B(_01251_),
    .Y(_05358_));
 OA211x2_ASAP7_75t_R _22812_ (.A1(net392),
    .A2(_05263_),
    .B(_05358_),
    .C(net307),
    .Y(_05359_));
 NAND2x1_ASAP7_75t_R _22813_ (.A(net392),
    .B(_01250_),
    .Y(_05360_));
 OA211x2_ASAP7_75t_R _22814_ (.A1(net392),
    .A2(_05266_),
    .B(_05360_),
    .C(net409),
    .Y(_05361_));
 OR3x1_ASAP7_75t_R _22815_ (.A(_13397_),
    .B(_05359_),
    .C(_05361_),
    .Y(_05362_));
 NAND2x1_ASAP7_75t_R _22816_ (.A(net395),
    .B(_01255_),
    .Y(_05363_));
 OA211x2_ASAP7_75t_R _22817_ (.A1(net395),
    .A2(_05283_),
    .B(_05363_),
    .C(net307),
    .Y(_05364_));
 NAND2x1_ASAP7_75t_R _22818_ (.A(net395),
    .B(_01254_),
    .Y(_05365_));
 OA211x2_ASAP7_75t_R _22819_ (.A1(net395),
    .A2(_05286_),
    .B(_05365_),
    .C(net409),
    .Y(_05366_));
 OR3x1_ASAP7_75t_R _22820_ (.A(net373),
    .B(_05364_),
    .C(_05366_),
    .Y(_05367_));
 AND4x1_ASAP7_75t_R _22821_ (.A(_05341_),
    .B(_05345_),
    .C(_05362_),
    .D(_05367_),
    .Y(_05368_));
 AO211x2_ASAP7_75t_R _22822_ (.A1(net366),
    .A2(_05346_),
    .B(_05357_),
    .C(_05368_),
    .Y(_05369_));
 INVx2_ASAP7_75t_R _22823_ (.A(_00229_),
    .Y(_05370_));
 AO222x2_ASAP7_75t_R _22824_ (.A1(_05326_),
    .A2(_13270_),
    .B1(_13563_),
    .B2(_05369_),
    .C1(_14503_),
    .C2(_05370_),
    .Y(_05371_));
 BUFx2_ASAP7_75t_R output227 (.A(net227),
    .Y(instr_addr_o[18]));
 INVx2_ASAP7_75t_R _22826_ (.A(_05371_),
    .Y(_18256_));
 XNOR2x2_ASAP7_75t_R _22827_ (.A(_01277_),
    .B(_01275_),
    .Y(_05372_));
 INVx3_ASAP7_75t_R _22828_ (.A(_05372_),
    .Y(net172));
 INVx1_ASAP7_75t_R _22829_ (.A(_01307_),
    .Y(_05373_));
 NAND2x1_ASAP7_75t_R _22830_ (.A(net348),
    .B(_01305_),
    .Y(_05374_));
 OA211x2_ASAP7_75t_R _22831_ (.A1(net348),
    .A2(_05373_),
    .B(_05374_),
    .C(net310),
    .Y(_05375_));
 INVx1_ASAP7_75t_R _22832_ (.A(_01306_),
    .Y(_05376_));
 NAND2x1_ASAP7_75t_R _22833_ (.A(net348),
    .B(_01304_),
    .Y(_05377_));
 OA211x2_ASAP7_75t_R _22834_ (.A1(net348),
    .A2(_05376_),
    .B(_05377_),
    .C(net361),
    .Y(_05378_));
 OR3x1_ASAP7_75t_R _22835_ (.A(net323),
    .B(_05375_),
    .C(_05378_),
    .Y(_05379_));
 AND2x2_ASAP7_75t_R _22836_ (.A(net347),
    .B(_01300_),
    .Y(_05380_));
 AO21x1_ASAP7_75t_R _22837_ (.A1(net312),
    .A2(_01302_),
    .B(_05380_),
    .Y(_05381_));
 AND2x2_ASAP7_75t_R _22838_ (.A(net347),
    .B(_01301_),
    .Y(_05382_));
 AO21x1_ASAP7_75t_R _22839_ (.A1(net312),
    .A2(_01303_),
    .B(_05382_),
    .Y(_05383_));
 AOI221x1_ASAP7_75t_R _22840_ (.A1(_13184_),
    .A2(_05381_),
    .B1(_05383_),
    .B2(_13164_),
    .C(_13976_),
    .Y(_05384_));
 AND2x2_ASAP7_75t_R _22841_ (.A(net350),
    .B(_01292_),
    .Y(_05385_));
 AO21x1_ASAP7_75t_R _22842_ (.A1(net312),
    .A2(_01294_),
    .B(_05385_),
    .Y(_05386_));
 AND2x2_ASAP7_75t_R _22843_ (.A(net347),
    .B(_01293_),
    .Y(_05387_));
 AO21x1_ASAP7_75t_R _22844_ (.A1(net312),
    .A2(_01295_),
    .B(_05387_),
    .Y(_05388_));
 OA21x2_ASAP7_75t_R _22845_ (.A1(net361),
    .A2(_05388_),
    .B(net323),
    .Y(_05389_));
 OAI21x1_ASAP7_75t_R _22846_ (.A1(net310),
    .A2(_05386_),
    .B(_05389_),
    .Y(_05390_));
 AND2x2_ASAP7_75t_R _22847_ (.A(net348),
    .B(_01297_),
    .Y(_05391_));
 AO21x1_ASAP7_75t_R _22848_ (.A1(net312),
    .A2(_01299_),
    .B(_05391_),
    .Y(_05392_));
 AND2x2_ASAP7_75t_R _22849_ (.A(net348),
    .B(_01296_),
    .Y(_05393_));
 AO21x1_ASAP7_75t_R _22850_ (.A1(net312),
    .A2(_01298_),
    .B(_05393_),
    .Y(_05394_));
 AOI221x1_ASAP7_75t_R _22851_ (.A1(_13124_),
    .A2(_05392_),
    .B1(_05394_),
    .B2(_13133_),
    .C(_13175_),
    .Y(_05395_));
 INVx1_ASAP7_75t_R _22852_ (.A(_01291_),
    .Y(_05396_));
 NAND2x1_ASAP7_75t_R _22853_ (.A(net349),
    .B(_01289_),
    .Y(_05397_));
 OA211x2_ASAP7_75t_R _22854_ (.A1(net349),
    .A2(_05396_),
    .B(_13124_),
    .C(_05397_),
    .Y(_05398_));
 INVx1_ASAP7_75t_R _22855_ (.A(_01290_),
    .Y(_05399_));
 NAND2x1_ASAP7_75t_R _22856_ (.A(net349),
    .B(_01288_),
    .Y(_05400_));
 OA211x2_ASAP7_75t_R _22857_ (.A1(net349),
    .A2(_05399_),
    .B(_13133_),
    .C(_05400_),
    .Y(_05401_));
 INVx1_ASAP7_75t_R _22858_ (.A(_01285_),
    .Y(_05402_));
 NAND2x1_ASAP7_75t_R _22859_ (.A(net312),
    .B(_01287_),
    .Y(_05403_));
 OA211x2_ASAP7_75t_R _22860_ (.A1(net312),
    .A2(_05402_),
    .B(_13164_),
    .C(_05403_),
    .Y(_05404_));
 INVx1_ASAP7_75t_R _22861_ (.A(_01286_),
    .Y(_05405_));
 NAND2x1_ASAP7_75t_R _22862_ (.A(net349),
    .B(_01284_),
    .Y(_05406_));
 OA211x2_ASAP7_75t_R _22863_ (.A1(net349),
    .A2(_05405_),
    .B(_13184_),
    .C(_05406_),
    .Y(_05407_));
 OR5x1_ASAP7_75t_R _22864_ (.A(net317),
    .B(_05398_),
    .C(_05401_),
    .D(_05404_),
    .E(_05407_),
    .Y(_05408_));
 AND2x2_ASAP7_75t_R _22865_ (.A(net349),
    .B(_01678_),
    .Y(_05409_));
 AO21x1_ASAP7_75t_R _22866_ (.A1(net312),
    .A2(_01279_),
    .B(_05409_),
    .Y(_05410_));
 OAI22x1_ASAP7_75t_R _22867_ (.A1(_01278_),
    .A2(_13586_),
    .B1(_05410_),
    .B2(net361),
    .Y(_05411_));
 INVx1_ASAP7_75t_R _22868_ (.A(_01282_),
    .Y(_05412_));
 NAND2x1_ASAP7_75t_R _22869_ (.A(net349),
    .B(_01280_),
    .Y(_05413_));
 OA211x2_ASAP7_75t_R _22870_ (.A1(net349),
    .A2(_05412_),
    .B(_05413_),
    .C(net361),
    .Y(_05414_));
 INVx1_ASAP7_75t_R _22871_ (.A(_01283_),
    .Y(_05415_));
 NAND2x1_ASAP7_75t_R _22872_ (.A(net349),
    .B(_01281_),
    .Y(_05416_));
 OA211x2_ASAP7_75t_R _22873_ (.A1(net349),
    .A2(_05415_),
    .B(_05416_),
    .C(net310),
    .Y(_05417_));
 OR3x1_ASAP7_75t_R _22874_ (.A(_14188_),
    .B(_05414_),
    .C(_05417_),
    .Y(_05418_));
 OA211x2_ASAP7_75t_R _22875_ (.A1(_13584_),
    .A2(_05411_),
    .B(_05418_),
    .C(net314),
    .Y(_05419_));
 AO222x2_ASAP7_75t_R _22876_ (.A1(_05379_),
    .A2(_05384_),
    .B1(_05390_),
    .B2(_05395_),
    .C1(_05408_),
    .C2(_05419_),
    .Y(_05420_));
 AND2x2_ASAP7_75t_R _22877_ (.A(_14597_),
    .B(_13299_),
    .Y(_05421_));
 NAND2x1_ASAP7_75t_R _22878_ (.A(_13298_),
    .B(_14436_),
    .Y(_05422_));
 AOI22x1_ASAP7_75t_R _22879_ (.A1(_13583_),
    .A2(_05420_),
    .B1(_05421_),
    .B2(_05422_),
    .Y(_17586_));
 INVx1_ASAP7_75t_R _22880_ (.A(_17586_),
    .Y(_17588_));
 NAND2x1_ASAP7_75t_R _22881_ (.A(net382),
    .B(_01280_),
    .Y(_05423_));
 OA211x2_ASAP7_75t_R _22882_ (.A1(net382),
    .A2(_05412_),
    .B(_05423_),
    .C(net404),
    .Y(_05424_));
 NAND2x1_ASAP7_75t_R _22883_ (.A(net382),
    .B(_01281_),
    .Y(_05425_));
 OA211x2_ASAP7_75t_R _22884_ (.A1(net382),
    .A2(_05415_),
    .B(_05425_),
    .C(net304),
    .Y(_05426_));
 OR3x1_ASAP7_75t_R _22885_ (.A(net298),
    .B(_05424_),
    .C(_05426_),
    .Y(_05427_));
 INVx1_ASAP7_75t_R _22886_ (.A(_01279_),
    .Y(_05428_));
 NAND2x1_ASAP7_75t_R _22887_ (.A(net404),
    .B(_01278_),
    .Y(_05429_));
 OA211x2_ASAP7_75t_R _22888_ (.A1(net404),
    .A2(_05428_),
    .B(_05429_),
    .C(net302),
    .Y(_05430_));
 INVx1_ASAP7_75t_R _22889_ (.A(_01678_),
    .Y(_05431_));
 AND3x1_ASAP7_75t_R _22890_ (.A(net304),
    .B(net382),
    .C(_05431_),
    .Y(_05432_));
 OR3x1_ASAP7_75t_R _22891_ (.A(net301),
    .B(_05430_),
    .C(_05432_),
    .Y(_05433_));
 AND3x1_ASAP7_75t_R _22892_ (.A(net363),
    .B(_05427_),
    .C(_05433_),
    .Y(_05434_));
 NAND2x1_ASAP7_75t_R _22893_ (.A(net382),
    .B(_01288_),
    .Y(_05435_));
 OA211x2_ASAP7_75t_R _22894_ (.A1(net382),
    .A2(_05399_),
    .B(_05435_),
    .C(_13397_),
    .Y(_05436_));
 NAND2x1_ASAP7_75t_R _22895_ (.A(net382),
    .B(_01284_),
    .Y(_05437_));
 OA211x2_ASAP7_75t_R _22896_ (.A1(net382),
    .A2(_05405_),
    .B(_05437_),
    .C(net369),
    .Y(_05438_));
 OR3x1_ASAP7_75t_R _22897_ (.A(net304),
    .B(_05436_),
    .C(_05438_),
    .Y(_05439_));
 NAND2x1_ASAP7_75t_R _22898_ (.A(net369),
    .B(_01287_),
    .Y(_05440_));
 OA211x2_ASAP7_75t_R _22899_ (.A1(net369),
    .A2(_05396_),
    .B(_05440_),
    .C(net303),
    .Y(_05441_));
 INVx1_ASAP7_75t_R _22900_ (.A(_01289_),
    .Y(_05442_));
 NAND2x1_ASAP7_75t_R _22901_ (.A(net369),
    .B(_01285_),
    .Y(_05443_));
 OA211x2_ASAP7_75t_R _22902_ (.A1(net369),
    .A2(_05442_),
    .B(_05443_),
    .C(net382),
    .Y(_05444_));
 OR3x1_ASAP7_75t_R _22903_ (.A(net404),
    .B(_05441_),
    .C(_05444_),
    .Y(_05445_));
 AO21x1_ASAP7_75t_R _22904_ (.A1(_05439_),
    .A2(_05445_),
    .B(net368),
    .Y(_05446_));
 NAND2x1_ASAP7_75t_R _22905_ (.A(net382),
    .B(_01305_),
    .Y(_05447_));
 OA211x2_ASAP7_75t_R _22906_ (.A1(net382),
    .A2(_05373_),
    .B(_05447_),
    .C(net304),
    .Y(_05448_));
 NAND2x1_ASAP7_75t_R _22907_ (.A(net383),
    .B(_01304_),
    .Y(_05449_));
 OA211x2_ASAP7_75t_R _22908_ (.A1(net383),
    .A2(_05376_),
    .B(_05449_),
    .C(net405),
    .Y(_05450_));
 OR3x1_ASAP7_75t_R _22909_ (.A(net373),
    .B(_05448_),
    .C(_05450_),
    .Y(_05451_));
 AND2x2_ASAP7_75t_R _22910_ (.A(net304),
    .B(net373),
    .Y(_05452_));
 AND2x2_ASAP7_75t_R _22911_ (.A(net383),
    .B(_01301_),
    .Y(_05453_));
 AO21x1_ASAP7_75t_R _22912_ (.A1(net302),
    .A2(_01303_),
    .B(_05453_),
    .Y(_05454_));
 NAND2x1_ASAP7_75t_R _22913_ (.A(_05452_),
    .B(_05454_),
    .Y(_05455_));
 AND2x2_ASAP7_75t_R _22914_ (.A(net405),
    .B(net373),
    .Y(_05456_));
 AND2x2_ASAP7_75t_R _22915_ (.A(net383),
    .B(_01300_),
    .Y(_05457_));
 AO21x1_ASAP7_75t_R _22916_ (.A1(net302),
    .A2(_01302_),
    .B(_05457_),
    .Y(_05458_));
 NAND2x1_ASAP7_75t_R _22917_ (.A(_05456_),
    .B(_05458_),
    .Y(_05459_));
 AND3x1_ASAP7_75t_R _22918_ (.A(_14571_),
    .B(_05455_),
    .C(_05459_),
    .Y(_05460_));
 AND2x2_ASAP7_75t_R _22919_ (.A(net383),
    .B(_01293_),
    .Y(_05461_));
 AO21x1_ASAP7_75t_R _22920_ (.A1(net302),
    .A2(_01295_),
    .B(_05461_),
    .Y(_05462_));
 NOR2x1_ASAP7_75t_R _22921_ (.A(net405),
    .B(net373),
    .Y(_05463_));
 AND2x2_ASAP7_75t_R _22922_ (.A(net382),
    .B(_01297_),
    .Y(_05464_));
 AO21x1_ASAP7_75t_R _22923_ (.A1(net302),
    .A2(_01299_),
    .B(_05464_),
    .Y(_05465_));
 AOI22x1_ASAP7_75t_R _22924_ (.A1(_05462_),
    .A2(_05452_),
    .B1(_05463_),
    .B2(_05465_),
    .Y(_05466_));
 AND2x2_ASAP7_75t_R _22925_ (.A(net382),
    .B(_01296_),
    .Y(_05467_));
 AOI21x1_ASAP7_75t_R _22926_ (.A1(net302),
    .A2(_01298_),
    .B(_05467_),
    .Y(_05468_));
 OR3x1_ASAP7_75t_R _22927_ (.A(net304),
    .B(net369),
    .C(_05468_),
    .Y(_05469_));
 AND2x2_ASAP7_75t_R _22928_ (.A(net383),
    .B(_01292_),
    .Y(_05470_));
 AO21x1_ASAP7_75t_R _22929_ (.A1(net302),
    .A2(_01294_),
    .B(_05470_),
    .Y(_05471_));
 NAND2x1_ASAP7_75t_R _22930_ (.A(_05456_),
    .B(_05471_),
    .Y(_05472_));
 AND4x1_ASAP7_75t_R _22931_ (.A(_04689_),
    .B(_05466_),
    .C(_05469_),
    .D(_05472_),
    .Y(_05473_));
 AO221x2_ASAP7_75t_R _22932_ (.A1(_05434_),
    .A2(_05446_),
    .B1(_05451_),
    .B2(_05460_),
    .C(_05473_),
    .Y(_05474_));
 BUFx2_ASAP7_75t_R output226 (.A(net226),
    .Y(instr_addr_o[17]));
 OAI21x1_ASAP7_75t_R _22934_ (.A1(_01610_),
    .A2(_13223_),
    .B(_13561_),
    .Y(_05476_));
 NAND2x1_ASAP7_75t_R _22935_ (.A(_00230_),
    .B(_13553_),
    .Y(_05477_));
 OA211x2_ASAP7_75t_R _22936_ (.A1(_13782_),
    .A2(_05474_),
    .B(_05476_),
    .C(_05477_),
    .Y(_05478_));
 BUFx2_ASAP7_75t_R output225 (.A(net225),
    .Y(instr_addr_o[16]));
 INVx1_ASAP7_75t_R _22938_ (.A(_05478_),
    .Y(_17587_));
 NAND3x2_ASAP7_75t_R _22939_ (.B(_13387_),
    .C(_17586_),
    .Y(_05479_),
    .A(net294));
 NOR2x1_ASAP7_75t_R _22940_ (.A(_00284_),
    .B(_05474_),
    .Y(_05480_));
 AO22x1_ASAP7_75t_R _22941_ (.A1(_13530_),
    .A2(_01308_),
    .B1(_02202_),
    .B2(_13533_),
    .Y(_05481_));
 OR3x1_ASAP7_75t_R _22942_ (.A(net295),
    .B(_13528_),
    .C(_05481_),
    .Y(_05482_));
 NAND2x1_ASAP7_75t_R _22943_ (.A(_13576_),
    .B(_13528_),
    .Y(_05483_));
 INVx1_ASAP7_75t_R _22944_ (.A(_05420_),
    .Y(_05484_));
 OA222x2_ASAP7_75t_R _22945_ (.A1(_13387_),
    .A2(_17586_),
    .B1(_05480_),
    .B2(_05482_),
    .C1(_05483_),
    .C2(_05484_),
    .Y(_05485_));
 OA21x2_ASAP7_75t_R _22946_ (.A1(_01078_),
    .A2(_01079_),
    .B(_02279_),
    .Y(_05486_));
 OR2x2_ASAP7_75t_R _22947_ (.A(_01143_),
    .B(_01111_),
    .Y(_05487_));
 OA21x2_ASAP7_75t_R _22948_ (.A1(_01143_),
    .A2(_01144_),
    .B(_02280_),
    .Y(_05488_));
 OA21x2_ASAP7_75t_R _22949_ (.A1(_05486_),
    .A2(_05487_),
    .B(_05488_),
    .Y(_05489_));
 OA21x2_ASAP7_75t_R _22950_ (.A1(_01209_),
    .A2(_01210_),
    .B(_02281_),
    .Y(_05490_));
 OA21x2_ASAP7_75t_R _22951_ (.A1(_01243_),
    .A2(_05490_),
    .B(_01276_),
    .Y(_05491_));
 OA21x2_ASAP7_75t_R _22952_ (.A1(_01275_),
    .A2(_05491_),
    .B(_01309_),
    .Y(_05492_));
 AND2x2_ASAP7_75t_R _22953_ (.A(_04608_),
    .B(_05492_),
    .Y(_05493_));
 OR2x2_ASAP7_75t_R _22954_ (.A(_16145_),
    .B(_04605_),
    .Y(_05494_));
 OR3x1_ASAP7_75t_R _22955_ (.A(_01078_),
    .B(_01046_),
    .C(_05487_),
    .Y(_05495_));
 OR4x1_ASAP7_75t_R _22956_ (.A(_01209_),
    .B(_01177_),
    .C(_01275_),
    .D(_01243_),
    .Y(_05496_));
 AO21x1_ASAP7_75t_R _22957_ (.A1(_05489_),
    .A2(_05495_),
    .B(_05496_),
    .Y(_05497_));
 AO32x2_ASAP7_75t_R _22958_ (.A1(_05489_),
    .A2(_05493_),
    .A3(_05494_),
    .B1(_05497_),
    .B2(_05492_),
    .Y(_05498_));
 AND2x2_ASAP7_75t_R _22959_ (.A(_05489_),
    .B(_05495_),
    .Y(_05499_));
 OR4x1_ASAP7_75t_R _22960_ (.A(_16140_),
    .B(_04605_),
    .C(_05496_),
    .D(_05499_),
    .Y(_05500_));
 AO21x2_ASAP7_75t_R _22961_ (.A1(_15413_),
    .A2(_15417_),
    .B(_05500_),
    .Y(_05501_));
 NAND2x2_ASAP7_75t_R _22962_ (.A(_05498_),
    .B(_05501_),
    .Y(_05502_));
 INVx4_ASAP7_75t_R _22963_ (.A(_01308_),
    .Y(_05503_));
 AND3x1_ASAP7_75t_R _22964_ (.A(_05503_),
    .B(_13576_),
    .C(_13533_),
    .Y(_05504_));
 AOI21x1_ASAP7_75t_R _22965_ (.A1(_05498_),
    .A2(_05501_),
    .B(_13576_),
    .Y(_05505_));
 OA21x2_ASAP7_75t_R _22966_ (.A1(_01308_),
    .A2(_13574_),
    .B(_13576_),
    .Y(_05506_));
 AND3x1_ASAP7_75t_R _22967_ (.A(_05498_),
    .B(_05501_),
    .C(_05506_),
    .Y(_05507_));
 AOI221x1_ASAP7_75t_R _22968_ (.A1(_05502_),
    .A2(_05504_),
    .B1(_05505_),
    .B2(_05478_),
    .C(_05507_),
    .Y(_05508_));
 OR3x2_ASAP7_75t_R _22969_ (.A(_13576_),
    .B(_05478_),
    .C(_05502_),
    .Y(_05509_));
 AOI22x1_ASAP7_75t_R _22970_ (.A1(_05479_),
    .A2(_05485_),
    .B1(_05508_),
    .B2(_05509_),
    .Y(_05510_));
 AND4x1_ASAP7_75t_R _22971_ (.A(_05479_),
    .B(_05485_),
    .C(_05508_),
    .D(_05509_),
    .Y(_05511_));
 OR2x6_ASAP7_75t_R _22972_ (.A(_05510_),
    .B(_05511_),
    .Y(_05512_));
 BUFx2_ASAP7_75t_R output224 (.A(net224),
    .Y(instr_addr_o[15]));
 CKINVDCx6p67_ASAP7_75t_R _22974_ (.A(_05512_),
    .Y(net173));
 BUFx2_ASAP7_75t_R output223 (.A(net223),
    .Y(instr_addr_o[14]));
 INVx1_ASAP7_75t_R _22976_ (.A(_02140_),
    .Y(\cs_registers_i.priv_lvl_q[0] ));
 INVx2_ASAP7_75t_R _22977_ (.A(_01314_),
    .Y(_05515_));
 INVx1_ASAP7_75t_R _22978_ (.A(_01874_),
    .Y(_05516_));
 OA21x2_ASAP7_75t_R _22979_ (.A1(_00283_),
    .A2(_13350_),
    .B(_13317_),
    .Y(_05517_));
 AND3x4_ASAP7_75t_R _22980_ (.A(_13313_),
    .B(_13550_),
    .C(_05517_),
    .Y(_05518_));
 NAND2x2_ASAP7_75t_R _22981_ (.A(_05516_),
    .B(_05518_),
    .Y(_05519_));
 NOR2x1_ASAP7_75t_R _22982_ (.A(_14628_),
    .B(_05519_),
    .Y(_05520_));
 AO21x1_ASAP7_75t_R _22983_ (.A1(_05515_),
    .A2(_14628_),
    .B(_05520_),
    .Y(_00001_));
 BUFx2_ASAP7_75t_R output222 (.A(net222),
    .Y(instr_addr_o[13]));
 AND4x2_ASAP7_75t_R _22985_ (.A(_00277_),
    .B(net59),
    .C(_01608_),
    .D(_01609_),
    .Y(_05522_));
 INVx2_ASAP7_75t_R _22986_ (.A(net25),
    .Y(_05523_));
 NAND2x2_ASAP7_75t_R _22987_ (.A(_05523_),
    .B(_01607_),
    .Y(_05524_));
 NAND2x2_ASAP7_75t_R _22988_ (.A(_05522_),
    .B(_05524_),
    .Y(_05525_));
 NOR2x1_ASAP7_75t_R _22989_ (.A(_01316_),
    .B(_05525_),
    .Y(\id_stage_i.controller_i.store_err_d ));
 AND3x1_ASAP7_75t_R _22990_ (.A(_01316_),
    .B(_05522_),
    .C(_05524_),
    .Y(\id_stage_i.controller_i.load_err_d ));
 INVx2_ASAP7_75t_R _22991_ (.A(_01716_),
    .Y(_05526_));
 AND4x2_ASAP7_75t_R _22992_ (.A(_01714_),
    .B(_14581_),
    .C(_05526_),
    .D(_01717_),
    .Y(_05527_));
 BUFx2_ASAP7_75t_R output221 (.A(net221),
    .Y(instr_addr_o[12]));
 BUFx2_ASAP7_75t_R output220 (.A(net220),
    .Y(instr_addr_o[11]));
 BUFx2_ASAP7_75t_R output219 (.A(net219),
    .Y(instr_addr_o[10]));
 OA21x2_ASAP7_75t_R _22996_ (.A1(_13269_),
    .A2(_13653_),
    .B(_13951_),
    .Y(_05531_));
 AO221x1_ASAP7_75t_R _22997_ (.A1(_00283_),
    .A2(_01742_),
    .B1(_13223_),
    .B2(_13248_),
    .C(_13275_),
    .Y(_05532_));
 AO21x1_ASAP7_75t_R _22998_ (.A1(_13298_),
    .A2(_14436_),
    .B(_05532_),
    .Y(_05533_));
 NOR2x2_ASAP7_75t_R _22999_ (.A(_01740_),
    .B(_01741_),
    .Y(_05534_));
 OA211x2_ASAP7_75t_R _23000_ (.A1(_14605_),
    .A2(_14607_),
    .B(_01847_),
    .C(_13567_),
    .Y(_05535_));
 AND3x2_ASAP7_75t_R _23001_ (.A(_01739_),
    .B(_05534_),
    .C(_05535_),
    .Y(_05536_));
 OA21x2_ASAP7_75t_R _23002_ (.A1(_14494_),
    .A2(_14495_),
    .B(_05536_),
    .Y(_05537_));
 AND4x2_ASAP7_75t_R _23003_ (.A(_13299_),
    .B(_05531_),
    .C(_05533_),
    .D(_05537_),
    .Y(_05538_));
 AND3x4_ASAP7_75t_R _23004_ (.A(_14083_),
    .B(_14139_),
    .C(_05538_),
    .Y(_05539_));
 BUFx2_ASAP7_75t_R output218 (.A(net218),
    .Y(data_we_o));
 BUFx2_ASAP7_75t_R output217 (.A(net217),
    .Y(data_wdata_o[9]));
 AND2x6_ASAP7_75t_R _23007_ (.A(_13302_),
    .B(_13658_),
    .Y(_05541_));
 OA21x2_ASAP7_75t_R _23008_ (.A1(_13298_),
    .A2(_14023_),
    .B(_05535_),
    .Y(_05542_));
 BUFx2_ASAP7_75t_R output216 (.A(net216),
    .Y(data_wdata_o[8]));
 AND3x1_ASAP7_75t_R _23010_ (.A(_13954_),
    .B(_05541_),
    .C(_05542_),
    .Y(_05544_));
 BUFx2_ASAP7_75t_R output215 (.A(net215),
    .Y(data_wdata_o[7]));
 BUFx2_ASAP7_75t_R output214 (.A(net214),
    .Y(data_wdata_o[6]));
 BUFx2_ASAP7_75t_R output213 (.A(net213),
    .Y(data_wdata_o[5]));
 INVx2_ASAP7_75t_R _23014_ (.A(_00184_),
    .Y(_05548_));
 CKINVDCx8_ASAP7_75t_R _23015_ (.A(_00385_),
    .Y(_05549_));
 AO33x2_ASAP7_75t_R _23016_ (.A1(_05548_),
    .A2(_13298_),
    .A3(_13952_),
    .B1(_13654_),
    .B2(_13281_),
    .B3(_05549_),
    .Y(_05550_));
 NAND2x1_ASAP7_75t_R _23017_ (.A(_01745_),
    .B(_13648_),
    .Y(_05551_));
 AO32x2_ASAP7_75t_R _23018_ (.A1(_13652_),
    .A2(_13653_),
    .A3(_13654_),
    .B1(_05551_),
    .B2(_13269_),
    .Y(_05552_));
 NOR3x2_ASAP7_75t_R _23019_ (.B(_05550_),
    .C(_05552_),
    .Y(_05553_),
    .A(_13583_));
 AND4x1_ASAP7_75t_R _23020_ (.A(_13955_),
    .B(_14026_),
    .C(_05535_),
    .D(_05553_),
    .Y(_05554_));
 OR3x1_ASAP7_75t_R _23021_ (.A(_13583_),
    .B(_05550_),
    .C(_05552_),
    .Y(_05555_));
 AO21x1_ASAP7_75t_R _23022_ (.A1(_13656_),
    .A2(_05555_),
    .B(_13955_),
    .Y(_05556_));
 AND3x2_ASAP7_75t_R _23023_ (.A(_00279_),
    .B(_00281_),
    .C(_00282_),
    .Y(_05557_));
 OR3x4_ASAP7_75t_R _23024_ (.A(_13547_),
    .B(_05557_),
    .C(_14608_),
    .Y(_05558_));
 BUFx2_ASAP7_75t_R output212 (.A(net212),
    .Y(data_wdata_o[4]));
 OR2x6_ASAP7_75t_R _23026_ (.A(_14024_),
    .B(_05558_),
    .Y(_05560_));
 BUFx2_ASAP7_75t_R output211 (.A(net211),
    .Y(data_wdata_o[3]));
 AO21x1_ASAP7_75t_R _23028_ (.A1(_13656_),
    .A2(_13955_),
    .B(_05560_),
    .Y(_05562_));
 BUFx2_ASAP7_75t_R output210 (.A(net210),
    .Y(data_wdata_o[31]));
 AND3x1_ASAP7_75t_R _23030_ (.A(_13302_),
    .B(_13658_),
    .C(_13954_),
    .Y(_05564_));
 AOI211x1_ASAP7_75t_R _23031_ (.A1(_13301_),
    .A2(_05556_),
    .B(_05562_),
    .C(_05564_),
    .Y(_05565_));
 OR3x1_ASAP7_75t_R _23032_ (.A(_05544_),
    .B(_05554_),
    .C(_05565_),
    .Y(_05566_));
 AND2x2_ASAP7_75t_R _23033_ (.A(_13301_),
    .B(_13656_),
    .Y(_05567_));
 INVx1_ASAP7_75t_R _23034_ (.A(_05567_),
    .Y(_05568_));
 NAND2x1_ASAP7_75t_R _23035_ (.A(_13658_),
    .B(_13954_),
    .Y(_05569_));
 AO22x1_ASAP7_75t_R _23036_ (.A1(_13954_),
    .A2(_05553_),
    .B1(_05568_),
    .B2(_05569_),
    .Y(_05570_));
 AND3x4_ASAP7_75t_R _23037_ (.A(_13306_),
    .B(_14138_),
    .C(_05535_),
    .Y(_05571_));
 AND2x4_ASAP7_75t_R _23038_ (.A(_14084_),
    .B(_05571_),
    .Y(_05572_));
 AND3x1_ASAP7_75t_R _23039_ (.A(_13954_),
    .B(_14026_),
    .C(_05535_),
    .Y(_05573_));
 AO33x2_ASAP7_75t_R _23040_ (.A1(_05542_),
    .A2(_05570_),
    .A3(_05572_),
    .B1(_05573_),
    .B2(_14139_),
    .B3(_05541_),
    .Y(_05574_));
 BUFx2_ASAP7_75t_R output209 (.A(net209),
    .Y(data_wdata_o[30]));
 AND2x4_ASAP7_75t_R _23042_ (.A(_14138_),
    .B(_05537_),
    .Y(_05576_));
 OR4x2_ASAP7_75t_R _23043_ (.A(_14168_),
    .B(_14196_),
    .C(_14226_),
    .D(_14254_),
    .Y(_05577_));
 AOI21x1_ASAP7_75t_R _23044_ (.A1(_13298_),
    .A2(_14436_),
    .B(_05532_),
    .Y(_05578_));
 AOI21x1_ASAP7_75t_R _23045_ (.A1(_13583_),
    .A2(_05577_),
    .B(_05578_),
    .Y(_05579_));
 AND2x2_ASAP7_75t_R _23046_ (.A(_14083_),
    .B(_14139_),
    .Y(_05580_));
 OR5x2_ASAP7_75t_R _23047_ (.A(_13583_),
    .B(_05550_),
    .C(_14024_),
    .D(_14022_),
    .E(_05552_),
    .Y(_05581_));
 OAI21x1_ASAP7_75t_R _23048_ (.A1(_13954_),
    .A2(_05581_),
    .B(_05535_),
    .Y(_05582_));
 BUFx2_ASAP7_75t_R output208 (.A(net208),
    .Y(data_wdata_o[2]));
 AND2x2_ASAP7_75t_R _23050_ (.A(_05580_),
    .B(_05582_),
    .Y(_05584_));
 BUFx2_ASAP7_75t_R output207 (.A(net207),
    .Y(data_wdata_o[29]));
 AND3x4_ASAP7_75t_R _23052_ (.A(_14083_),
    .B(_14140_),
    .C(_05579_),
    .Y(_05586_));
 NOR2x2_ASAP7_75t_R _23053_ (.A(_05558_),
    .B(_05586_),
    .Y(_05587_));
 OR4x2_ASAP7_75t_R _23054_ (.A(_13302_),
    .B(net289),
    .C(_13954_),
    .D(_05560_),
    .Y(_05588_));
 NOR2x1_ASAP7_75t_R _23055_ (.A(_05587_),
    .B(_05588_),
    .Y(_05589_));
 AO21x1_ASAP7_75t_R _23056_ (.A1(_05579_),
    .A2(_05584_),
    .B(_05589_),
    .Y(_05590_));
 AO222x2_ASAP7_75t_R _23057_ (.A1(_05539_),
    .A2(_05566_),
    .B1(_05574_),
    .B2(_05538_),
    .C1(_05576_),
    .C2(_05590_),
    .Y(_05591_));
 AND2x2_ASAP7_75t_R _23058_ (.A(_13954_),
    .B(_14025_),
    .Y(_05592_));
 AND2x2_ASAP7_75t_R _23059_ (.A(_13301_),
    .B(_13658_),
    .Y(_05593_));
 OA211x2_ASAP7_75t_R _23060_ (.A1(_13302_),
    .A2(_05553_),
    .B(_14026_),
    .C(_13955_),
    .Y(_05594_));
 AO21x1_ASAP7_75t_R _23061_ (.A1(_05592_),
    .A2(_05593_),
    .B(_05594_),
    .Y(_05595_));
 AND2x2_ASAP7_75t_R _23062_ (.A(_13955_),
    .B(_14025_),
    .Y(_05596_));
 NAND2x1_ASAP7_75t_R _23063_ (.A(_05535_),
    .B(_05581_),
    .Y(_05597_));
 AO21x1_ASAP7_75t_R _23064_ (.A1(_05541_),
    .A2(_05596_),
    .B(_05597_),
    .Y(_05598_));
 OA21x2_ASAP7_75t_R _23065_ (.A1(_13269_),
    .A2(_13653_),
    .B(_05536_),
    .Y(_05599_));
 OA21x2_ASAP7_75t_R _23066_ (.A1(_14496_),
    .A2(_14491_),
    .B(_05599_),
    .Y(_05600_));
 AND2x2_ASAP7_75t_R _23067_ (.A(_05579_),
    .B(_05600_),
    .Y(_05601_));
 AND4x1_ASAP7_75t_R _23068_ (.A(_14084_),
    .B(_14140_),
    .C(_05535_),
    .D(_05601_),
    .Y(_05602_));
 AO32x1_ASAP7_75t_R _23069_ (.A1(_05538_),
    .A2(_05572_),
    .A3(_05595_),
    .B1(_05598_),
    .B2(_05602_),
    .Y(_05603_));
 NAND2x1_ASAP7_75t_R _23070_ (.A(_13227_),
    .B(_13567_),
    .Y(_05604_));
 NOR2x2_ASAP7_75t_R _23071_ (.A(_14168_),
    .B(_14196_),
    .Y(_05605_));
 AO32x2_ASAP7_75t_R _23072_ (.A1(_00283_),
    .A2(_14199_),
    .A3(_14138_),
    .B1(_05605_),
    .B2(_14255_),
    .Y(_05606_));
 BUFx2_ASAP7_75t_R output206 (.A(net206),
    .Y(data_wdata_o[28]));
 AND5x1_ASAP7_75t_R _23074_ (.A(_14024_),
    .B(_05535_),
    .C(_05576_),
    .D(_05572_),
    .E(_05606_),
    .Y(_05608_));
 AND4x2_ASAP7_75t_R _23075_ (.A(_14084_),
    .B(_14140_),
    .C(_05579_),
    .D(_05535_),
    .Y(_05609_));
 AND3x1_ASAP7_75t_R _23076_ (.A(_13369_),
    .B(_05534_),
    .C(_05535_),
    .Y(_05610_));
 OA211x2_ASAP7_75t_R _23077_ (.A1(_13269_),
    .A2(_13653_),
    .B(_05610_),
    .C(_13951_),
    .Y(_05611_));
 BUFx2_ASAP7_75t_R output205 (.A(net205),
    .Y(data_wdata_o[27]));
 AND3x1_ASAP7_75t_R _23079_ (.A(_18162_),
    .B(_05553_),
    .C(_05611_),
    .Y(_05613_));
 AND4x1_ASAP7_75t_R _23080_ (.A(_13954_),
    .B(_05542_),
    .C(_05609_),
    .D(_05613_),
    .Y(_05614_));
 AND4x1_ASAP7_75t_R _23081_ (.A(_13954_),
    .B(_14026_),
    .C(_14140_),
    .D(_05600_),
    .Y(_05615_));
 NOR2x1_ASAP7_75t_R _23082_ (.A(_14082_),
    .B(_05558_),
    .Y(_05616_));
 AND5x1_ASAP7_75t_R _23083_ (.A(_13955_),
    .B(_14025_),
    .C(_05576_),
    .D(_05571_),
    .E(_05616_),
    .Y(_05617_));
 OA21x2_ASAP7_75t_R _23084_ (.A1(_05615_),
    .A2(_05617_),
    .B(_05606_),
    .Y(_05618_));
 OR4x1_ASAP7_75t_R _23085_ (.A(_05604_),
    .B(_05608_),
    .C(_05614_),
    .D(_05618_),
    .Y(_05619_));
 NAND2x1_ASAP7_75t_R _23086_ (.A(_13955_),
    .B(_14026_),
    .Y(_05620_));
 OAI21x1_ASAP7_75t_R _23087_ (.A1(_14496_),
    .A2(_14491_),
    .B(_05599_),
    .Y(_05621_));
 OR3x1_ASAP7_75t_R _23088_ (.A(_13658_),
    .B(_05620_),
    .C(_05621_),
    .Y(_05622_));
 NOR2x1_ASAP7_75t_R _23089_ (.A(_05587_),
    .B(_05622_),
    .Y(_05623_));
 AO21x1_ASAP7_75t_R _23090_ (.A1(_13955_),
    .A2(_14025_),
    .B(_05558_),
    .Y(_05624_));
 AOI211x1_ASAP7_75t_R _23091_ (.A1(_13306_),
    .A2(_14138_),
    .B(_05558_),
    .C(_14082_),
    .Y(_05625_));
 AND3x2_ASAP7_75t_R _23092_ (.A(_01742_),
    .B(_13299_),
    .C(_14142_),
    .Y(_05626_));
 AND5x2_ASAP7_75t_R _23093_ (.A(_13299_),
    .B(_05531_),
    .C(_05537_),
    .D(_05625_),
    .E(_05626_),
    .Y(_05627_));
 AND2x2_ASAP7_75t_R _23094_ (.A(_05624_),
    .B(_05627_),
    .Y(_05628_));
 AND3x4_ASAP7_75t_R _23095_ (.A(_01742_),
    .B(_14142_),
    .C(_05537_),
    .Y(_05629_));
 AND2x6_ASAP7_75t_R _23096_ (.A(_05625_),
    .B(_05629_),
    .Y(_05630_));
 AO21x1_ASAP7_75t_R _23097_ (.A1(_14083_),
    .A2(_14140_),
    .B(_05558_),
    .Y(_05631_));
 AND2x6_ASAP7_75t_R _23098_ (.A(_05538_),
    .B(_05631_),
    .Y(_05632_));
 AO32x1_ASAP7_75t_R _23099_ (.A1(_05553_),
    .A2(_05592_),
    .A3(_05630_),
    .B1(_05632_),
    .B2(_05597_),
    .Y(_05633_));
 OR5x1_ASAP7_75t_R _23100_ (.A(_05603_),
    .B(_05619_),
    .C(_05623_),
    .D(_05628_),
    .E(_05633_),
    .Y(_05634_));
 NAND2x1_ASAP7_75t_R _23101_ (.A(_14026_),
    .B(_05535_),
    .Y(_05635_));
 AND2x2_ASAP7_75t_R _23102_ (.A(net289),
    .B(_13954_),
    .Y(_05636_));
 OR3x1_ASAP7_75t_R _23103_ (.A(_05635_),
    .B(_05593_),
    .C(_05636_),
    .Y(_05637_));
 AND2x2_ASAP7_75t_R _23104_ (.A(_14026_),
    .B(_05535_),
    .Y(_05638_));
 AO21x1_ASAP7_75t_R _23105_ (.A1(_13955_),
    .A2(_05553_),
    .B(_05564_),
    .Y(_05639_));
 OR3x1_ASAP7_75t_R _23106_ (.A(_05558_),
    .B(_05638_),
    .C(_05639_),
    .Y(_05640_));
 AND4x1_ASAP7_75t_R _23107_ (.A(_05538_),
    .B(_05572_),
    .C(_05637_),
    .D(_05640_),
    .Y(_05641_));
 AND3x1_ASAP7_75t_R _23108_ (.A(_13955_),
    .B(_14026_),
    .C(_05555_),
    .Y(_05642_));
 OAI22x1_ASAP7_75t_R _23109_ (.A1(_13301_),
    .A2(_13656_),
    .B1(_05592_),
    .B2(_05642_),
    .Y(_05643_));
 OR3x1_ASAP7_75t_R _23110_ (.A(_13302_),
    .B(_13658_),
    .C(_14026_),
    .Y(_05644_));
 AND2x2_ASAP7_75t_R _23111_ (.A(_13954_),
    .B(_05560_),
    .Y(_05645_));
 OAI21x1_ASAP7_75t_R _23112_ (.A1(_05596_),
    .A2(_05645_),
    .B(_05541_),
    .Y(_05646_));
 AND5x1_ASAP7_75t_R _23113_ (.A(_05643_),
    .B(_05600_),
    .C(_05609_),
    .D(_05644_),
    .E(_05646_),
    .Y(_05647_));
 AND3x1_ASAP7_75t_R _23114_ (.A(_13954_),
    .B(_05576_),
    .C(_05542_),
    .Y(_05648_));
 OR4x1_ASAP7_75t_R _23115_ (.A(_13954_),
    .B(_14025_),
    .C(_05558_),
    .D(_05621_),
    .Y(_05649_));
 INVx1_ASAP7_75t_R _23116_ (.A(_05649_),
    .Y(_05650_));
 AND3x1_ASAP7_75t_R _23117_ (.A(_05535_),
    .B(_05586_),
    .C(_05593_),
    .Y(_05651_));
 OA21x2_ASAP7_75t_R _23118_ (.A1(_05648_),
    .A2(_05650_),
    .B(_05651_),
    .Y(_05652_));
 NOR2x2_ASAP7_75t_R _23119_ (.A(_14226_),
    .B(_14254_),
    .Y(_05653_));
 AO21x1_ASAP7_75t_R _23120_ (.A1(_13223_),
    .A2(_13248_),
    .B(_01742_),
    .Y(_05654_));
 OA33x2_ASAP7_75t_R _23121_ (.A1(_13299_),
    .A2(_05605_),
    .A3(_05653_),
    .B1(_05654_),
    .B2(_14437_),
    .B3(_00283_),
    .Y(_05655_));
 NAND2x1_ASAP7_75t_R _23122_ (.A(_14497_),
    .B(_05611_),
    .Y(_05656_));
 NOR2x1_ASAP7_75t_R _23123_ (.A(_05655_),
    .B(_05656_),
    .Y(_05657_));
 AND2x2_ASAP7_75t_R _23124_ (.A(_13955_),
    .B(_05542_),
    .Y(_05658_));
 AND4x1_ASAP7_75t_R _23125_ (.A(_13301_),
    .B(_05631_),
    .C(_05657_),
    .D(_05658_),
    .Y(_05659_));
 OR3x1_ASAP7_75t_R _23126_ (.A(_13955_),
    .B(_14025_),
    .C(_05558_),
    .Y(_05660_));
 AND2x2_ASAP7_75t_R _23127_ (.A(_05600_),
    .B(_05606_),
    .Y(_05661_));
 AND5x1_ASAP7_75t_R _23128_ (.A(_13306_),
    .B(_14138_),
    .C(_14497_),
    .D(_05536_),
    .E(_05606_),
    .Y(_05662_));
 AO32x1_ASAP7_75t_R _23129_ (.A1(_14140_),
    .A2(_05660_),
    .A3(_05661_),
    .B1(_05662_),
    .B2(_05542_),
    .Y(_05663_));
 XNOR2x1_ASAP7_75t_R _23130_ (.B(_13656_),
    .Y(_05664_),
    .A(_13302_));
 AND4x1_ASAP7_75t_R _23131_ (.A(_14140_),
    .B(_05592_),
    .C(_05664_),
    .D(_05601_),
    .Y(_05665_));
 AO21x1_ASAP7_75t_R _23132_ (.A1(_14084_),
    .A2(_05663_),
    .B(_05665_),
    .Y(_05666_));
 AND2x2_ASAP7_75t_R _23133_ (.A(_14083_),
    .B(_14140_),
    .Y(_05667_));
 AND2x2_ASAP7_75t_R _23134_ (.A(_05667_),
    .B(_05601_),
    .Y(_05668_));
 AO21x1_ASAP7_75t_R _23135_ (.A1(_13656_),
    .A2(_05596_),
    .B(_05558_),
    .Y(_05669_));
 OR3x1_ASAP7_75t_R _23136_ (.A(_13954_),
    .B(_05560_),
    .C(_05553_),
    .Y(_05670_));
 AND3x1_ASAP7_75t_R _23137_ (.A(_01739_),
    .B(_14138_),
    .C(_05534_),
    .Y(_05671_));
 OA21x2_ASAP7_75t_R _23138_ (.A1(_14394_),
    .A2(_14407_),
    .B(_14433_),
    .Y(_05672_));
 AND4x1_ASAP7_75t_R _23139_ (.A(_13583_),
    .B(_14316_),
    .C(_14373_),
    .D(_05672_),
    .Y(_05673_));
 OA21x2_ASAP7_75t_R _23140_ (.A1(_05671_),
    .A2(_05673_),
    .B(_18162_),
    .Y(_05674_));
 AND4x1_ASAP7_75t_R _23141_ (.A(_05660_),
    .B(_05606_),
    .C(_05625_),
    .D(_05674_),
    .Y(_05675_));
 BUFx2_ASAP7_75t_R output204 (.A(net204),
    .Y(data_wdata_o[26]));
 INVx4_ASAP7_75t_R _23143_ (.A(_01311_),
    .Y(_05677_));
 AO32x1_ASAP7_75t_R _23144_ (.A1(_00283_),
    .A2(_14199_),
    .A3(_13299_),
    .B1(_05605_),
    .B2(_14255_),
    .Y(_05678_));
 AND5x2_ASAP7_75t_R _23145_ (.A(_14084_),
    .B(_14497_),
    .C(_05571_),
    .D(_05611_),
    .E(_05678_),
    .Y(_05679_));
 AND3x1_ASAP7_75t_R _23146_ (.A(_13955_),
    .B(_14026_),
    .C(_05600_),
    .Y(_05680_));
 AO33x2_ASAP7_75t_R _23147_ (.A1(_05677_),
    .A2(_05624_),
    .A3(_05679_),
    .B1(_05680_),
    .B2(_05664_),
    .B3(_05609_),
    .Y(_05681_));
 AO221x1_ASAP7_75t_R _23148_ (.A1(_05668_),
    .A2(_05669_),
    .B1(_05670_),
    .B2(_05675_),
    .C(_05681_),
    .Y(_05682_));
 OR5x1_ASAP7_75t_R _23149_ (.A(_05647_),
    .B(_05652_),
    .C(_05659_),
    .D(_05666_),
    .E(_05682_),
    .Y(_05683_));
 NAND2x2_ASAP7_75t_R _23150_ (.A(_05580_),
    .B(_05538_),
    .Y(_05684_));
 NAND2x1_ASAP7_75t_R _23151_ (.A(net289),
    .B(_13955_),
    .Y(_05685_));
 AOI21x1_ASAP7_75t_R _23152_ (.A1(_05539_),
    .A2(_05685_),
    .B(_13302_),
    .Y(_05686_));
 AOI211x1_ASAP7_75t_R _23153_ (.A1(_05684_),
    .A2(_05569_),
    .B(_05635_),
    .C(_05686_),
    .Y(_05687_));
 OR4x1_ASAP7_75t_R _23154_ (.A(_13301_),
    .B(_13656_),
    .C(_13955_),
    .D(_05602_),
    .Y(_05688_));
 AND4x1_ASAP7_75t_R _23155_ (.A(_13658_),
    .B(_05573_),
    .C(_05667_),
    .D(_05601_),
    .Y(_05689_));
 OA21x2_ASAP7_75t_R _23156_ (.A1(_05675_),
    .A2(_05689_),
    .B(_13302_),
    .Y(_05690_));
 AO21x1_ASAP7_75t_R _23157_ (.A1(_05687_),
    .A2(_05688_),
    .B(_05690_),
    .Y(_05691_));
 XNOR2x1_ASAP7_75t_R _23158_ (.B(_05541_),
    .Y(_05692_),
    .A(_13955_));
 AND3x1_ASAP7_75t_R _23159_ (.A(_05542_),
    .B(_05667_),
    .C(_05601_),
    .Y(_05693_));
 AO21x1_ASAP7_75t_R _23160_ (.A1(_13954_),
    .A2(_05567_),
    .B(_05541_),
    .Y(_05694_));
 AO32x1_ASAP7_75t_R _23161_ (.A1(_05638_),
    .A2(_05668_),
    .A3(_05692_),
    .B1(_05693_),
    .B2(_05694_),
    .Y(_05695_));
 OR5x2_ASAP7_75t_R _23162_ (.A(_05634_),
    .B(_05641_),
    .C(_05683_),
    .D(_05691_),
    .E(_05695_),
    .Y(_05696_));
 OR2x2_ASAP7_75t_R _23163_ (.A(_05591_),
    .B(_05696_),
    .Y(_05697_));
 AND2x2_ASAP7_75t_R _23164_ (.A(_13227_),
    .B(_13567_),
    .Y(_05698_));
 AND3x1_ASAP7_75t_R _23165_ (.A(_02288_),
    .B(_14585_),
    .C(_05535_),
    .Y(_05699_));
 OR2x2_ASAP7_75t_R _23166_ (.A(_01313_),
    .B(_02284_),
    .Y(_05700_));
 INVx1_ASAP7_75t_R _23167_ (.A(_02285_),
    .Y(_05701_));
 OAI21x1_ASAP7_75t_R _23168_ (.A1(_05701_),
    .A2(_02284_),
    .B(_02283_),
    .Y(_05702_));
 AO32x2_ASAP7_75t_R _23169_ (.A1(_18155_),
    .A2(_18162_),
    .A3(_05699_),
    .B1(_05700_),
    .B2(_05702_),
    .Y(_05703_));
 OR5x2_ASAP7_75t_R _23170_ (.A(_01317_),
    .B(_00172_),
    .C(_13245_),
    .D(_13546_),
    .E(_13550_),
    .Y(_05704_));
 OR3x4_ASAP7_75t_R _23171_ (.A(_14600_),
    .B(_14599_),
    .C(_05704_),
    .Y(_05705_));
 BUFx2_ASAP7_75t_R output203 (.A(net203),
    .Y(data_wdata_o[25]));
 BUFx2_ASAP7_75t_R output202 (.A(net202),
    .Y(data_wdata_o[24]));
 NOR2x1_ASAP7_75t_R _23174_ (.A(_17592_),
    .B(_02140_),
    .Y(_05708_));
 NAND2x1_ASAP7_75t_R _23175_ (.A(net309),
    .B(_01745_),
    .Y(_05709_));
 OR4x1_ASAP7_75t_R _23176_ (.A(_14375_),
    .B(_01741_),
    .C(_14188_),
    .D(_05709_),
    .Y(_05710_));
 OR3x2_ASAP7_75t_R _23177_ (.A(_14596_),
    .B(_05704_),
    .C(_05710_),
    .Y(_05711_));
 OR3x4_ASAP7_75t_R _23178_ (.A(_14596_),
    .B(_14600_),
    .C(_05704_),
    .Y(_05712_));
 BUFx2_ASAP7_75t_R output201 (.A(net201),
    .Y(data_wdata_o[23]));
 OA21x2_ASAP7_75t_R _23180_ (.A1(_01997_),
    .A2(_05711_),
    .B(_05712_),
    .Y(_05714_));
 OAI22x1_ASAP7_75t_R _23181_ (.A1(_05677_),
    .A2(_05705_),
    .B1(_05708_),
    .B2(_05714_),
    .Y(_05715_));
 AOI21x1_ASAP7_75t_R _23182_ (.A1(_05698_),
    .A2(_05703_),
    .B(_05715_),
    .Y(_05716_));
 OA211x2_ASAP7_75t_R _23183_ (.A1(_01317_),
    .A2(_14625_),
    .B(_05697_),
    .C(_05716_),
    .Y(_05717_));
 NOR2x1_ASAP7_75t_R _23184_ (.A(_05527_),
    .B(_05717_),
    .Y(\id_stage_i.controller_i.illegal_insn_d ));
 BUFx2_ASAP7_75t_R output200 (.A(net200),
    .Y(data_wdata_o[22]));
 INVx1_ASAP7_75t_R _23186_ (.A(_01721_),
    .Y(_05719_));
 AND3x1_ASAP7_75t_R _23187_ (.A(_00280_),
    .B(_00283_),
    .C(_14595_),
    .Y(_05720_));
 AND4x1_ASAP7_75t_R _23188_ (.A(_01740_),
    .B(_01741_),
    .C(_05557_),
    .D(_13933_),
    .Y(_05721_));
 AND4x1_ASAP7_75t_R _23189_ (.A(_00245_),
    .B(_13772_),
    .C(_05720_),
    .D(_05721_),
    .Y(_05722_));
 NOR2x2_ASAP7_75t_R _23190_ (.A(_05719_),
    .B(_05722_),
    .Y(_05723_));
 AO21x1_ASAP7_75t_R _23191_ (.A1(_14625_),
    .A2(_05723_),
    .B(_01317_),
    .Y(_05724_));
 AND2x2_ASAP7_75t_R _23192_ (.A(_05716_),
    .B(_05724_),
    .Y(_05725_));
 AND2x2_ASAP7_75t_R _23193_ (.A(_05697_),
    .B(_05725_),
    .Y(_05726_));
 NOR2x1_ASAP7_75t_R _23194_ (.A(_05527_),
    .B(_05726_),
    .Y(\id_stage_i.controller_i.exc_req_d ));
 BUFx2_ASAP7_75t_R output199 (.A(net199),
    .Y(data_wdata_o[21]));
 BUFx2_ASAP7_75t_R output198 (.A(net198),
    .Y(data_wdata_o[20]));
 AND2x6_ASAP7_75t_R _23197_ (.A(_14585_),
    .B(_14625_),
    .Y(_05729_));
 AND3x4_ASAP7_75t_R _23198_ (.A(_01713_),
    .B(_14615_),
    .C(_05729_),
    .Y(_05730_));
 NAND2x2_ASAP7_75t_R _23199_ (.A(_01608_),
    .B(_05730_),
    .Y(_05731_));
 NAND2x1_ASAP7_75t_R _23200_ (.A(_00277_),
    .B(net26),
    .Y(_05732_));
 AO21x2_ASAP7_75t_R _23201_ (.A1(_01609_),
    .A2(_05731_),
    .B(_05732_),
    .Y(_05733_));
 INVx2_ASAP7_75t_R _23202_ (.A(_05733_),
    .Y(_05734_));
 OR2x2_ASAP7_75t_R _23203_ (.A(_13273_),
    .B(_13545_),
    .Y(_05735_));
 OR3x1_ASAP7_75t_R _23204_ (.A(_13350_),
    .B(_05735_),
    .C(_05733_),
    .Y(_05736_));
 OAI21x1_ASAP7_75t_R _23205_ (.A1(_01731_),
    .A2(_05734_),
    .B(_05736_),
    .Y(_00007_));
 BUFx2_ASAP7_75t_R output197 (.A(net197),
    .Y(data_wdata_o[1]));
 INVx4_ASAP7_75t_R _23207_ (.A(_01730_),
    .Y(_05738_));
 AND2x2_ASAP7_75t_R _23208_ (.A(_00282_),
    .B(_14615_),
    .Y(_05739_));
 AND3x1_ASAP7_75t_R _23209_ (.A(_00281_),
    .B(_05734_),
    .C(_05739_),
    .Y(_05740_));
 AO21x1_ASAP7_75t_R _23210_ (.A1(_05738_),
    .A2(_05733_),
    .B(_05740_),
    .Y(_00006_));
 INVx2_ASAP7_75t_R _23211_ (.A(_01357_),
    .Y(_05741_));
 BUFx2_ASAP7_75t_R output196 (.A(net196),
    .Y(data_wdata_o[19]));
 AND2x6_ASAP7_75t_R _23213_ (.A(_13325_),
    .B(_13313_),
    .Y(_05743_));
 BUFx2_ASAP7_75t_R output195 (.A(net195),
    .Y(data_wdata_o[18]));
 AND2x6_ASAP7_75t_R _23215_ (.A(_13317_),
    .B(_05743_),
    .Y(_05745_));
 BUFx2_ASAP7_75t_R output194 (.A(net194),
    .Y(data_wdata_o[17]));
 NAND2x2_ASAP7_75t_R _23217_ (.A(_05729_),
    .B(_05745_),
    .Y(_05747_));
 BUFx2_ASAP7_75t_R output193 (.A(net193),
    .Y(data_wdata_o[16]));
 BUFx2_ASAP7_75t_R output192 (.A(net192),
    .Y(data_wdata_o[15]));
 NAND2x2_ASAP7_75t_R _23220_ (.A(_01322_),
    .B(_17607_),
    .Y(_05750_));
 INVx3_ASAP7_75t_R _23221_ (.A(_01318_),
    .Y(_05751_));
 OR2x4_ASAP7_75t_R _23222_ (.A(_01319_),
    .B(_05751_),
    .Y(_05752_));
 OR3x1_ASAP7_75t_R _23223_ (.A(_05747_),
    .B(_05750_),
    .C(_05752_),
    .Y(_05753_));
 BUFx2_ASAP7_75t_R output191 (.A(net191),
    .Y(data_wdata_o[14]));
 NOR2x2_ASAP7_75t_R _23225_ (.A(_01873_),
    .B(_05747_),
    .Y(_05755_));
 BUFx2_ASAP7_75t_R output190 (.A(net190),
    .Y(data_wdata_o[13]));
 AO21x1_ASAP7_75t_R _23227_ (.A1(_05741_),
    .A2(_05753_),
    .B(_05755_),
    .Y(_00005_));
 AND3x4_ASAP7_75t_R _23228_ (.A(_14585_),
    .B(_14625_),
    .C(_05745_),
    .Y(_05757_));
 BUFx2_ASAP7_75t_R output189 (.A(net189),
    .Y(data_wdata_o[12]));
 BUFx2_ASAP7_75t_R output188 (.A(net188),
    .Y(data_wdata_o[11]));
 CKINVDCx8_ASAP7_75t_R _23231_ (.A(net163),
    .Y(_05760_));
 INVx3_ASAP7_75t_R _23232_ (.A(_00676_),
    .Y(net178));
 OR4x1_ASAP7_75t_R _23233_ (.A(net176),
    .B(net180),
    .C(net152),
    .D(_18337_),
    .Y(_05761_));
 OR5x2_ASAP7_75t_R _23234_ (.A(net174),
    .B(net154),
    .C(net158),
    .D(net156),
    .E(_05761_),
    .Y(_05762_));
 OR4x1_ASAP7_75t_R _23235_ (.A(net164),
    .B(net166),
    .C(net168),
    .D(net170),
    .Y(_05763_));
 OR5x1_ASAP7_75t_R _23236_ (.A(net178),
    .B(net257),
    .C(net255),
    .D(_05762_),
    .E(_05763_),
    .Y(_05764_));
 INVx1_ASAP7_75t_R _23237_ (.A(_05764_),
    .Y(_05765_));
 XOR2x2_ASAP7_75t_R _23238_ (.A(_02264_),
    .B(_02223_),
    .Y(_05766_));
 XOR2x2_ASAP7_75t_R _23239_ (.A(_02262_),
    .B(_02222_),
    .Y(_05767_));
 XOR2x2_ASAP7_75t_R _23240_ (.A(_02224_),
    .B(_02266_),
    .Y(_05768_));
 AND5x1_ASAP7_75t_R _23241_ (.A(_05372_),
    .B(_05765_),
    .C(_05766_),
    .D(_05767_),
    .E(_05768_),
    .Y(_05769_));
 XNOR2x2_ASAP7_75t_R _23242_ (.A(_00818_),
    .B(_02275_),
    .Y(_05770_));
 XOR2x2_ASAP7_75t_R _23243_ (.A(_02272_),
    .B(_02226_),
    .Y(_05771_));
 XOR2x2_ASAP7_75t_R _23244_ (.A(_02270_),
    .B(_02225_),
    .Y(_05772_));
 XNOR2x2_ASAP7_75t_R _23245_ (.A(_00679_),
    .B(_02268_),
    .Y(_05773_));
 AND4x1_ASAP7_75t_R _23246_ (.A(_05770_),
    .B(_05771_),
    .C(_05772_),
    .D(_05773_),
    .Y(_05774_));
 AND5x1_ASAP7_75t_R _23247_ (.A(_15557_),
    .B(_16020_),
    .C(_04937_),
    .D(_05154_),
    .E(_05774_),
    .Y(_05775_));
 AND5x2_ASAP7_75t_R _23248_ (.A(_16260_),
    .B(_05760_),
    .C(_04719_),
    .D(_05769_),
    .E(_05775_),
    .Y(_05776_));
 OA21x2_ASAP7_75t_R _23249_ (.A1(_05510_),
    .A2(_05511_),
    .B(_05776_),
    .Y(_05777_));
 INVx2_ASAP7_75t_R _23250_ (.A(_01872_),
    .Y(_05778_));
 NAND2x1_ASAP7_75t_R _23251_ (.A(_05778_),
    .B(_05757_),
    .Y(_05779_));
 OAI22x1_ASAP7_75t_R _23252_ (.A1(_00284_),
    .A2(_05757_),
    .B1(_05777_),
    .B2(_05779_),
    .Y(_00004_));
 BUFx2_ASAP7_75t_R output187 (.A(net187),
    .Y(data_wdata_o[10]));
 AO21x1_ASAP7_75t_R _23254_ (.A1(_05778_),
    .A2(_05777_),
    .B(_13530_),
    .Y(_05781_));
 NAND2x1_ASAP7_75t_R _23255_ (.A(_01728_),
    .B(_05747_),
    .Y(_05782_));
 OA21x2_ASAP7_75t_R _23256_ (.A1(_05747_),
    .A2(_05781_),
    .B(_05782_),
    .Y(_00003_));
 BUFx2_ASAP7_75t_R output186 (.A(net186),
    .Y(data_wdata_o[0]));
 BUFx2_ASAP7_75t_R output185 (.A(net185),
    .Y(data_req_o));
 BUFx2_ASAP7_75t_R output184 (.A(net184),
    .Y(data_be_o[3]));
 OR4x1_ASAP7_75t_R _23260_ (.A(_01357_),
    .B(_05747_),
    .C(_05750_),
    .D(_05752_),
    .Y(_05786_));
 OAI21x1_ASAP7_75t_R _23261_ (.A1(_01727_),
    .A2(_05757_),
    .B(_05786_),
    .Y(_00002_));
 INVx3_ASAP7_75t_R _23262_ (.A(_05767_),
    .Y(net171));
 INVx4_ASAP7_75t_R _23263_ (.A(_05766_),
    .Y(net175));
 INVx3_ASAP7_75t_R _23264_ (.A(_05768_),
    .Y(net177));
 INVx3_ASAP7_75t_R _23265_ (.A(_05773_),
    .Y(net179));
 INVx2_ASAP7_75t_R _23266_ (.A(_05772_),
    .Y(net151));
 INVx3_ASAP7_75t_R _23267_ (.A(_05771_),
    .Y(net153));
 INVx2_ASAP7_75t_R _23268_ (.A(_05770_),
    .Y(net157));
 AND3x4_ASAP7_75t_R _23269_ (.A(_13238_),
    .B(_14615_),
    .C(_14625_),
    .Y(net218));
 INVx4_ASAP7_75t_R _23270_ (.A(_17600_),
    .Y(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ));
 INVx1_ASAP7_75t_R _23271_ (.A(_02291_),
    .Y(_17603_));
 INVx2_ASAP7_75t_R _23272_ (.A(net280),
    .Y(_16503_));
 INVx8_ASAP7_75t_R _23273_ (.A(net279),
    .Y(_16499_));
 BUFx2_ASAP7_75t_R output183 (.A(net183),
    .Y(data_be_o[2]));
 AND2x6_ASAP7_75t_R _23275_ (.A(_01314_),
    .B(_01875_),
    .Y(_05788_));
 BUFx2_ASAP7_75t_R output182 (.A(net182),
    .Y(data_be_o[1]));
 OR2x2_ASAP7_75t_R _23277_ (.A(_01874_),
    .B(_05518_),
    .Y(_05790_));
 AND2x6_ASAP7_75t_R _23278_ (.A(_05788_),
    .B(_05790_),
    .Y(_05791_));
 BUFx2_ASAP7_75t_R output181 (.A(net181),
    .Y(data_be_o[0]));
 BUFx2_ASAP7_75t_R output180 (.A(net180),
    .Y(data_addr_o[9]));
 OAI22x1_ASAP7_75t_R _23281_ (.A1(_00324_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_00816_),
    .Y(_17608_));
 NAND2x2_ASAP7_75t_R _23282_ (.A(_01314_),
    .B(_01875_),
    .Y(_05794_));
 AND3x1_ASAP7_75t_R _23283_ (.A(_15699_),
    .B(_15730_),
    .C(_05794_),
    .Y(_05795_));
 AO21x2_ASAP7_75t_R _23284_ (.A1(_13640_),
    .A2(_05788_),
    .B(_05795_),
    .Y(_05796_));
 BUFx2_ASAP7_75t_R output179 (.A(net179),
    .Y(data_addr_o[8]));
 AND2x6_ASAP7_75t_R _23286_ (.A(_01314_),
    .B(_01874_),
    .Y(_05798_));
 BUFx2_ASAP7_75t_R output178 (.A(net178),
    .Y(data_addr_o[7]));
 NAND2x2_ASAP7_75t_R _23288_ (.A(_01314_),
    .B(_01874_),
    .Y(_05800_));
 BUFx2_ASAP7_75t_R output177 (.A(net177),
    .Y(data_addr_o[6]));
 AND3x1_ASAP7_75t_R _23290_ (.A(_15754_),
    .B(_15777_),
    .C(_05800_),
    .Y(_05802_));
 AO21x2_ASAP7_75t_R _23291_ (.A1(_13758_),
    .A2(_05798_),
    .B(_05802_),
    .Y(_05803_));
 BUFx2_ASAP7_75t_R output176 (.A(net176),
    .Y(data_addr_o[5]));
 AND2x2_ASAP7_75t_R _23293_ (.A(_05796_),
    .B(_05803_),
    .Y(_17609_));
 OAI22x1_ASAP7_75t_R _23294_ (.A1(_00291_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_00849_),
    .Y(_17615_));
 BUFx2_ASAP7_75t_R output175 (.A(net175),
    .Y(data_addr_o[4]));
 OAI22x1_ASAP7_75t_R _23296_ (.A1(_00663_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_00881_),
    .Y(_17622_));
 AND3x1_ASAP7_75t_R _23297_ (.A(_15935_),
    .B(_15970_),
    .C(_05794_),
    .Y(_05806_));
 AO21x2_ASAP7_75t_R _23298_ (.A1(_13943_),
    .A2(_05788_),
    .B(_05806_),
    .Y(_05807_));
 BUFx2_ASAP7_75t_R output174 (.A(net275),
    .Y(data_addr_o[3]));
 BUFx2_ASAP7_75t_R output173 (.A(net173),
    .Y(data_addr_o[31]));
 NAND2x1_ASAP7_75t_R _23301_ (.A(_05803_),
    .B(_05807_),
    .Y(_16546_));
 OAI22x1_ASAP7_75t_R _23302_ (.A1(_00665_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_00914_),
    .Y(_17626_));
 BUFx2_ASAP7_75t_R output172 (.A(net172),
    .Y(data_addr_o[30]));
 AND3x1_ASAP7_75t_R _23304_ (.A(_16050_),
    .B(_16082_),
    .C(_05794_),
    .Y(_05811_));
 AO21x2_ASAP7_75t_R _23305_ (.A1(_14019_),
    .A2(_05788_),
    .B(_05811_),
    .Y(_05812_));
 BUFx2_ASAP7_75t_R output171 (.A(net171),
    .Y(data_addr_o[2]));
 AND2x2_ASAP7_75t_R _23307_ (.A(_05803_),
    .B(_05812_),
    .Y(_17627_));
 OR2x2_ASAP7_75t_R _23308_ (.A(_15890_),
    .B(_05798_),
    .Y(_05814_));
 OA21x2_ASAP7_75t_R _23309_ (.A1(_13523_),
    .A2(_05800_),
    .B(_05814_),
    .Y(_05815_));
 BUFx2_ASAP7_75t_R output170 (.A(net2117),
    .Y(data_addr_o[29]));
 NAND2x1_ASAP7_75t_R _23311_ (.A(_05807_),
    .B(_05815_),
    .Y(_16549_));
 BUFx2_ASAP7_75t_R output169 (.A(net169),
    .Y(data_addr_o[28]));
 OAI22x1_ASAP7_75t_R _23313_ (.A1(_00668_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_00946_),
    .Y(_17641_));
 AND3x1_ASAP7_75t_R _23314_ (.A(_15994_),
    .B(_16017_),
    .C(_05800_),
    .Y(_05818_));
 AO21x2_ASAP7_75t_R _23315_ (.A1(_14684_),
    .A2(_05798_),
    .B(_05818_),
    .Y(_05819_));
 BUFx2_ASAP7_75t_R output168 (.A(net168),
    .Y(data_addr_o[27]));
 NAND2x1_ASAP7_75t_R _23317_ (.A(_05807_),
    .B(_05819_),
    .Y(_16556_));
 OAI22x1_ASAP7_75t_R _23318_ (.A1(_00670_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_00979_),
    .Y(_17651_));
 AND3x1_ASAP7_75t_R _23319_ (.A(_16292_),
    .B(_16323_),
    .C(_05794_),
    .Y(_05821_));
 AO21x2_ASAP7_75t_R _23320_ (.A1(_14137_),
    .A2(_05788_),
    .B(_05821_),
    .Y(_05822_));
 BUFx2_ASAP7_75t_R output167 (.A(net167),
    .Y(data_addr_o[26]));
 AND2x2_ASAP7_75t_R _23322_ (.A(_05803_),
    .B(_05822_),
    .Y(_16566_));
 AND2x2_ASAP7_75t_R _23323_ (.A(_14080_),
    .B(_05788_),
    .Y(_05824_));
 AO21x2_ASAP7_75t_R _23324_ (.A1(_16204_),
    .A2(_05794_),
    .B(_05824_),
    .Y(_05825_));
 BUFx2_ASAP7_75t_R output166 (.A(net166),
    .Y(data_addr_o[25]));
 AND2x2_ASAP7_75t_R _23326_ (.A(_05815_),
    .B(_05825_),
    .Y(_16567_));
 AND2x2_ASAP7_75t_R _23327_ (.A(_05812_),
    .B(_05819_),
    .Y(_16568_));
 OR2x2_ASAP7_75t_R _23328_ (.A(_14752_),
    .B(_05800_),
    .Y(_05827_));
 OA21x2_ASAP7_75t_R _23329_ (.A1(_16132_),
    .A2(_05798_),
    .B(_05827_),
    .Y(_05828_));
 BUFx2_ASAP7_75t_R output165 (.A(net165),
    .Y(data_addr_o[24]));
 NAND2x1_ASAP7_75t_R _23331_ (.A(_05807_),
    .B(_05828_),
    .Y(_16570_));
 BUFx2_ASAP7_75t_R output164 (.A(net164),
    .Y(data_addr_o[23]));
 OAI22x1_ASAP7_75t_R _23333_ (.A1(_00672_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_01011_),
    .Y(_17657_));
 AND3x1_ASAP7_75t_R _23334_ (.A(_16399_),
    .B(_16432_),
    .C(_05794_),
    .Y(_05831_));
 AO21x2_ASAP7_75t_R _23335_ (.A1(_14197_),
    .A2(_05788_),
    .B(_05831_),
    .Y(_05832_));
 BUFx2_ASAP7_75t_R output163 (.A(net163),
    .Y(data_addr_o[22]));
 AND2x2_ASAP7_75t_R _23337_ (.A(_05803_),
    .B(_05832_),
    .Y(_17654_));
 AND2x2_ASAP7_75t_R _23338_ (.A(_05815_),
    .B(_05822_),
    .Y(_16587_));
 AND2x2_ASAP7_75t_R _23339_ (.A(_05819_),
    .B(_05825_),
    .Y(_16588_));
 AND2x2_ASAP7_75t_R _23340_ (.A(_05812_),
    .B(_05828_),
    .Y(_16589_));
 AND3x1_ASAP7_75t_R _23341_ (.A(_16230_),
    .B(_16255_),
    .C(_05800_),
    .Y(_05834_));
 AO21x2_ASAP7_75t_R _23342_ (.A1(_14820_),
    .A2(_05798_),
    .B(_05834_),
    .Y(_05835_));
 BUFx2_ASAP7_75t_R output162 (.A(net255),
    .Y(data_addr_o[21]));
 NAND2x1_ASAP7_75t_R _23344_ (.A(_05807_),
    .B(_05835_),
    .Y(_16591_));
 BUFx2_ASAP7_75t_R output161 (.A(net161),
    .Y(data_addr_o[20]));
 OAI22x1_ASAP7_75t_R _23346_ (.A1(_00674_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_01045_),
    .Y(_17669_));
 OR2x4_ASAP7_75t_R _23347_ (.A(_14226_),
    .B(_14254_),
    .Y(_05838_));
 AND2x2_ASAP7_75t_R _23348_ (.A(_05838_),
    .B(_05788_),
    .Y(_05839_));
 AO21x2_ASAP7_75t_R _23349_ (.A1(_04547_),
    .A2(_05794_),
    .B(_05839_),
    .Y(_05840_));
 BUFx2_ASAP7_75t_R output160 (.A(net160),
    .Y(data_addr_o[19]));
 AND2x2_ASAP7_75t_R _23351_ (.A(_05803_),
    .B(_05840_),
    .Y(_17663_));
 AND2x2_ASAP7_75t_R _23352_ (.A(_05815_),
    .B(_05832_),
    .Y(_17664_));
 AND2x2_ASAP7_75t_R _23353_ (.A(_05819_),
    .B(_05822_),
    .Y(_16606_));
 AND2x2_ASAP7_75t_R _23354_ (.A(_05825_),
    .B(_05828_),
    .Y(_16607_));
 AND2x2_ASAP7_75t_R _23355_ (.A(_05812_),
    .B(_05835_),
    .Y(_16608_));
 OR2x2_ASAP7_75t_R _23356_ (.A(_14873_),
    .B(_05800_),
    .Y(_05842_));
 OA21x2_ASAP7_75t_R _23357_ (.A1(_16372_),
    .A2(_05798_),
    .B(_05842_),
    .Y(_05843_));
 BUFx2_ASAP7_75t_R output159 (.A(net159),
    .Y(data_addr_o[18]));
 NAND2x1_ASAP7_75t_R _23359_ (.A(_05807_),
    .B(_05843_),
    .Y(_16610_));
 OAI22x1_ASAP7_75t_R _23360_ (.A1(_00677_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_01077_),
    .Y(_17676_));
 AND3x1_ASAP7_75t_R _23361_ (.A(_04635_),
    .B(_04666_),
    .C(_05794_),
    .Y(_05845_));
 AO21x2_ASAP7_75t_R _23362_ (.A1(_14316_),
    .A2(_05788_),
    .B(_05845_),
    .Y(_05846_));
 BUFx2_ASAP7_75t_R output158 (.A(net158),
    .Y(data_addr_o[17]));
 BUFx2_ASAP7_75t_R output157 (.A(net157),
    .Y(data_addr_o[16]));
 NAND2x1_ASAP7_75t_R _23365_ (.A(_05803_),
    .B(_05846_),
    .Y(_16624_));
 AND2x2_ASAP7_75t_R _23366_ (.A(_05822_),
    .B(_05828_),
    .Y(_16628_));
 AND2x2_ASAP7_75t_R _23367_ (.A(_05825_),
    .B(_05835_),
    .Y(_16629_));
 AND2x2_ASAP7_75t_R _23368_ (.A(_05812_),
    .B(_05843_),
    .Y(_16630_));
 AO22x2_ASAP7_75t_R _23369_ (.A1(_16446_),
    .A2(_16455_),
    .B1(_16466_),
    .B2(_16477_),
    .Y(_05849_));
 OR2x2_ASAP7_75t_R _23370_ (.A(_05849_),
    .B(_05798_),
    .Y(_05850_));
 OA21x2_ASAP7_75t_R _23371_ (.A1(_14936_),
    .A2(_05800_),
    .B(_05850_),
    .Y(_05851_));
 BUFx2_ASAP7_75t_R output156 (.A(net156),
    .Y(data_addr_o[15]));
 NAND2x1_ASAP7_75t_R _23373_ (.A(_05807_),
    .B(_05851_),
    .Y(_16636_));
 OAI22x1_ASAP7_75t_R _23374_ (.A1(_00680_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_01110_),
    .Y(_17681_));
 INVx2_ASAP7_75t_R _23375_ (.A(_04780_),
    .Y(_05853_));
 AND2x2_ASAP7_75t_R _23376_ (.A(_14373_),
    .B(_05788_),
    .Y(_05854_));
 AO21x2_ASAP7_75t_R _23377_ (.A1(_05853_),
    .A2(_05794_),
    .B(_05854_),
    .Y(_05855_));
 BUFx2_ASAP7_75t_R output155 (.A(net155),
    .Y(data_addr_o[14]));
 AND2x2_ASAP7_75t_R _23379_ (.A(_05803_),
    .B(_05855_),
    .Y(_17682_));
 NAND2x1_ASAP7_75t_R _23380_ (.A(_05815_),
    .B(_05846_),
    .Y(_16654_));
 AND2x2_ASAP7_75t_R _23381_ (.A(_05822_),
    .B(_05835_),
    .Y(_16659_));
 AND2x2_ASAP7_75t_R _23382_ (.A(_05825_),
    .B(_05843_),
    .Y(_16660_));
 AND2x2_ASAP7_75t_R _23383_ (.A(_05812_),
    .B(_05851_),
    .Y(_16661_));
 AND3x1_ASAP7_75t_R _23384_ (.A(_14961_),
    .B(_14989_),
    .C(_05798_),
    .Y(_05857_));
 AO21x2_ASAP7_75t_R _23385_ (.A1(_04595_),
    .A2(_05800_),
    .B(_05857_),
    .Y(_05858_));
 BUFx2_ASAP7_75t_R output154 (.A(net154),
    .Y(data_addr_o[13]));
 NAND2x1_ASAP7_75t_R _23387_ (.A(_05807_),
    .B(_05858_),
    .Y(_16663_));
 BUFx2_ASAP7_75t_R output153 (.A(net153),
    .Y(data_addr_o[12]));
 BUFx2_ASAP7_75t_R output152 (.A(net152),
    .Y(data_addr_o[11]));
 OAI22x1_ASAP7_75t_R _23390_ (.A1(_00682_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_01142_),
    .Y(_17698_));
 NAND2x1_ASAP7_75t_R _23391_ (.A(_05819_),
    .B(_05846_),
    .Y(_16678_));
 AND2x2_ASAP7_75t_R _23392_ (.A(_05822_),
    .B(_05843_),
    .Y(_16683_));
 AND2x2_ASAP7_75t_R _23393_ (.A(_05825_),
    .B(_05851_),
    .Y(_16684_));
 AND2x2_ASAP7_75t_R _23394_ (.A(_05812_),
    .B(_05858_),
    .Y(_16685_));
 AND2x2_ASAP7_75t_R _23395_ (.A(_15042_),
    .B(_05798_),
    .Y(_05862_));
 AO21x2_ASAP7_75t_R _23396_ (.A1(_04715_),
    .A2(_05800_),
    .B(_05862_),
    .Y(_05863_));
 BUFx2_ASAP7_75t_R output151 (.A(net151),
    .Y(data_addr_o[10]));
 BUFx2_ASAP7_75t_R output150 (.A(net150),
    .Y(core_sleep_o));
 NAND2x1_ASAP7_75t_R _23399_ (.A(_05807_),
    .B(_05863_),
    .Y(_16691_));
 OAI22x1_ASAP7_75t_R _23400_ (.A1(_00684_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_01176_),
    .Y(_17710_));
 AND3x1_ASAP7_75t_R _23401_ (.A(_04964_),
    .B(_04995_),
    .C(_05794_),
    .Y(_05866_));
 AO21x2_ASAP7_75t_R _23402_ (.A1(_14489_),
    .A2(_05788_),
    .B(_05866_),
    .Y(_05867_));
 BUFx2_ASAP7_75t_R input149 (.A(test_en_i),
    .Y(net149));
 BUFx16f_ASAP7_75t_R input148 (.A(rst_ni),
    .Y(net148));
 NAND2x1_ASAP7_75t_R _23405_ (.A(_05803_),
    .B(_05867_),
    .Y(_16708_));
 NAND2x1_ASAP7_75t_R _23406_ (.A(_05828_),
    .B(_05846_),
    .Y(_16711_));
 AND2x2_ASAP7_75t_R _23407_ (.A(_05822_),
    .B(_05851_),
    .Y(_16716_));
 AND2x2_ASAP7_75t_R _23408_ (.A(_05825_),
    .B(_05858_),
    .Y(_16717_));
 AND2x2_ASAP7_75t_R _23409_ (.A(_05812_),
    .B(_05863_),
    .Y(_16718_));
 OR2x2_ASAP7_75t_R _23410_ (.A(_15096_),
    .B(_05800_),
    .Y(_05870_));
 OA21x2_ASAP7_75t_R _23411_ (.A1(_04828_),
    .A2(_05798_),
    .B(_05870_),
    .Y(_05871_));
 BUFx2_ASAP7_75t_R input147 (.A(irq_timer_i),
    .Y(net147));
 BUFx2_ASAP7_75t_R input146 (.A(irq_software_i),
    .Y(net146));
 NAND2x1_ASAP7_75t_R _23414_ (.A(_05807_),
    .B(_05871_),
    .Y(_16724_));
 OAI22x1_ASAP7_75t_R _23415_ (.A1(_00686_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_01208_),
    .Y(_17724_));
 OR2x2_ASAP7_75t_R _23416_ (.A(_15266_),
    .B(_05794_),
    .Y(_05874_));
 OAI21x1_ASAP7_75t_R _23417_ (.A1(_05105_),
    .A2(_05788_),
    .B(_05874_),
    .Y(_05875_));
 BUFx3_ASAP7_75t_R input145 (.A(irq_nm_i),
    .Y(net145));
 AND2x2_ASAP7_75t_R _23419_ (.A(_05803_),
    .B(_05875_),
    .Y(_17725_));
 NAND2x1_ASAP7_75t_R _23420_ (.A(_05815_),
    .B(_05867_),
    .Y(_16740_));
 NAND2x1_ASAP7_75t_R _23421_ (.A(_05835_),
    .B(_05846_),
    .Y(_16743_));
 AND2x2_ASAP7_75t_R _23422_ (.A(_05822_),
    .B(_05858_),
    .Y(_16748_));
 AND2x2_ASAP7_75t_R _23423_ (.A(_05825_),
    .B(_05863_),
    .Y(_16749_));
 AND2x2_ASAP7_75t_R _23424_ (.A(_05812_),
    .B(_05871_),
    .Y(_16750_));
 AND3x1_ASAP7_75t_R _23425_ (.A(_04910_),
    .B(_04934_),
    .C(_05800_),
    .Y(_05877_));
 AO21x2_ASAP7_75t_R _23426_ (.A1(_15157_),
    .A2(_05798_),
    .B(_05877_),
    .Y(_05878_));
 BUFx2_ASAP7_75t_R input144 (.A(irq_fast_i[9]),
    .Y(net144));
 BUFx2_ASAP7_75t_R input143 (.A(irq_fast_i[8]),
    .Y(net143));
 NAND2x1_ASAP7_75t_R _23429_ (.A(_05807_),
    .B(_05878_),
    .Y(_16758_));
 BUFx2_ASAP7_75t_R input142 (.A(irq_fast_i[7]),
    .Y(net142));
 OAI22x1_ASAP7_75t_R _23431_ (.A1(_00718_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_01242_),
    .Y(_17745_));
 NAND2x1_ASAP7_75t_R _23432_ (.A(_05819_),
    .B(_05867_),
    .Y(_16777_));
 NAND2x1_ASAP7_75t_R _23433_ (.A(_05843_),
    .B(_05846_),
    .Y(_16785_));
 AND2x2_ASAP7_75t_R _23434_ (.A(_05822_),
    .B(_05863_),
    .Y(_16790_));
 AND2x2_ASAP7_75t_R _23435_ (.A(_05825_),
    .B(_05871_),
    .Y(_16791_));
 AND2x2_ASAP7_75t_R _23436_ (.A(_05812_),
    .B(_05878_),
    .Y(_16789_));
 AND3x1_ASAP7_75t_R _23437_ (.A(_05020_),
    .B(_05043_),
    .C(_05800_),
    .Y(_05882_));
 AO21x2_ASAP7_75t_R _23438_ (.A1(_14574_),
    .A2(_05798_),
    .B(_05882_),
    .Y(_05883_));
 BUFx2_ASAP7_75t_R input141 (.A(irq_fast_i[6]),
    .Y(net141));
 BUFx2_ASAP7_75t_R input140 (.A(irq_fast_i[5]),
    .Y(net140));
 NAND2x1_ASAP7_75t_R _23441_ (.A(_05807_),
    .B(_05883_),
    .Y(_16799_));
 BUFx2_ASAP7_75t_R input139 (.A(irq_fast_i[4]),
    .Y(net139));
 OAI22x1_ASAP7_75t_R _23443_ (.A1(_00750_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_01274_),
    .Y(_17761_));
 INVx2_ASAP7_75t_R _23444_ (.A(_15507_),
    .Y(_05887_));
 AND3x1_ASAP7_75t_R _23445_ (.A(_05291_),
    .B(_05322_),
    .C(_05794_),
    .Y(_05888_));
 AO21x2_ASAP7_75t_R _23446_ (.A1(_05887_),
    .A2(_05788_),
    .B(_05888_),
    .Y(_05889_));
 BUFx2_ASAP7_75t_R input138 (.A(irq_fast_i[3]),
    .Y(net138));
 NAND2x1_ASAP7_75t_R _23448_ (.A(_05803_),
    .B(_05889_),
    .Y(_16812_));
 NAND2x1_ASAP7_75t_R _23449_ (.A(_05828_),
    .B(_05867_),
    .Y(_16818_));
 NAND2x1_ASAP7_75t_R _23450_ (.A(_05846_),
    .B(_05851_),
    .Y(_16828_));
 AND2x2_ASAP7_75t_R _23451_ (.A(_05822_),
    .B(_05871_),
    .Y(_16831_));
 AND2x2_ASAP7_75t_R _23452_ (.A(_05825_),
    .B(_05878_),
    .Y(_16833_));
 AND2x2_ASAP7_75t_R _23453_ (.A(_05812_),
    .B(_05883_),
    .Y(_16832_));
 AO22x2_ASAP7_75t_R _23454_ (.A1(_05119_),
    .A2(_05128_),
    .B1(_05139_),
    .B2(_05150_),
    .Y(_05891_));
 NAND2x1_ASAP7_75t_R _23455_ (.A(_13878_),
    .B(_05798_),
    .Y(_05892_));
 OA21x2_ASAP7_75t_R _23456_ (.A1(_05891_),
    .A2(_05798_),
    .B(_05892_),
    .Y(_05893_));
 BUFx2_ASAP7_75t_R input137 (.A(irq_fast_i[2]),
    .Y(net137));
 BUFx2_ASAP7_75t_R input136 (.A(irq_fast_i[1]),
    .Y(net136));
 NAND2x1_ASAP7_75t_R _23459_ (.A(_05807_),
    .B(_05893_),
    .Y(_16845_));
 OAI22x1_ASAP7_75t_R _23460_ (.A1(_00783_),
    .A2(_05519_),
    .B1(_05791_),
    .B2(_01308_),
    .Y(_17777_));
 BUFx2_ASAP7_75t_R input135 (.A(irq_fast_i[14]),
    .Y(net135));
 OR2x2_ASAP7_75t_R _23462_ (.A(_05420_),
    .B(_05788_),
    .Y(_05897_));
 OA21x2_ASAP7_75t_R _23463_ (.A1(_15617_),
    .A2(_05794_),
    .B(_05897_),
    .Y(_05898_));
 BUFx2_ASAP7_75t_R input134 (.A(irq_fast_i[13]),
    .Y(net134));
 AND2x2_ASAP7_75t_R _23465_ (.A(_05803_),
    .B(_05898_),
    .Y(_17778_));
 AND2x2_ASAP7_75t_R _23466_ (.A(_05815_),
    .B(_05889_),
    .Y(_16860_));
 OR2x2_ASAP7_75t_R _23467_ (.A(_15352_),
    .B(_05794_),
    .Y(_05900_));
 OAI21x1_ASAP7_75t_R _23468_ (.A1(_05213_),
    .A2(_05788_),
    .B(_05900_),
    .Y(_05901_));
 BUFx2_ASAP7_75t_R input133 (.A(irq_fast_i[12]),
    .Y(net133));
 AND2x2_ASAP7_75t_R _23470_ (.A(_05819_),
    .B(_05901_),
    .Y(_16861_));
 AND2x2_ASAP7_75t_R _23471_ (.A(_05828_),
    .B(_05875_),
    .Y(_16862_));
 NAND2x1_ASAP7_75t_R _23472_ (.A(_05835_),
    .B(_05867_),
    .Y(_16866_));
 NAND2x1_ASAP7_75t_R _23473_ (.A(_05846_),
    .B(_05858_),
    .Y(_16875_));
 AND2x2_ASAP7_75t_R _23474_ (.A(_05822_),
    .B(_05878_),
    .Y(_16878_));
 AND2x2_ASAP7_75t_R _23475_ (.A(_05825_),
    .B(_05883_),
    .Y(_16879_));
 AND2x2_ASAP7_75t_R _23476_ (.A(_05812_),
    .B(_05893_),
    .Y(_16880_));
 AND3x1_ASAP7_75t_R _23477_ (.A(_05239_),
    .B(_05260_),
    .C(_05800_),
    .Y(_05903_));
 AO21x2_ASAP7_75t_R _23478_ (.A1(_15401_),
    .A2(_05798_),
    .B(_05903_),
    .Y(_05904_));
 BUFx2_ASAP7_75t_R input132 (.A(irq_fast_i[11]),
    .Y(net132));
 BUFx2_ASAP7_75t_R input131 (.A(irq_fast_i[10]),
    .Y(net131));
 NAND2x1_ASAP7_75t_R _23481_ (.A(_05807_),
    .B(_05904_),
    .Y(_16890_));
 NAND2x2_ASAP7_75t_R _23482_ (.A(_13261_),
    .B(_13263_),
    .Y(_05907_));
 OA21x2_ASAP7_75t_R _23483_ (.A1(_14141_),
    .A2(_05907_),
    .B(_13327_),
    .Y(_05908_));
 NOR2x2_ASAP7_75t_R _23484_ (.A(_13318_),
    .B(_05908_),
    .Y(_05909_));
 NAND2x2_ASAP7_75t_R _23485_ (.A(_05420_),
    .B(_05909_),
    .Y(_05910_));
 OR2x6_ASAP7_75t_R _23486_ (.A(_05788_),
    .B(_05910_),
    .Y(_05911_));
 BUFx2_ASAP7_75t_R input130 (.A(irq_fast_i[0]),
    .Y(net130));
 BUFx2_ASAP7_75t_R input129 (.A(irq_external_i),
    .Y(net129));
 AND2x2_ASAP7_75t_R _23489_ (.A(_05815_),
    .B(_05898_),
    .Y(_16907_));
 AND2x2_ASAP7_75t_R _23490_ (.A(_05819_),
    .B(_05889_),
    .Y(_16908_));
 AND2x2_ASAP7_75t_R _23491_ (.A(_05828_),
    .B(_05901_),
    .Y(_16909_));
 NAND2x1_ASAP7_75t_R _23492_ (.A(_05835_),
    .B(_05875_),
    .Y(_16914_));
 BUFx2_ASAP7_75t_R input128 (.A(instr_rvalid_i),
    .Y(net128));
 NAND2x1_ASAP7_75t_R _23494_ (.A(_05855_),
    .B(_05858_),
    .Y(_16923_));
 AND2x2_ASAP7_75t_R _23495_ (.A(_05832_),
    .B(_05878_),
    .Y(_16928_));
 AND2x2_ASAP7_75t_R _23496_ (.A(_05822_),
    .B(_05883_),
    .Y(_16929_));
 AND2x2_ASAP7_75t_R _23497_ (.A(_05825_),
    .B(_05893_),
    .Y(_16930_));
 NAND2x1_ASAP7_75t_R _23498_ (.A(_05812_),
    .B(_05904_),
    .Y(_16940_));
 NAND2x1_ASAP7_75t_R _23499_ (.A(_00281_),
    .B(_13344_),
    .Y(_05914_));
 AOI21x1_ASAP7_75t_R _23500_ (.A1(_05907_),
    .A2(_05914_),
    .B(_13318_),
    .Y(_05915_));
 AND3x4_ASAP7_75t_R _23501_ (.A(_05474_),
    .B(_05800_),
    .C(_05915_),
    .Y(_05916_));
 BUFx2_ASAP7_75t_R input127 (.A(instr_rdata_i[9]),
    .Y(net127));
 BUFx2_ASAP7_75t_R input126 (.A(instr_rdata_i[8]),
    .Y(net126));
 NAND2x2_ASAP7_75t_R _23504_ (.A(_05796_),
    .B(_05916_),
    .Y(_16995_));
 INVx2_ASAP7_75t_R _23505_ (.A(_16995_),
    .Y(_16948_));
 OA22x2_ASAP7_75t_R _23506_ (.A1(_01314_),
    .A2(_00034_),
    .B1(_05519_),
    .B2(_00849_),
    .Y(_16958_));
 AND2x2_ASAP7_75t_R _23507_ (.A(_05828_),
    .B(_05889_),
    .Y(_16963_));
 AND2x2_ASAP7_75t_R _23508_ (.A(_05835_),
    .B(_05901_),
    .Y(_16964_));
 AND2x2_ASAP7_75t_R _23509_ (.A(_05843_),
    .B(_05875_),
    .Y(_16965_));
 NAND2x1_ASAP7_75t_R _23510_ (.A(_05851_),
    .B(_05867_),
    .Y(_16969_));
 NAND2x1_ASAP7_75t_R _23511_ (.A(_05846_),
    .B(_05871_),
    .Y(_16980_));
 AND2x2_ASAP7_75t_R _23512_ (.A(_05822_),
    .B(_05893_),
    .Y(_16985_));
 AND2x2_ASAP7_75t_R _23513_ (.A(_05825_),
    .B(_05904_),
    .Y(_16986_));
 NAND2x1_ASAP7_75t_R _23514_ (.A(_15555_),
    .B(_05798_),
    .Y(_05919_));
 OA21x2_ASAP7_75t_R _23515_ (.A1(_05369_),
    .A2(_05798_),
    .B(_05919_),
    .Y(_05920_));
 BUFx2_ASAP7_75t_R input125 (.A(instr_rdata_i[7]),
    .Y(net125));
 AND2x2_ASAP7_75t_R _23517_ (.A(_05812_),
    .B(_05920_),
    .Y(_16987_));
 BUFx3_ASAP7_75t_R input124 (.A(instr_rdata_i[6]),
    .Y(net124));
 OR2x2_ASAP7_75t_R _23519_ (.A(_15665_),
    .B(_05800_),
    .Y(_05923_));
 OA21x2_ASAP7_75t_R _23520_ (.A1(_05474_),
    .A2(_05798_),
    .B(_05923_),
    .Y(_05924_));
 BUFx2_ASAP7_75t_R input123 (.A(instr_rdata_i[5]),
    .Y(net123));
 BUFx2_ASAP7_75t_R input122 (.A(instr_rdata_i[4]),
    .Y(net122));
 NAND2x1_ASAP7_75t_R _23523_ (.A(_05807_),
    .B(_05924_),
    .Y(_16996_));
 NOR2x1_ASAP7_75t_R _23524_ (.A(_13217_),
    .B(_05794_),
    .Y(_05927_));
 AO21x2_ASAP7_75t_R _23525_ (.A1(_15841_),
    .A2(_05794_),
    .B(_05927_),
    .Y(_05928_));
 BUFx3_ASAP7_75t_R input121 (.A(instr_rdata_i[3]),
    .Y(net121));
 NAND2x1_ASAP7_75t_R _23527_ (.A(_05916_),
    .B(_05928_),
    .Y(_16997_));
 INVx1_ASAP7_75t_R _23528_ (.A(_16997_),
    .Y(_17044_));
 AO21x2_ASAP7_75t_R _23529_ (.A1(_05907_),
    .A2(_05914_),
    .B(_13318_),
    .Y(_05930_));
 OR3x4_ASAP7_75t_R _23530_ (.A(_01314_),
    .B(_00034_),
    .C(_05930_),
    .Y(_05931_));
 BUFx2_ASAP7_75t_R input120 (.A(instr_rdata_i[31]),
    .Y(net120));
 OA21x2_ASAP7_75t_R _23532_ (.A1(_00881_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17008_));
 AND2x2_ASAP7_75t_R _23533_ (.A(_05835_),
    .B(_05889_),
    .Y(_17013_));
 AND2x2_ASAP7_75t_R _23534_ (.A(_05843_),
    .B(_05901_),
    .Y(_17014_));
 AND2x2_ASAP7_75t_R _23535_ (.A(_05851_),
    .B(_05875_),
    .Y(_17015_));
 NAND2x1_ASAP7_75t_R _23536_ (.A(_05858_),
    .B(_05867_),
    .Y(_17019_));
 NAND2x1_ASAP7_75t_R _23537_ (.A(_05846_),
    .B(_05878_),
    .Y(_17029_));
 NAND2x1_ASAP7_75t_R _23538_ (.A(_05822_),
    .B(_05904_),
    .Y(_17034_));
 AND2x2_ASAP7_75t_R _23539_ (.A(_05807_),
    .B(_05916_),
    .Y(_17045_));
 OA21x2_ASAP7_75t_R _23540_ (.A1(_00914_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17059_));
 AND2x2_ASAP7_75t_R _23541_ (.A(_05843_),
    .B(_05889_),
    .Y(_17064_));
 AND2x2_ASAP7_75t_R _23542_ (.A(_05851_),
    .B(_05901_),
    .Y(_17065_));
 AND2x2_ASAP7_75t_R _23543_ (.A(_05858_),
    .B(_05875_),
    .Y(_17066_));
 NAND2x1_ASAP7_75t_R _23544_ (.A(_05863_),
    .B(_05867_),
    .Y(_17070_));
 NAND2x1_ASAP7_75t_R _23545_ (.A(_05846_),
    .B(_05883_),
    .Y(_17080_));
 BUFx2_ASAP7_75t_R input119 (.A(instr_rdata_i[30]),
    .Y(net119));
 NAND2x1_ASAP7_75t_R _23547_ (.A(_05822_),
    .B(_05920_),
    .Y(_17085_));
 NAND2x2_ASAP7_75t_R _23548_ (.A(_05812_),
    .B(_05916_),
    .Y(_17087_));
 INVx1_ASAP7_75t_R _23549_ (.A(_17087_),
    .Y(_17174_));
 OA21x2_ASAP7_75t_R _23550_ (.A1(_00946_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17103_));
 AND2x2_ASAP7_75t_R _23551_ (.A(_05851_),
    .B(_05889_),
    .Y(_17108_));
 AND2x2_ASAP7_75t_R _23552_ (.A(_05858_),
    .B(_05901_),
    .Y(_17109_));
 AND2x2_ASAP7_75t_R _23553_ (.A(_05863_),
    .B(_05875_),
    .Y(_17110_));
 NAND2x1_ASAP7_75t_R _23554_ (.A(_05867_),
    .B(_05871_),
    .Y(_17114_));
 NAND2x1_ASAP7_75t_R _23555_ (.A(_05846_),
    .B(_05893_),
    .Y(_17124_));
 NAND2x1_ASAP7_75t_R _23556_ (.A(_05822_),
    .B(_05924_),
    .Y(_17129_));
 NAND2x1_ASAP7_75t_R _23557_ (.A(_05825_),
    .B(_05916_),
    .Y(_17130_));
 INVx1_ASAP7_75t_R _23558_ (.A(_17130_),
    .Y(_17175_));
 OA21x2_ASAP7_75t_R _23559_ (.A1(_00979_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17147_));
 NAND2x1_ASAP7_75t_R _23560_ (.A(_05858_),
    .B(_05889_),
    .Y(_17152_));
 NAND2x1_ASAP7_75t_R _23561_ (.A(_05867_),
    .B(_05878_),
    .Y(_17159_));
 NAND2x1_ASAP7_75t_R _23562_ (.A(_05846_),
    .B(_05904_),
    .Y(_17169_));
 AND2x2_ASAP7_75t_R _23563_ (.A(_05822_),
    .B(_05916_),
    .Y(_17176_));
 BUFx2_ASAP7_75t_R input118 (.A(instr_rdata_i[2]),
    .Y(net118));
 OA21x2_ASAP7_75t_R _23565_ (.A1(_01011_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17195_));
 NAND2x1_ASAP7_75t_R _23566_ (.A(_05863_),
    .B(_05889_),
    .Y(_17200_));
 NAND2x1_ASAP7_75t_R _23567_ (.A(_05867_),
    .B(_05883_),
    .Y(_17207_));
 NAND2x1_ASAP7_75t_R _23568_ (.A(_05846_),
    .B(_05920_),
    .Y(_17216_));
 NAND2x2_ASAP7_75t_R _23569_ (.A(_05832_),
    .B(_05916_),
    .Y(_17218_));
 INVx1_ASAP7_75t_R _23570_ (.A(_17218_),
    .Y(_17295_));
 OA21x2_ASAP7_75t_R _23571_ (.A1(_01045_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17238_));
 NAND2x1_ASAP7_75t_R _23572_ (.A(_05871_),
    .B(_05889_),
    .Y(_17243_));
 NAND2x1_ASAP7_75t_R _23573_ (.A(_05867_),
    .B(_05893_),
    .Y(_17250_));
 NAND2x1_ASAP7_75t_R _23574_ (.A(_05846_),
    .B(_05924_),
    .Y(_17259_));
 NAND2x1_ASAP7_75t_R _23575_ (.A(_05840_),
    .B(_05916_),
    .Y(_17260_));
 INVx1_ASAP7_75t_R _23576_ (.A(_17260_),
    .Y(_17296_));
 OA21x2_ASAP7_75t_R _23577_ (.A1(_01077_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17274_));
 NAND2x1_ASAP7_75t_R _23578_ (.A(_05878_),
    .B(_05889_),
    .Y(_17279_));
 NAND2x1_ASAP7_75t_R _23579_ (.A(_05867_),
    .B(_05904_),
    .Y(_17286_));
 AND2x2_ASAP7_75t_R _23580_ (.A(_05846_),
    .B(_05916_),
    .Y(_17297_));
 OA21x2_ASAP7_75t_R _23581_ (.A1(_01110_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17316_));
 NAND2x1_ASAP7_75t_R _23582_ (.A(_05883_),
    .B(_05889_),
    .Y(_17321_));
 NAND2x1_ASAP7_75t_R _23583_ (.A(_05867_),
    .B(_05920_),
    .Y(_17328_));
 NAND2x2_ASAP7_75t_R _23584_ (.A(_05855_),
    .B(_05916_),
    .Y(_17330_));
 INVx1_ASAP7_75t_R _23585_ (.A(_17330_),
    .Y(_17394_));
 OA21x2_ASAP7_75t_R _23586_ (.A1(_01142_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17350_));
 NAND2x1_ASAP7_75t_R _23587_ (.A(_05889_),
    .B(_05893_),
    .Y(_17355_));
 NAND2x1_ASAP7_75t_R _23588_ (.A(_05867_),
    .B(_05924_),
    .Y(_17362_));
 AND3x1_ASAP7_75t_R _23589_ (.A(_04856_),
    .B(_04887_),
    .C(_05794_),
    .Y(_05935_));
 AO21x2_ASAP7_75t_R _23590_ (.A1(_14434_),
    .A2(_05788_),
    .B(_05935_),
    .Y(_05936_));
 BUFx2_ASAP7_75t_R input117 (.A(instr_rdata_i[29]),
    .Y(net117));
 NAND2x1_ASAP7_75t_R _23592_ (.A(_05916_),
    .B(_05936_),
    .Y(_17363_));
 INVx1_ASAP7_75t_R _23593_ (.A(_17363_),
    .Y(_17395_));
 OA21x2_ASAP7_75t_R _23594_ (.A1(_01176_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17382_));
 NAND2x1_ASAP7_75t_R _23595_ (.A(_05889_),
    .B(_05904_),
    .Y(_17387_));
 AND2x2_ASAP7_75t_R _23596_ (.A(_05867_),
    .B(_05916_),
    .Y(_17396_));
 OA21x2_ASAP7_75t_R _23597_ (.A1(_01208_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17412_));
 NAND2x1_ASAP7_75t_R _23598_ (.A(_05889_),
    .B(_05920_),
    .Y(_17417_));
 NAND2x2_ASAP7_75t_R _23599_ (.A(_05875_),
    .B(_05916_),
    .Y(_17419_));
 INVx1_ASAP7_75t_R _23600_ (.A(_17419_),
    .Y(_17466_));
 OA21x2_ASAP7_75t_R _23601_ (.A1(_01242_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17440_));
 NAND2x1_ASAP7_75t_R _23602_ (.A(_05889_),
    .B(_05924_),
    .Y(_17445_));
 NAND2x1_ASAP7_75t_R _23603_ (.A(_05901_),
    .B(_05916_),
    .Y(_17446_));
 INVx1_ASAP7_75t_R _23604_ (.A(_17446_),
    .Y(_17467_));
 OA21x2_ASAP7_75t_R _23605_ (.A1(_01274_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17462_));
 AND2x2_ASAP7_75t_R _23606_ (.A(_05889_),
    .B(_05916_),
    .Y(_17468_));
 OA21x2_ASAP7_75t_R _23607_ (.A1(_01308_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17492_));
 OA21x2_ASAP7_75t_R _23608_ (.A1(_01677_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_17517_));
 INVx1_ASAP7_75t_R _23609_ (.A(_17650_),
    .Y(_16555_));
 OA21x2_ASAP7_75t_R _23610_ (.A1(_01375_),
    .A2(_16555_),
    .B(_01386_),
    .Y(_05938_));
 OA21x2_ASAP7_75t_R _23611_ (.A1(_01385_),
    .A2(_05938_),
    .B(_02313_),
    .Y(_05939_));
 AND3x1_ASAP7_75t_R _23612_ (.A(_01427_),
    .B(_02326_),
    .C(_02322_),
    .Y(_05940_));
 OA211x2_ASAP7_75t_R _23613_ (.A1(_01398_),
    .A2(_05939_),
    .B(_05940_),
    .C(_01411_),
    .Y(_05941_));
 AO21x1_ASAP7_75t_R _23614_ (.A1(_01410_),
    .A2(_02322_),
    .B(_01420_),
    .Y(_05942_));
 AO21x1_ASAP7_75t_R _23615_ (.A1(_01427_),
    .A2(_05942_),
    .B(_01426_),
    .Y(_05943_));
 AO21x1_ASAP7_75t_R _23616_ (.A1(_02326_),
    .A2(_05943_),
    .B(_01432_),
    .Y(_05944_));
 OA21x2_ASAP7_75t_R _23617_ (.A1(_05941_),
    .A2(_05944_),
    .B(_01437_),
    .Y(_05945_));
 OA21x2_ASAP7_75t_R _23618_ (.A1(_01436_),
    .A2(_05945_),
    .B(_02330_),
    .Y(_05946_));
 OR3x1_ASAP7_75t_R _23619_ (.A(_00015_),
    .B(_00009_),
    .C(_00019_),
    .Y(_05947_));
 OR2x2_ASAP7_75t_R _23620_ (.A(_00015_),
    .B(_00016_),
    .Y(_05948_));
 AO21x1_ASAP7_75t_R _23621_ (.A1(_02336_),
    .A2(_05948_),
    .B(_00019_),
    .Y(_05949_));
 AND3x1_ASAP7_75t_R _23622_ (.A(_00025_),
    .B(_00032_),
    .C(_02342_),
    .Y(_05950_));
 OA211x2_ASAP7_75t_R _23623_ (.A1(_05946_),
    .A2(_05947_),
    .B(_05949_),
    .C(_05950_),
    .Y(_05951_));
 AND3x1_ASAP7_75t_R _23624_ (.A(_00024_),
    .B(_00032_),
    .C(_02342_),
    .Y(_05952_));
 AO21x1_ASAP7_75t_R _23625_ (.A1(_00032_),
    .A2(_00029_),
    .B(_05952_),
    .Y(_05953_));
 OR3x1_ASAP7_75t_R _23626_ (.A(_00031_),
    .B(_00038_),
    .C(_00036_),
    .Y(_05954_));
 OR3x1_ASAP7_75t_R _23627_ (.A(_00038_),
    .B(_00036_),
    .C(_02344_),
    .Y(_05955_));
 OA21x2_ASAP7_75t_R _23628_ (.A1(_00038_),
    .A2(_00039_),
    .B(_05955_),
    .Y(_05956_));
 OA31x2_ASAP7_75t_R _23629_ (.A1(_05951_),
    .A2(_05953_),
    .A3(_05954_),
    .B1(_05956_),
    .Y(_05957_));
 AND3x1_ASAP7_75t_R _23630_ (.A(_00045_),
    .B(_02347_),
    .C(_02350_),
    .Y(_05958_));
 AND3x1_ASAP7_75t_R _23631_ (.A(_00045_),
    .B(_00041_),
    .C(_02350_),
    .Y(_05959_));
 AO21x1_ASAP7_75t_R _23632_ (.A1(_00044_),
    .A2(_02350_),
    .B(_05959_),
    .Y(_05960_));
 AO21x1_ASAP7_75t_R _23633_ (.A1(_05957_),
    .A2(_05958_),
    .B(_05960_),
    .Y(_05961_));
 OR3x1_ASAP7_75t_R _23634_ (.A(_00052_),
    .B(_00049_),
    .C(_00054_),
    .Y(_05962_));
 OR2x2_ASAP7_75t_R _23635_ (.A(_00052_),
    .B(_00053_),
    .Y(_05963_));
 AO21x1_ASAP7_75t_R _23636_ (.A1(_02353_),
    .A2(_05963_),
    .B(_00054_),
    .Y(_05964_));
 OA21x2_ASAP7_75t_R _23637_ (.A1(_05961_),
    .A2(_05962_),
    .B(_05964_),
    .Y(_05965_));
 AND3x1_ASAP7_75t_R _23638_ (.A(_00056_),
    .B(_00059_),
    .C(_02354_),
    .Y(_05966_));
 AND3x1_ASAP7_75t_R _23639_ (.A(_00055_),
    .B(_00059_),
    .C(_02354_),
    .Y(_05967_));
 AO221x1_ASAP7_75t_R _23640_ (.A1(_00059_),
    .A2(_00057_),
    .B1(_05965_),
    .B2(_05966_),
    .C(_05967_),
    .Y(_05968_));
 OA21x2_ASAP7_75t_R _23641_ (.A1(_00058_),
    .A2(_05968_),
    .B(_02355_),
    .Y(_05969_));
 OA21x2_ASAP7_75t_R _23642_ (.A1(_00060_),
    .A2(_05969_),
    .B(_00062_),
    .Y(_05970_));
 OA21x2_ASAP7_75t_R _23643_ (.A1(_00061_),
    .A2(_05970_),
    .B(_02356_),
    .Y(_05971_));
 OA21x2_ASAP7_75t_R _23644_ (.A1(_00063_),
    .A2(_05971_),
    .B(_00065_),
    .Y(_05972_));
 OA21x2_ASAP7_75t_R _23645_ (.A1(_00064_),
    .A2(_05972_),
    .B(_00067_),
    .Y(_17532_));
 CKINVDCx14_ASAP7_75t_R _23646_ (.A(_00051_),
    .Y(_17268_));
 CKINVDCx12_ASAP7_75t_R _23647_ (.A(_02352_),
    .Y(_17308_));
 INVx1_ASAP7_75t_R _23648_ (.A(_02357_),
    .Y(_18106_));
 INVx1_ASAP7_75t_R _23649_ (.A(_02064_),
    .Y(\cs_registers_i.mhpmcounter[2][34] ));
 INVx1_ASAP7_75t_R _23650_ (.A(_02170_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[34] ));
 INVx1_ASAP7_75t_R _23651_ (.A(_01486_),
    .Y(\cs_registers_i.mhpmcounter[2][2] ));
 INVx1_ASAP7_75t_R _23652_ (.A(_01517_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[2] ));
 INVx1_ASAP7_75t_R _23653_ (.A(_02062_),
    .Y(\cs_registers_i.mhpmcounter[2][36] ));
 INVx1_ASAP7_75t_R _23654_ (.A(_02168_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[36] ));
 INVx1_ASAP7_75t_R _23655_ (.A(_01484_),
    .Y(\cs_registers_i.mhpmcounter[2][4] ));
 INVx1_ASAP7_75t_R _23656_ (.A(_01515_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[4] ));
 INVx1_ASAP7_75t_R _23657_ (.A(_02060_),
    .Y(\cs_registers_i.mhpmcounter[2][38] ));
 INVx1_ASAP7_75t_R _23658_ (.A(_02166_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[38] ));
 INVx1_ASAP7_75t_R _23659_ (.A(_01482_),
    .Y(\cs_registers_i.mhpmcounter[2][6] ));
 INVx1_ASAP7_75t_R _23660_ (.A(_01513_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[6] ));
 INVx1_ASAP7_75t_R _23661_ (.A(_02058_),
    .Y(\cs_registers_i.mhpmcounter[2][40] ));
 INVx1_ASAP7_75t_R _23662_ (.A(_02164_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[40] ));
 INVx1_ASAP7_75t_R _23663_ (.A(_01480_),
    .Y(\cs_registers_i.mhpmcounter[2][8] ));
 INVx1_ASAP7_75t_R _23664_ (.A(_01511_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[8] ));
 INVx1_ASAP7_75t_R _23665_ (.A(_02056_),
    .Y(\cs_registers_i.mhpmcounter[2][42] ));
 INVx1_ASAP7_75t_R _23666_ (.A(_02162_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[42] ));
 INVx1_ASAP7_75t_R _23667_ (.A(_01478_),
    .Y(\cs_registers_i.mhpmcounter[2][10] ));
 INVx1_ASAP7_75t_R _23668_ (.A(_01509_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[10] ));
 INVx1_ASAP7_75t_R _23669_ (.A(_02052_),
    .Y(\cs_registers_i.mhpmcounter[2][46] ));
 INVx1_ASAP7_75t_R _23670_ (.A(_02158_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[46] ));
 INVx1_ASAP7_75t_R _23671_ (.A(_01474_),
    .Y(\cs_registers_i.mhpmcounter[2][14] ));
 INVx1_ASAP7_75t_R _23672_ (.A(_01505_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[14] ));
 INVx1_ASAP7_75t_R _23673_ (.A(_02050_),
    .Y(\cs_registers_i.mhpmcounter[2][48] ));
 INVx1_ASAP7_75t_R _23674_ (.A(_02156_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[48] ));
 INVx1_ASAP7_75t_R _23675_ (.A(_01472_),
    .Y(\cs_registers_i.mhpmcounter[2][16] ));
 INVx1_ASAP7_75t_R _23676_ (.A(_01503_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[16] ));
 INVx1_ASAP7_75t_R _23677_ (.A(_02048_),
    .Y(\cs_registers_i.mhpmcounter[2][50] ));
 INVx1_ASAP7_75t_R _23678_ (.A(_02154_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[50] ));
 INVx1_ASAP7_75t_R _23679_ (.A(_01470_),
    .Y(\cs_registers_i.mhpmcounter[2][18] ));
 INVx1_ASAP7_75t_R _23680_ (.A(_01501_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[18] ));
 INVx1_ASAP7_75t_R _23681_ (.A(_02046_),
    .Y(\cs_registers_i.mhpmcounter[2][52] ));
 INVx1_ASAP7_75t_R _23682_ (.A(_02152_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[52] ));
 INVx1_ASAP7_75t_R _23683_ (.A(_01468_),
    .Y(\cs_registers_i.mhpmcounter[2][20] ));
 INVx1_ASAP7_75t_R _23684_ (.A(_01499_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[20] ));
 INVx1_ASAP7_75t_R _23685_ (.A(_02044_),
    .Y(\cs_registers_i.mhpmcounter[2][54] ));
 INVx1_ASAP7_75t_R _23686_ (.A(_02150_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[54] ));
 INVx1_ASAP7_75t_R _23687_ (.A(_01466_),
    .Y(\cs_registers_i.mhpmcounter[2][22] ));
 INVx1_ASAP7_75t_R _23688_ (.A(_01497_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[22] ));
 INVx1_ASAP7_75t_R _23689_ (.A(_02042_),
    .Y(\cs_registers_i.mhpmcounter[2][56] ));
 INVx1_ASAP7_75t_R _23690_ (.A(_02148_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[56] ));
 INVx1_ASAP7_75t_R _23691_ (.A(_01464_),
    .Y(\cs_registers_i.mhpmcounter[2][24] ));
 INVx1_ASAP7_75t_R _23692_ (.A(_01495_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[24] ));
 INVx1_ASAP7_75t_R _23693_ (.A(_02040_),
    .Y(\cs_registers_i.mhpmcounter[2][58] ));
 INVx1_ASAP7_75t_R _23694_ (.A(_02146_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[58] ));
 INVx1_ASAP7_75t_R _23695_ (.A(_01462_),
    .Y(\cs_registers_i.mhpmcounter[2][26] ));
 INVx1_ASAP7_75t_R _23696_ (.A(_01493_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[26] ));
 INVx1_ASAP7_75t_R _23697_ (.A(_02038_),
    .Y(\cs_registers_i.mhpmcounter[2][60] ));
 INVx1_ASAP7_75t_R _23698_ (.A(_02144_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[60] ));
 INVx1_ASAP7_75t_R _23699_ (.A(_01460_),
    .Y(\cs_registers_i.mhpmcounter[2][28] ));
 INVx1_ASAP7_75t_R _23700_ (.A(_01491_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[28] ));
 INVx1_ASAP7_75t_R _23701_ (.A(_02036_),
    .Y(\cs_registers_i.mhpmcounter[2][62] ));
 INVx1_ASAP7_75t_R _23702_ (.A(_02142_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[62] ));
 INVx1_ASAP7_75t_R _23703_ (.A(_01458_),
    .Y(\cs_registers_i.mhpmcounter[2][30] ));
 INVx1_ASAP7_75t_R _23704_ (.A(_01489_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[30] ));
 INVx1_ASAP7_75t_R _23705_ (.A(_02391_),
    .Y(_18260_));
 OR3x1_ASAP7_75t_R _23706_ (.A(_01485_),
    .B(_01486_),
    .C(_02391_),
    .Y(_05973_));
 INVx1_ASAP7_75t_R _23707_ (.A(_05973_),
    .Y(_18261_));
 OR5x2_ASAP7_75t_R _23708_ (.A(_01483_),
    .B(_01484_),
    .C(_01485_),
    .D(_01486_),
    .E(_02391_),
    .Y(_05974_));
 INVx1_ASAP7_75t_R _23709_ (.A(_05974_),
    .Y(_18262_));
 OR3x2_ASAP7_75t_R _23710_ (.A(_01481_),
    .B(_01482_),
    .C(_05974_),
    .Y(_05975_));
 INVx1_ASAP7_75t_R _23711_ (.A(_05975_),
    .Y(_18263_));
 OR2x2_ASAP7_75t_R _23712_ (.A(_01479_),
    .B(_01480_),
    .Y(_05976_));
 OR2x2_ASAP7_75t_R _23713_ (.A(_05975_),
    .B(_05976_),
    .Y(_05977_));
 INVx1_ASAP7_75t_R _23714_ (.A(_05977_),
    .Y(_18264_));
 OR2x2_ASAP7_75t_R _23715_ (.A(_01477_),
    .B(_01478_),
    .Y(_05978_));
 OR3x1_ASAP7_75t_R _23716_ (.A(_05975_),
    .B(_05976_),
    .C(_05978_),
    .Y(_05979_));
 INVx1_ASAP7_75t_R _23717_ (.A(_05979_),
    .Y(_18265_));
 OR2x2_ASAP7_75t_R _23718_ (.A(_01475_),
    .B(_01476_),
    .Y(_05980_));
 NOR2x1_ASAP7_75t_R _23719_ (.A(_05979_),
    .B(_05980_),
    .Y(_18266_));
 OR2x2_ASAP7_75t_R _23720_ (.A(_01473_),
    .B(_01474_),
    .Y(_05981_));
 OR5x2_ASAP7_75t_R _23721_ (.A(_05975_),
    .B(_05976_),
    .C(_05978_),
    .D(_05980_),
    .E(_05981_),
    .Y(_05982_));
 INVx1_ASAP7_75t_R _23722_ (.A(_05982_),
    .Y(_18267_));
 OR3x1_ASAP7_75t_R _23723_ (.A(_01471_),
    .B(_01472_),
    .C(_05982_),
    .Y(_05983_));
 INVx1_ASAP7_75t_R _23724_ (.A(_05983_),
    .Y(_18268_));
 OR5x1_ASAP7_75t_R _23725_ (.A(_01469_),
    .B(_01470_),
    .C(_01471_),
    .D(_01472_),
    .E(_05982_),
    .Y(_05984_));
 INVx1_ASAP7_75t_R _23726_ (.A(_05984_),
    .Y(_18269_));
 INVx1_ASAP7_75t_R _23727_ (.A(_01467_),
    .Y(_05985_));
 AND3x1_ASAP7_75t_R _23728_ (.A(_05985_),
    .B(\cs_registers_i.mhpmcounter[2][20] ),
    .C(_18269_),
    .Y(_18270_));
 OR5x2_ASAP7_75t_R _23729_ (.A(_01465_),
    .B(_01466_),
    .C(_01467_),
    .D(_01468_),
    .E(_05984_),
    .Y(_05986_));
 INVx1_ASAP7_75t_R _23730_ (.A(_05986_),
    .Y(_18271_));
 OR3x1_ASAP7_75t_R _23731_ (.A(_01463_),
    .B(_01464_),
    .C(_05986_),
    .Y(_05987_));
 INVx1_ASAP7_75t_R _23732_ (.A(_05987_),
    .Y(_18272_));
 OR5x2_ASAP7_75t_R _23733_ (.A(_01461_),
    .B(_01462_),
    .C(_01463_),
    .D(_01464_),
    .E(_05986_),
    .Y(_05988_));
 INVx1_ASAP7_75t_R _23734_ (.A(_05988_),
    .Y(_18273_));
 INVx1_ASAP7_75t_R _23735_ (.A(_01459_),
    .Y(_05989_));
 AND3x1_ASAP7_75t_R _23736_ (.A(_05989_),
    .B(\cs_registers_i.mhpmcounter[2][28] ),
    .C(_18273_),
    .Y(_18274_));
 OR5x2_ASAP7_75t_R _23737_ (.A(_01457_),
    .B(_01458_),
    .C(_01459_),
    .D(_01460_),
    .E(_05988_),
    .Y(_05990_));
 INVx1_ASAP7_75t_R _23738_ (.A(_05990_),
    .Y(_18275_));
 INVx1_ASAP7_75t_R _23739_ (.A(_02065_),
    .Y(_05991_));
 AND3x1_ASAP7_75t_R _23740_ (.A(_05991_),
    .B(\cs_registers_i.mhpmcounter[2][32] ),
    .C(_18275_),
    .Y(_18276_));
 OR5x2_ASAP7_75t_R _23741_ (.A(_02063_),
    .B(_02064_),
    .C(_02065_),
    .D(_02066_),
    .E(_05990_),
    .Y(_05992_));
 INVx1_ASAP7_75t_R _23742_ (.A(_05992_),
    .Y(_18277_));
 INVx1_ASAP7_75t_R _23743_ (.A(_02061_),
    .Y(_05993_));
 AND3x1_ASAP7_75t_R _23744_ (.A(_05993_),
    .B(\cs_registers_i.mhpmcounter[2][36] ),
    .C(_18277_),
    .Y(_18278_));
 OR5x2_ASAP7_75t_R _23745_ (.A(_02059_),
    .B(_02060_),
    .C(_02061_),
    .D(_02062_),
    .E(_05992_),
    .Y(_05994_));
 INVx1_ASAP7_75t_R _23746_ (.A(_05994_),
    .Y(_18279_));
 OR3x1_ASAP7_75t_R _23747_ (.A(_02057_),
    .B(_02058_),
    .C(_05994_),
    .Y(_05995_));
 INVx1_ASAP7_75t_R _23748_ (.A(_05995_),
    .Y(_18280_));
 OR5x1_ASAP7_75t_R _23749_ (.A(_02055_),
    .B(_02056_),
    .C(_02057_),
    .D(_02058_),
    .E(_05994_),
    .Y(_05996_));
 INVx1_ASAP7_75t_R _23750_ (.A(_05996_),
    .Y(_18281_));
 INVx1_ASAP7_75t_R _23751_ (.A(_02053_),
    .Y(_05997_));
 AND3x1_ASAP7_75t_R _23752_ (.A(_05997_),
    .B(\cs_registers_i.mhpmcounter[2][44] ),
    .C(_18281_),
    .Y(_18282_));
 OR5x2_ASAP7_75t_R _23753_ (.A(_02051_),
    .B(_02052_),
    .C(_02053_),
    .D(_02054_),
    .E(_05996_),
    .Y(_05998_));
 INVx1_ASAP7_75t_R _23754_ (.A(_05998_),
    .Y(_18283_));
 OR3x1_ASAP7_75t_R _23755_ (.A(_02049_),
    .B(_02050_),
    .C(_05998_),
    .Y(_05999_));
 INVx1_ASAP7_75t_R _23756_ (.A(_05999_),
    .Y(_18284_));
 OR3x1_ASAP7_75t_R _23757_ (.A(_02047_),
    .B(_02048_),
    .C(_05999_),
    .Y(_06000_));
 INVx1_ASAP7_75t_R _23758_ (.A(_06000_),
    .Y(_18285_));
 OR3x1_ASAP7_75t_R _23759_ (.A(_02045_),
    .B(_02046_),
    .C(_06000_),
    .Y(_06001_));
 INVx1_ASAP7_75t_R _23760_ (.A(_06001_),
    .Y(_18286_));
 OR5x2_ASAP7_75t_R _23761_ (.A(_02043_),
    .B(_02044_),
    .C(_02045_),
    .D(_02046_),
    .E(_06000_),
    .Y(_06002_));
 INVx1_ASAP7_75t_R _23762_ (.A(_06002_),
    .Y(_18287_));
 OR3x1_ASAP7_75t_R _23763_ (.A(_02041_),
    .B(_02042_),
    .C(_06002_),
    .Y(_06003_));
 INVx1_ASAP7_75t_R _23764_ (.A(_06003_),
    .Y(_18288_));
 OR5x2_ASAP7_75t_R _23765_ (.A(_02039_),
    .B(_02040_),
    .C(_02041_),
    .D(_02042_),
    .E(_06002_),
    .Y(_06004_));
 INVx1_ASAP7_75t_R _23766_ (.A(_06004_),
    .Y(_18289_));
 NOR3x1_ASAP7_75t_R _23767_ (.A(_02037_),
    .B(_02038_),
    .C(_06004_),
    .Y(_18290_));
 INVx1_ASAP7_75t_R _23768_ (.A(_02455_),
    .Y(_18291_));
 OR3x1_ASAP7_75t_R _23769_ (.A(_01516_),
    .B(_01517_),
    .C(_02455_),
    .Y(_06005_));
 INVx1_ASAP7_75t_R _23770_ (.A(_06005_),
    .Y(_18292_));
 OR5x2_ASAP7_75t_R _23771_ (.A(_01514_),
    .B(_01515_),
    .C(_01516_),
    .D(_01517_),
    .E(_02455_),
    .Y(_06006_));
 INVx1_ASAP7_75t_R _23772_ (.A(_06006_),
    .Y(_18293_));
 OR3x2_ASAP7_75t_R _23773_ (.A(_01512_),
    .B(_01513_),
    .C(_06006_),
    .Y(_06007_));
 INVx1_ASAP7_75t_R _23774_ (.A(_06007_),
    .Y(_18294_));
 OR3x1_ASAP7_75t_R _23775_ (.A(_01510_),
    .B(_01511_),
    .C(_06007_),
    .Y(_06008_));
 INVx1_ASAP7_75t_R _23776_ (.A(_06008_),
    .Y(_18295_));
 OR5x2_ASAP7_75t_R _23777_ (.A(_01508_),
    .B(_01509_),
    .C(_01510_),
    .D(_01511_),
    .E(_06007_),
    .Y(_06009_));
 INVx1_ASAP7_75t_R _23778_ (.A(_06009_),
    .Y(_18296_));
 INVx1_ASAP7_75t_R _23779_ (.A(_01506_),
    .Y(_06010_));
 AND3x1_ASAP7_75t_R _23780_ (.A(_06010_),
    .B(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .C(_18296_),
    .Y(_18297_));
 OR5x2_ASAP7_75t_R _23781_ (.A(_01504_),
    .B(_01505_),
    .C(_01506_),
    .D(_01507_),
    .E(_06009_),
    .Y(_06011_));
 INVx1_ASAP7_75t_R _23782_ (.A(_06011_),
    .Y(_18298_));
 OR2x2_ASAP7_75t_R _23783_ (.A(_01502_),
    .B(_01503_),
    .Y(_06012_));
 OR2x2_ASAP7_75t_R _23784_ (.A(_06011_),
    .B(_06012_),
    .Y(_06013_));
 INVx1_ASAP7_75t_R _23785_ (.A(_06013_),
    .Y(_18299_));
 OR3x1_ASAP7_75t_R _23786_ (.A(_01500_),
    .B(_01501_),
    .C(_06013_),
    .Y(_06014_));
 INVx1_ASAP7_75t_R _23787_ (.A(_06014_),
    .Y(_18300_));
 OR2x2_ASAP7_75t_R _23788_ (.A(_01498_),
    .B(_01499_),
    .Y(_06015_));
 OR5x2_ASAP7_75t_R _23789_ (.A(_01500_),
    .B(_01501_),
    .C(_06011_),
    .D(_06012_),
    .E(_06015_),
    .Y(_06016_));
 INVx1_ASAP7_75t_R _23790_ (.A(_06016_),
    .Y(_18301_));
 OR2x2_ASAP7_75t_R _23791_ (.A(_01496_),
    .B(_01497_),
    .Y(_06017_));
 OR2x2_ASAP7_75t_R _23792_ (.A(_06016_),
    .B(_06017_),
    .Y(_06018_));
 INVx1_ASAP7_75t_R _23793_ (.A(_06018_),
    .Y(_18302_));
 OR2x2_ASAP7_75t_R _23794_ (.A(_01494_),
    .B(_01495_),
    .Y(_06019_));
 OR3x1_ASAP7_75t_R _23795_ (.A(_06016_),
    .B(_06017_),
    .C(_06019_),
    .Y(_06020_));
 INVx1_ASAP7_75t_R _23796_ (.A(_06020_),
    .Y(_18303_));
 OR2x2_ASAP7_75t_R _23797_ (.A(_01492_),
    .B(_01493_),
    .Y(_06021_));
 OR2x2_ASAP7_75t_R _23798_ (.A(_06020_),
    .B(_06021_),
    .Y(_06022_));
 INVx1_ASAP7_75t_R _23799_ (.A(_06022_),
    .Y(_18304_));
 OR2x2_ASAP7_75t_R _23800_ (.A(_01490_),
    .B(_01491_),
    .Y(_06023_));
 OR5x2_ASAP7_75t_R _23801_ (.A(_06016_),
    .B(_06017_),
    .C(_06019_),
    .D(_06021_),
    .E(_06023_),
    .Y(_06024_));
 INVx1_ASAP7_75t_R _23802_ (.A(_06024_),
    .Y(_18305_));
 OR3x4_ASAP7_75t_R _23803_ (.A(_01488_),
    .B(_01489_),
    .C(_06024_),
    .Y(_06025_));
 INVx1_ASAP7_75t_R _23804_ (.A(_06025_),
    .Y(_18306_));
 OR3x1_ASAP7_75t_R _23805_ (.A(_02171_),
    .B(_02172_),
    .C(_06025_),
    .Y(_06026_));
 INVx1_ASAP7_75t_R _23806_ (.A(_06026_),
    .Y(_18307_));
 OR4x1_ASAP7_75t_R _23807_ (.A(_02169_),
    .B(_02170_),
    .C(_02171_),
    .D(_02172_),
    .Y(_06027_));
 NOR2x1_ASAP7_75t_R _23808_ (.A(_06025_),
    .B(_06027_),
    .Y(_18308_));
 OR3x1_ASAP7_75t_R _23809_ (.A(_02167_),
    .B(_02168_),
    .C(_06027_),
    .Y(_06028_));
 NOR2x1_ASAP7_75t_R _23810_ (.A(_06025_),
    .B(_06028_),
    .Y(_18309_));
 OR2x2_ASAP7_75t_R _23811_ (.A(_02165_),
    .B(_02166_),
    .Y(_06029_));
 OR5x2_ASAP7_75t_R _23812_ (.A(_01488_),
    .B(_01489_),
    .C(_06024_),
    .D(_06028_),
    .E(_06029_),
    .Y(_06030_));
 INVx1_ASAP7_75t_R _23813_ (.A(_06030_),
    .Y(_18310_));
 NOR3x2_ASAP7_75t_R _23814_ (.B(_02164_),
    .C(_06030_),
    .Y(_18311_),
    .A(_02163_));
 NOR2x2_ASAP7_75t_R _23815_ (.A(_02161_),
    .B(_02162_),
    .Y(_06031_));
 AND2x2_ASAP7_75t_R _23816_ (.A(_18311_),
    .B(_06031_),
    .Y(_18312_));
 NOR2x1_ASAP7_75t_R _23817_ (.A(_02159_),
    .B(_02160_),
    .Y(_06032_));
 AND3x1_ASAP7_75t_R _23818_ (.A(_18311_),
    .B(_06031_),
    .C(_06032_),
    .Y(_18313_));
 INVx1_ASAP7_75t_R _23819_ (.A(_02157_),
    .Y(_06033_));
 AND5x2_ASAP7_75t_R _23820_ (.A(_06033_),
    .B(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .C(_18311_),
    .D(_06031_),
    .E(_06032_),
    .Y(_18314_));
 INVx1_ASAP7_75t_R _23821_ (.A(_02155_),
    .Y(_06034_));
 AND3x2_ASAP7_75t_R _23822_ (.A(_06034_),
    .B(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .C(_18314_),
    .Y(_18315_));
 NOR2x1_ASAP7_75t_R _23823_ (.A(_02153_),
    .B(_02154_),
    .Y(_06035_));
 NAND2x1_ASAP7_75t_R _23824_ (.A(_18315_),
    .B(_06035_),
    .Y(_06036_));
 INVx1_ASAP7_75t_R _23825_ (.A(_06036_),
    .Y(_18316_));
 OR3x4_ASAP7_75t_R _23826_ (.A(_02151_),
    .B(_02152_),
    .C(_06036_),
    .Y(_06037_));
 INVx1_ASAP7_75t_R _23827_ (.A(_06037_),
    .Y(_18317_));
 NOR3x2_ASAP7_75t_R _23828_ (.B(_02150_),
    .C(_06037_),
    .Y(_18318_),
    .A(_02149_));
 INVx1_ASAP7_75t_R _23829_ (.A(_02147_),
    .Y(_06038_));
 AND3x1_ASAP7_75t_R _23830_ (.A(_06038_),
    .B(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .C(_18318_),
    .Y(_18319_));
 INVx1_ASAP7_75t_R _23831_ (.A(_02145_),
    .Y(_06039_));
 AND3x1_ASAP7_75t_R _23832_ (.A(_06039_),
    .B(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .C(_18319_),
    .Y(_18320_));
 INVx1_ASAP7_75t_R _23833_ (.A(_02143_),
    .Y(_06040_));
 AND3x1_ASAP7_75t_R _23834_ (.A(_06040_),
    .B(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .C(_18320_),
    .Y(_18321_));
 INVx1_ASAP7_75t_R _23835_ (.A(_01606_),
    .Y(\cs_registers_i.pc_if_i[3] ));
 INVx1_ASAP7_75t_R _23836_ (.A(_01604_),
    .Y(\cs_registers_i.pc_if_i[5] ));
 INVx1_ASAP7_75t_R _23837_ (.A(_01602_),
    .Y(\cs_registers_i.pc_if_i[7] ));
 INVx1_ASAP7_75t_R _23838_ (.A(_01600_),
    .Y(\cs_registers_i.pc_if_i[9] ));
 INVx1_ASAP7_75t_R _23839_ (.A(_01598_),
    .Y(\cs_registers_i.pc_if_i[11] ));
 INVx1_ASAP7_75t_R _23840_ (.A(_01596_),
    .Y(\cs_registers_i.pc_if_i[13] ));
 INVx1_ASAP7_75t_R _23841_ (.A(_01594_),
    .Y(\cs_registers_i.pc_if_i[15] ));
 INVx1_ASAP7_75t_R _23842_ (.A(_01592_),
    .Y(\cs_registers_i.pc_if_i[17] ));
 INVx1_ASAP7_75t_R _23843_ (.A(_01590_),
    .Y(\cs_registers_i.pc_if_i[19] ));
 INVx1_ASAP7_75t_R _23844_ (.A(_01588_),
    .Y(\cs_registers_i.pc_if_i[21] ));
 INVx1_ASAP7_75t_R _23845_ (.A(_01586_),
    .Y(\cs_registers_i.pc_if_i[23] ));
 INVx1_ASAP7_75t_R _23846_ (.A(_01584_),
    .Y(\cs_registers_i.pc_if_i[25] ));
 INVx1_ASAP7_75t_R _23847_ (.A(_01582_),
    .Y(\cs_registers_i.pc_if_i[27] ));
 INVx1_ASAP7_75t_R _23848_ (.A(_01580_),
    .Y(\cs_registers_i.pc_if_i[29] ));
 INVx1_ASAP7_75t_R _23849_ (.A(_02519_),
    .Y(_18322_));
 OR3x1_ASAP7_75t_R _23850_ (.A(_00170_),
    .B(_00174_),
    .C(_02519_),
    .Y(_06041_));
 INVx1_ASAP7_75t_R _23851_ (.A(_06041_),
    .Y(_18323_));
 OR5x2_ASAP7_75t_R _23852_ (.A(_00170_),
    .B(_00174_),
    .C(_00177_),
    .D(_00180_),
    .E(_02519_),
    .Y(_06042_));
 INVx1_ASAP7_75t_R _23853_ (.A(_06042_),
    .Y(_18324_));
 OR3x1_ASAP7_75t_R _23854_ (.A(_00182_),
    .B(_00186_),
    .C(_06042_),
    .Y(_06043_));
 INVx1_ASAP7_75t_R _23855_ (.A(_06043_),
    .Y(_18325_));
 OR3x1_ASAP7_75t_R _23856_ (.A(_00189_),
    .B(_00193_),
    .C(_06043_),
    .Y(_06044_));
 INVx1_ASAP7_75t_R _23857_ (.A(_06044_),
    .Y(_18326_));
 OR5x2_ASAP7_75t_R _23858_ (.A(_00189_),
    .B(_00193_),
    .C(_00196_),
    .D(_00199_),
    .E(_06043_),
    .Y(_06045_));
 INVx1_ASAP7_75t_R _23859_ (.A(_06045_),
    .Y(_18327_));
 OR3x1_ASAP7_75t_R _23860_ (.A(_00201_),
    .B(_00204_),
    .C(_06045_),
    .Y(_06046_));
 INVx1_ASAP7_75t_R _23861_ (.A(_06046_),
    .Y(_18328_));
 OR3x1_ASAP7_75t_R _23862_ (.A(_00206_),
    .B(_00208_),
    .C(_06046_),
    .Y(_06047_));
 INVx1_ASAP7_75t_R _23863_ (.A(_06047_),
    .Y(_18329_));
 OR3x1_ASAP7_75t_R _23864_ (.A(_00209_),
    .B(_00211_),
    .C(_06047_),
    .Y(_06048_));
 INVx1_ASAP7_75t_R _23865_ (.A(_06048_),
    .Y(_18330_));
 OR3x1_ASAP7_75t_R _23866_ (.A(_00212_),
    .B(_00214_),
    .C(_06048_),
    .Y(_06049_));
 INVx1_ASAP7_75t_R _23867_ (.A(_06049_),
    .Y(_18331_));
 OR3x1_ASAP7_75t_R _23868_ (.A(_00215_),
    .B(_00217_),
    .C(_06049_),
    .Y(_06050_));
 INVx1_ASAP7_75t_R _23869_ (.A(_06050_),
    .Y(_18332_));
 OR3x1_ASAP7_75t_R _23870_ (.A(_00218_),
    .B(_00220_),
    .C(_06050_),
    .Y(_06051_));
 INVx1_ASAP7_75t_R _23871_ (.A(_06051_),
    .Y(_18333_));
 OR3x1_ASAP7_75t_R _23872_ (.A(_00221_),
    .B(_00223_),
    .C(_06051_),
    .Y(_06052_));
 INVx1_ASAP7_75t_R _23873_ (.A(_06052_),
    .Y(_18334_));
 OR3x1_ASAP7_75t_R _23874_ (.A(_00224_),
    .B(_00226_),
    .C(_06052_),
    .Y(_06053_));
 INVx1_ASAP7_75t_R _23875_ (.A(_06053_),
    .Y(_18335_));
 BUFx2_ASAP7_75t_R input116 (.A(instr_rdata_i[28]),
    .Y(net116));
 BUFx2_ASAP7_75t_R input115 (.A(instr_rdata_i[27]),
    .Y(net115));
 BUFx2_ASAP7_75t_R input114 (.A(instr_rdata_i[26]),
    .Y(net114));
 BUFx2_ASAP7_75t_R input113 (.A(instr_rdata_i[25]),
    .Y(net113));
 BUFx2_ASAP7_75t_R input112 (.A(instr_rdata_i[24]),
    .Y(net112));
 BUFx2_ASAP7_75t_R input111 (.A(instr_rdata_i[23]),
    .Y(net111));
 INVx1_ASAP7_75t_R _23882_ (.A(_14316_),
    .Y(_06060_));
 OA222x2_ASAP7_75t_R _23883_ (.A1(net276),
    .A2(_15731_),
    .B1(_04668_),
    .B2(_00232_),
    .C1(_02537_),
    .C2(_06060_),
    .Y(_06061_));
 NAND2x1_ASAP7_75t_R _23884_ (.A(_18337_),
    .B(_06061_),
    .Y(_06062_));
 OA21x2_ASAP7_75t_R _23885_ (.A1(_18337_),
    .A2(_13640_),
    .B(_06062_),
    .Y(net186));
 AND2x2_ASAP7_75t_R _23886_ (.A(_13196_),
    .B(_13216_),
    .Y(_06063_));
 NAND3x2_ASAP7_75t_R _23887_ (.B(_13177_),
    .C(_06063_),
    .Y(_06064_),
    .A(_13151_));
 CKINVDCx8_ASAP7_75t_R _23888_ (.A(_00232_),
    .Y(_06065_));
 BUFx2_ASAP7_75t_R input110 (.A(instr_rdata_i[22]),
    .Y(net110));
 CKINVDCx6p67_ASAP7_75t_R _23890_ (.A(net277),
    .Y(_06067_));
 CKINVDCx8_ASAP7_75t_R _23891_ (.A(net276),
    .Y(_06068_));
 BUFx2_ASAP7_75t_R input109 (.A(instr_rdata_i[21]),
    .Y(net109));
 CKINVDCx20_ASAP7_75t_R _23893_ (.A(net274),
    .Y(_06070_));
 BUFx2_ASAP7_75t_R input108 (.A(instr_rdata_i[20]),
    .Y(net108));
 AO221x1_ASAP7_75t_R _23895_ (.A1(_06067_),
    .A2(_14373_),
    .B1(_15841_),
    .B2(_06068_),
    .C(_06070_),
    .Y(_06072_));
 AO21x1_ASAP7_75t_R _23896_ (.A1(_06065_),
    .A2(_05853_),
    .B(_06072_),
    .Y(_06073_));
 OA21x2_ASAP7_75t_R _23897_ (.A1(net273),
    .A2(_06064_),
    .B(_06073_),
    .Y(net197));
 BUFx3_ASAP7_75t_R input107 (.A(instr_rdata_i[1]),
    .Y(net107));
 BUFx2_ASAP7_75t_R input106 (.A(instr_rdata_i[19]),
    .Y(net106));
 OA21x2_ASAP7_75t_R _23900_ (.A1(_02537_),
    .A2(_05672_),
    .B(_18337_),
    .Y(_06076_));
 OA21x2_ASAP7_75t_R _23901_ (.A1(net276),
    .A2(_15971_),
    .B(_06076_),
    .Y(_06077_));
 OAI21x1_ASAP7_75t_R _23902_ (.A1(_00232_),
    .A2(_04888_),
    .B(_06077_),
    .Y(_06078_));
 OA21x2_ASAP7_75t_R _23903_ (.A1(_18337_),
    .A2(_13943_),
    .B(_06078_),
    .Y(net208));
 BUFx2_ASAP7_75t_R input105 (.A(instr_rdata_i[18]),
    .Y(net105));
 OA222x2_ASAP7_75t_R _23905_ (.A1(net276),
    .A2(_16083_),
    .B1(_04996_),
    .B2(_00232_),
    .C1(_02537_),
    .C2(_15160_),
    .Y(_06080_));
 NOR2x1_ASAP7_75t_R _23906_ (.A(_06070_),
    .B(_06080_),
    .Y(_06081_));
 AO21x2_ASAP7_75t_R _23907_ (.A1(_06070_),
    .A2(_14019_),
    .B(_06081_),
    .Y(net211));
 OA222x2_ASAP7_75t_R _23908_ (.A1(net276),
    .A2(_16205_),
    .B1(_05105_),
    .B2(_00232_),
    .C1(net277),
    .C2(_15266_),
    .Y(_06082_));
 NAND2x1_ASAP7_75t_R _23909_ (.A(net273),
    .B(_06082_),
    .Y(_06083_));
 OA21x2_ASAP7_75t_R _23910_ (.A1(net273),
    .A2(_14080_),
    .B(_06083_),
    .Y(net212));
 OA222x2_ASAP7_75t_R _23911_ (.A1(_00231_),
    .A2(_16324_),
    .B1(_05213_),
    .B2(_00232_),
    .C1(_02537_),
    .C2(_15352_),
    .Y(_06084_));
 NAND2x1_ASAP7_75t_R _23912_ (.A(_18337_),
    .B(_06084_),
    .Y(_06085_));
 OA21x2_ASAP7_75t_R _23913_ (.A1(_18337_),
    .A2(_14137_),
    .B(_06085_),
    .Y(net213));
 BUFx3_ASAP7_75t_R input104 (.A(instr_rdata_i[17]),
    .Y(net104));
 OA222x2_ASAP7_75t_R _23915_ (.A1(net276),
    .A2(_16433_),
    .B1(_05323_),
    .B2(_00232_),
    .C1(net277),
    .C2(_15507_),
    .Y(_06087_));
 NAND2x1_ASAP7_75t_R _23916_ (.A(net273),
    .B(_06087_),
    .Y(_06088_));
 OA21x2_ASAP7_75t_R _23917_ (.A1(net273),
    .A2(_14197_),
    .B(_06088_),
    .Y(net214));
 BUFx2_ASAP7_75t_R input103 (.A(instr_rdata_i[16]),
    .Y(net103));
 AO221x1_ASAP7_75t_R _23919_ (.A1(_06068_),
    .A2(_04547_),
    .B1(_05420_),
    .B2(_06065_),
    .C(_06070_),
    .Y(_06090_));
 AO21x1_ASAP7_75t_R _23920_ (.A1(_06067_),
    .A2(_15617_),
    .B(_06090_),
    .Y(_06091_));
 OA21x2_ASAP7_75t_R _23921_ (.A1(net273),
    .A2(_05838_),
    .B(_06091_),
    .Y(net215));
 BUFx2_ASAP7_75t_R input102 (.A(instr_rdata_i[15]),
    .Y(net102));
 NAND2x1_ASAP7_75t_R _23923_ (.A(_06065_),
    .B(_13640_),
    .Y(_06093_));
 OA211x2_ASAP7_75t_R _23924_ (.A1(net277),
    .A2(_15731_),
    .B(_06093_),
    .C(net273),
    .Y(_06094_));
 OAI21x1_ASAP7_75t_R _23925_ (.A1(net276),
    .A2(_04668_),
    .B(_06094_),
    .Y(_06095_));
 OA21x2_ASAP7_75t_R _23926_ (.A1(net273),
    .A2(_14316_),
    .B(_06095_),
    .Y(net216));
 AO221x1_ASAP7_75t_R _23927_ (.A1(_06065_),
    .A2(_06064_),
    .B1(_15841_),
    .B2(_06067_),
    .C(_06070_),
    .Y(_06096_));
 AND3x1_ASAP7_75t_R _23928_ (.A(_06068_),
    .B(_04748_),
    .C(_04779_),
    .Y(_06097_));
 OA22x2_ASAP7_75t_R _23929_ (.A1(net273),
    .A2(_14373_),
    .B1(_06096_),
    .B2(_06097_),
    .Y(net217));
 AOI221x1_ASAP7_75t_R _23930_ (.A1(_13614_),
    .A2(_13896_),
    .B1(_13923_),
    .B2(net314),
    .C(_13942_),
    .Y(_06098_));
 OA21x2_ASAP7_75t_R _23931_ (.A1(_00232_),
    .A2(_06098_),
    .B(net273),
    .Y(_06099_));
 OA21x2_ASAP7_75t_R _23932_ (.A1(net277),
    .A2(_15971_),
    .B(_06099_),
    .Y(_06100_));
 OAI21x1_ASAP7_75t_R _23933_ (.A1(net276),
    .A2(_04888_),
    .B(_06100_),
    .Y(_06101_));
 OA21x2_ASAP7_75t_R _23934_ (.A1(net273),
    .A2(_14434_),
    .B(_06101_),
    .Y(net187));
 INVx1_ASAP7_75t_R _23935_ (.A(_14019_),
    .Y(_06102_));
 OA222x2_ASAP7_75t_R _23936_ (.A1(_00232_),
    .A2(_06102_),
    .B1(_16083_),
    .B2(_02537_),
    .C1(_04996_),
    .C2(_00231_),
    .Y(_06103_));
 NAND2x1_ASAP7_75t_R _23937_ (.A(_18337_),
    .B(_06103_),
    .Y(_06104_));
 OA21x2_ASAP7_75t_R _23938_ (.A1(_18337_),
    .A2(_14489_),
    .B(_06104_),
    .Y(net188));
 BUFx2_ASAP7_75t_R input101 (.A(instr_rdata_i[14]),
    .Y(net101));
 AOI221x1_ASAP7_75t_R _23940_ (.A1(_06065_),
    .A2(_14080_),
    .B1(_16204_),
    .B2(_06067_),
    .C(_06070_),
    .Y(_06106_));
 OA21x2_ASAP7_75t_R _23941_ (.A1(net276),
    .A2(_05105_),
    .B(_06106_),
    .Y(_06107_));
 AOI21x1_ASAP7_75t_R _23942_ (.A1(_06070_),
    .A2(_15266_),
    .B(_06107_),
    .Y(net189));
 INVx2_ASAP7_75t_R _23943_ (.A(_14137_),
    .Y(_06108_));
 OA222x2_ASAP7_75t_R _23944_ (.A1(_00232_),
    .A2(_06108_),
    .B1(_16324_),
    .B2(_02537_),
    .C1(_05213_),
    .C2(_00231_),
    .Y(_06109_));
 OR2x2_ASAP7_75t_R _23945_ (.A(_18337_),
    .B(_15352_),
    .Y(_06110_));
 OAI21x1_ASAP7_75t_R _23946_ (.A1(_06070_),
    .A2(_06109_),
    .B(_06110_),
    .Y(net190));
 OA222x2_ASAP7_75t_R _23947_ (.A1(_00232_),
    .A2(_05605_),
    .B1(_16433_),
    .B2(net277),
    .C1(_05323_),
    .C2(net276),
    .Y(_06111_));
 NOR2x1_ASAP7_75t_R _23948_ (.A(_06070_),
    .B(_06111_),
    .Y(_06112_));
 AO21x2_ASAP7_75t_R _23949_ (.A1(_06070_),
    .A2(_05887_),
    .B(_06112_),
    .Y(net191));
 AO221x1_ASAP7_75t_R _23950_ (.A1(_06065_),
    .A2(_05838_),
    .B1(_05420_),
    .B2(_06068_),
    .C(_06070_),
    .Y(_06113_));
 AO21x1_ASAP7_75t_R _23951_ (.A1(_06067_),
    .A2(_04547_),
    .B(_06113_),
    .Y(_06114_));
 OA21x2_ASAP7_75t_R _23952_ (.A1(_18337_),
    .A2(_15617_),
    .B(_06114_),
    .Y(net192));
 AO222x2_ASAP7_75t_R _23953_ (.A1(_06068_),
    .A2(_13640_),
    .B1(_14316_),
    .B2(_06065_),
    .C1(_04667_),
    .C2(_06067_),
    .Y(_06115_));
 AND3x1_ASAP7_75t_R _23954_ (.A(_06070_),
    .B(_15699_),
    .C(_15730_),
    .Y(_06116_));
 AO21x2_ASAP7_75t_R _23955_ (.A1(net274),
    .A2(_06115_),
    .B(_06116_),
    .Y(net193));
 AOI22x1_ASAP7_75t_R _23956_ (.A1(_06068_),
    .A2(_06064_),
    .B1(_14373_),
    .B2(_06065_),
    .Y(_06117_));
 OA211x2_ASAP7_75t_R _23957_ (.A1(net277),
    .A2(_04780_),
    .B(_06117_),
    .C(net273),
    .Y(_06118_));
 AOI21x1_ASAP7_75t_R _23958_ (.A1(_06070_),
    .A2(_15842_),
    .B(_06118_),
    .Y(net194));
 AOI22x1_ASAP7_75t_R _23959_ (.A1(_06068_),
    .A2(_13943_),
    .B1(_14434_),
    .B2(_06065_),
    .Y(_06119_));
 OA211x2_ASAP7_75t_R _23960_ (.A1(_02537_),
    .A2(_04888_),
    .B(_06119_),
    .C(_18337_),
    .Y(_06120_));
 AOI21x1_ASAP7_75t_R _23961_ (.A1(_06070_),
    .A2(_15971_),
    .B(_06120_),
    .Y(net195));
 AOI22x1_ASAP7_75t_R _23962_ (.A1(_06068_),
    .A2(_14019_),
    .B1(_14489_),
    .B2(_06065_),
    .Y(_06121_));
 OA211x2_ASAP7_75t_R _23963_ (.A1(_02537_),
    .A2(_04996_),
    .B(_06121_),
    .C(_18337_),
    .Y(_06122_));
 AOI21x1_ASAP7_75t_R _23964_ (.A1(_06070_),
    .A2(_16083_),
    .B(_06122_),
    .Y(net196));
 INVx1_ASAP7_75t_R _23965_ (.A(_14080_),
    .Y(_06123_));
 OA222x2_ASAP7_75t_R _23966_ (.A1(net276),
    .A2(_06123_),
    .B1(_15266_),
    .B2(_00232_),
    .C1(_05105_),
    .C2(net277),
    .Y(_06124_));
 NOR2x1_ASAP7_75t_R _23967_ (.A(_06070_),
    .B(_06124_),
    .Y(_06125_));
 AO21x1_ASAP7_75t_R _23968_ (.A1(_06070_),
    .A2(_16204_),
    .B(_06125_),
    .Y(net198));
 OA222x2_ASAP7_75t_R _23969_ (.A1(_00231_),
    .A2(_06108_),
    .B1(_15352_),
    .B2(_00232_),
    .C1(_05213_),
    .C2(_02537_),
    .Y(_06126_));
 OR2x2_ASAP7_75t_R _23970_ (.A(_18337_),
    .B(_16324_),
    .Y(_06127_));
 OAI21x1_ASAP7_75t_R _23971_ (.A1(_06070_),
    .A2(_06126_),
    .B(_06127_),
    .Y(net199));
 OA222x2_ASAP7_75t_R _23972_ (.A1(net276),
    .A2(_05605_),
    .B1(_15507_),
    .B2(_00232_),
    .C1(_05323_),
    .C2(net277),
    .Y(_06128_));
 OR2x2_ASAP7_75t_R _23973_ (.A(_06070_),
    .B(_06128_),
    .Y(_06129_));
 OAI21x1_ASAP7_75t_R _23974_ (.A1(net273),
    .A2(_16433_),
    .B(_06129_),
    .Y(net200));
 AO221x1_ASAP7_75t_R _23975_ (.A1(_06068_),
    .A2(_05838_),
    .B1(_05420_),
    .B2(_06067_),
    .C(_06070_),
    .Y(_06130_));
 AO21x1_ASAP7_75t_R _23976_ (.A1(_06065_),
    .A2(_15617_),
    .B(_06130_),
    .Y(_06131_));
 OA21x2_ASAP7_75t_R _23977_ (.A1(_18337_),
    .A2(_04547_),
    .B(_06131_),
    .Y(net201));
 AOI22x1_ASAP7_75t_R _23978_ (.A1(_06067_),
    .A2(_13640_),
    .B1(_14316_),
    .B2(_06068_),
    .Y(_06132_));
 OA211x2_ASAP7_75t_R _23979_ (.A1(_00232_),
    .A2(_15731_),
    .B(_06132_),
    .C(net273),
    .Y(_06133_));
 AOI21x1_ASAP7_75t_R _23980_ (.A1(_06070_),
    .A2(_04668_),
    .B(_06133_),
    .Y(net202));
 AO221x1_ASAP7_75t_R _23981_ (.A1(_06067_),
    .A2(_06064_),
    .B1(_14373_),
    .B2(_06068_),
    .C(_06070_),
    .Y(_06134_));
 AO21x1_ASAP7_75t_R _23982_ (.A1(_06065_),
    .A2(_15841_),
    .B(_06134_),
    .Y(_06135_));
 OA21x2_ASAP7_75t_R _23983_ (.A1(net273),
    .A2(_05853_),
    .B(_06135_),
    .Y(net203));
 AOI22x1_ASAP7_75t_R _23984_ (.A1(_06067_),
    .A2(_13943_),
    .B1(_14434_),
    .B2(_06068_),
    .Y(_06136_));
 OA211x2_ASAP7_75t_R _23985_ (.A1(_00232_),
    .A2(_15971_),
    .B(_06136_),
    .C(net273),
    .Y(_06137_));
 AOI21x1_ASAP7_75t_R _23986_ (.A1(_06070_),
    .A2(_04888_),
    .B(_06137_),
    .Y(net204));
 AOI22x1_ASAP7_75t_R _23987_ (.A1(_06067_),
    .A2(_14019_),
    .B1(_14489_),
    .B2(_06068_),
    .Y(_06138_));
 OA211x2_ASAP7_75t_R _23988_ (.A1(_00232_),
    .A2(_16083_),
    .B(_06138_),
    .C(_18337_),
    .Y(_06139_));
 AOI21x1_ASAP7_75t_R _23989_ (.A1(_06070_),
    .A2(_04996_),
    .B(_06139_),
    .Y(net205));
 OA222x2_ASAP7_75t_R _23990_ (.A1(net276),
    .A2(_15266_),
    .B1(_16205_),
    .B2(_00232_),
    .C1(net277),
    .C2(_06123_),
    .Y(_06140_));
 OR2x2_ASAP7_75t_R _23991_ (.A(net273),
    .B(_05105_),
    .Y(_06141_));
 OAI21x1_ASAP7_75t_R _23992_ (.A1(_06070_),
    .A2(_06140_),
    .B(_06141_),
    .Y(net206));
 OA222x2_ASAP7_75t_R _23993_ (.A1(_00231_),
    .A2(_15352_),
    .B1(_16324_),
    .B2(_00232_),
    .C1(_02537_),
    .C2(_06108_),
    .Y(_06142_));
 OR2x2_ASAP7_75t_R _23994_ (.A(_18337_),
    .B(_05213_),
    .Y(_06143_));
 OAI21x1_ASAP7_75t_R _23995_ (.A1(_06070_),
    .A2(_06142_),
    .B(_06143_),
    .Y(net207));
 OA222x2_ASAP7_75t_R _23996_ (.A1(net276),
    .A2(_15507_),
    .B1(_16433_),
    .B2(_00232_),
    .C1(net277),
    .C2(_05605_),
    .Y(_06144_));
 OR2x2_ASAP7_75t_R _23997_ (.A(net273),
    .B(_05323_),
    .Y(_06145_));
 OAI21x1_ASAP7_75t_R _23998_ (.A1(_06070_),
    .A2(_06144_),
    .B(_06145_),
    .Y(net209));
 AO21x1_ASAP7_75t_R _23999_ (.A1(_06067_),
    .A2(_05838_),
    .B(_06070_),
    .Y(_06146_));
 AO221x1_ASAP7_75t_R _24000_ (.A1(_06068_),
    .A2(_15617_),
    .B1(_04547_),
    .B2(_06065_),
    .C(_06146_),
    .Y(_06147_));
 OA21x2_ASAP7_75t_R _24001_ (.A1(net273),
    .A2(_05420_),
    .B(_06147_),
    .Y(net210));
 NAND2x2_ASAP7_75t_R _24002_ (.A(_00282_),
    .B(_14615_),
    .Y(_06148_));
 AND2x2_ASAP7_75t_R _24003_ (.A(_13261_),
    .B(_02534_),
    .Y(_06149_));
 AO21x1_ASAP7_75t_R _24004_ (.A1(_00281_),
    .A2(_06070_),
    .B(_06149_),
    .Y(_06150_));
 NAND2x1_ASAP7_75t_R _24005_ (.A(_02535_),
    .B(_06148_),
    .Y(_06151_));
 OA21x2_ASAP7_75t_R _24006_ (.A1(_06148_),
    .A2(_06150_),
    .B(_06151_),
    .Y(net181));
 INVx1_ASAP7_75t_R _24007_ (.A(_02536_),
    .Y(_06152_));
 NAND2x1_ASAP7_75t_R _24008_ (.A(_13261_),
    .B(_00233_),
    .Y(_06153_));
 OA211x2_ASAP7_75t_R _24009_ (.A1(_13261_),
    .A2(_06065_),
    .B(_05739_),
    .C(_06153_),
    .Y(_06154_));
 AO21x2_ASAP7_75t_R _24010_ (.A1(_06152_),
    .A2(_06148_),
    .B(_06154_),
    .Y(net182));
 OR3x1_ASAP7_75t_R _24011_ (.A(_13283_),
    .B(_00281_),
    .C(_00235_),
    .Y(_06155_));
 OAI21x1_ASAP7_75t_R _24012_ (.A1(_13261_),
    .A2(net276),
    .B(_06155_),
    .Y(_06156_));
 NAND2x1_ASAP7_75t_R _24013_ (.A(_13283_),
    .B(_02537_),
    .Y(_06157_));
 OA211x2_ASAP7_75t_R _24014_ (.A1(_13283_),
    .A2(_00234_),
    .B(_06148_),
    .C(_06157_),
    .Y(_06158_));
 AO21x2_ASAP7_75t_R _24015_ (.A1(_05739_),
    .A2(_06156_),
    .B(_06158_),
    .Y(net183));
 NAND2x1_ASAP7_75t_R _24016_ (.A(_13261_),
    .B(_00236_),
    .Y(_06159_));
 OA211x2_ASAP7_75t_R _24017_ (.A1(_13261_),
    .A2(_06067_),
    .B(_05739_),
    .C(_06159_),
    .Y(_06160_));
 AO21x2_ASAP7_75t_R _24018_ (.A1(_18336_),
    .A2(_06148_),
    .B(_06160_),
    .Y(net184));
 OR2x2_ASAP7_75t_R _24019_ (.A(_13218_),
    .B(_05730_),
    .Y(_06161_));
 AND2x2_ASAP7_75t_R _24020_ (.A(_00277_),
    .B(_06161_),
    .Y(net185));
 AO32x2_ASAP7_75t_R _24021_ (.A1(_13261_),
    .A2(_13263_),
    .A3(_13267_),
    .B1(_13271_),
    .B2(_13235_),
    .Y(_06162_));
 NAND3x1_ASAP7_75t_R _24022_ (.A(_01713_),
    .B(_14585_),
    .C(_06162_),
    .Y(_06163_));
 OA31x2_ASAP7_75t_R _24023_ (.A1(_14592_),
    .A2(_14624_),
    .A3(_06163_),
    .B1(_01710_),
    .Y(_06164_));
 OR2x6_ASAP7_75t_R _24024_ (.A(_01317_),
    .B(_01721_),
    .Y(_06165_));
 NAND2x1_ASAP7_75t_R _24025_ (.A(_14584_),
    .B(_06165_),
    .Y(_06166_));
 AND3x4_ASAP7_75t_R _24026_ (.A(_01719_),
    .B(_01724_),
    .C(_01725_),
    .Y(_06167_));
 NAND2x1_ASAP7_75t_R _24027_ (.A(_17592_),
    .B(_02140_),
    .Y(_06168_));
 OR3x1_ASAP7_75t_R _24028_ (.A(_02030_),
    .B(_17592_),
    .C(_02140_),
    .Y(_06169_));
 OA21x2_ASAP7_75t_R _24029_ (.A1(_02032_),
    .A2(_06168_),
    .B(_06169_),
    .Y(_06170_));
 AND2x2_ASAP7_75t_R _24030_ (.A(_01311_),
    .B(_06170_),
    .Y(_06171_));
 NOR2x2_ASAP7_75t_R _24031_ (.A(_01317_),
    .B(_01721_),
    .Y(_06172_));
 OR3x1_ASAP7_75t_R _24032_ (.A(net360),
    .B(_13127_),
    .C(_06172_),
    .Y(_06173_));
 INVx4_ASAP7_75t_R _24033_ (.A(_01312_),
    .Y(_06174_));
 NAND2x1_ASAP7_75t_R _24034_ (.A(_01740_),
    .B(_01741_),
    .Y(_06175_));
 OR5x1_ASAP7_75t_R _24035_ (.A(_06174_),
    .B(_06175_),
    .C(_13584_),
    .D(_14596_),
    .E(_05704_),
    .Y(_06176_));
 OR4x2_ASAP7_75t_R _24036_ (.A(_06167_),
    .B(_06171_),
    .C(_06173_),
    .D(_06176_),
    .Y(_06177_));
 NAND2x1_ASAP7_75t_R _24037_ (.A(_05527_),
    .B(_06177_),
    .Y(_06178_));
 AND3x1_ASAP7_75t_R _24038_ (.A(_05705_),
    .B(_05712_),
    .C(_06167_),
    .Y(_06179_));
 INVx1_ASAP7_75t_R _24039_ (.A(_01714_),
    .Y(_06180_));
 NAND2x2_ASAP7_75t_R _24040_ (.A(_01715_),
    .B(_01716_),
    .Y(_06181_));
 BUFx2_ASAP7_75t_R input100 (.A(instr_rdata_i[13]),
    .Y(net100));
 INVx1_ASAP7_75t_R _24042_ (.A(net60),
    .Y(_06183_));
 AND2x2_ASAP7_75t_R _24043_ (.A(_06183_),
    .B(_02034_),
    .Y(_06184_));
 OR2x2_ASAP7_75t_R _24044_ (.A(_01714_),
    .B(_06181_),
    .Y(_06185_));
 AO21x1_ASAP7_75t_R _24045_ (.A1(_01717_),
    .A2(_06184_),
    .B(_06185_),
    .Y(_06186_));
 OA21x2_ASAP7_75t_R _24046_ (.A1(_06180_),
    .A2(_06181_),
    .B(_06186_),
    .Y(_06187_));
 NOR2x1_ASAP7_75t_R _24047_ (.A(_01716_),
    .B(_01717_),
    .Y(_06188_));
 AND3x4_ASAP7_75t_R _24048_ (.A(_01714_),
    .B(_14581_),
    .C(_06188_),
    .Y(_06189_));
 INVx2_ASAP7_75t_R _24049_ (.A(_01453_),
    .Y(_06190_));
 OA211x2_ASAP7_75t_R _24050_ (.A1(net145),
    .A2(_06190_),
    .B(_01718_),
    .C(_01311_),
    .Y(_06191_));
 NAND2x2_ASAP7_75t_R _24051_ (.A(_06189_),
    .B(_06191_),
    .Y(_06192_));
 INVx1_ASAP7_75t_R _24052_ (.A(_01960_),
    .Y(_06193_));
 INVx1_ASAP7_75t_R _24053_ (.A(_01961_),
    .Y(_06194_));
 AO22x2_ASAP7_75t_R _24054_ (.A1(net138),
    .A2(_06193_),
    .B1(_06194_),
    .B2(net137),
    .Y(_06195_));
 INVx1_ASAP7_75t_R _24055_ (.A(_01962_),
    .Y(_06196_));
 INVx1_ASAP7_75t_R _24056_ (.A(_01963_),
    .Y(_06197_));
 AO22x1_ASAP7_75t_R _24057_ (.A1(net136),
    .A2(_06196_),
    .B1(_06197_),
    .B2(net130),
    .Y(_06198_));
 INVx1_ASAP7_75t_R _24058_ (.A(_01956_),
    .Y(_06199_));
 INVx1_ASAP7_75t_R _24059_ (.A(_01957_),
    .Y(_06200_));
 AO22x1_ASAP7_75t_R _24060_ (.A1(net142),
    .A2(_06199_),
    .B1(_06200_),
    .B2(net141),
    .Y(_06201_));
 INVx2_ASAP7_75t_R _24061_ (.A(_01958_),
    .Y(_06202_));
 INVx1_ASAP7_75t_R _24062_ (.A(_01959_),
    .Y(_06203_));
 AO22x1_ASAP7_75t_R _24063_ (.A1(net140),
    .A2(_06202_),
    .B1(_06203_),
    .B2(net139),
    .Y(_06204_));
 OR4x2_ASAP7_75t_R _24064_ (.A(_06195_),
    .B(_06198_),
    .C(_06201_),
    .D(_06204_),
    .Y(_06205_));
 INVx2_ASAP7_75t_R _24065_ (.A(_01949_),
    .Y(_06206_));
 INVx1_ASAP7_75t_R _24066_ (.A(_01951_),
    .Y(_06207_));
 INVx1_ASAP7_75t_R _24067_ (.A(_01950_),
    .Y(_06208_));
 AND2x2_ASAP7_75t_R _24068_ (.A(net134),
    .B(_06208_),
    .Y(_06209_));
 AO221x2_ASAP7_75t_R _24069_ (.A1(net135),
    .A2(_06206_),
    .B1(_06207_),
    .B2(net133),
    .C(_06209_),
    .Y(_06210_));
 INVx2_ASAP7_75t_R _24070_ (.A(_01946_),
    .Y(_06211_));
 INVx1_ASAP7_75t_R _24071_ (.A(_01948_),
    .Y(_06212_));
 AO22x1_ASAP7_75t_R _24072_ (.A1(net146),
    .A2(_06211_),
    .B1(_06212_),
    .B2(net129),
    .Y(_06213_));
 INVx1_ASAP7_75t_R _24073_ (.A(_01947_),
    .Y(_06214_));
 AO21x1_ASAP7_75t_R _24074_ (.A1(net147),
    .A2(_06214_),
    .B(net145),
    .Y(_06215_));
 INVx1_ASAP7_75t_R _24075_ (.A(_01954_),
    .Y(_06216_));
 INVx1_ASAP7_75t_R _24076_ (.A(_01955_),
    .Y(_06217_));
 AO22x1_ASAP7_75t_R _24077_ (.A1(net144),
    .A2(_06216_),
    .B1(_06217_),
    .B2(net143),
    .Y(_06218_));
 INVx1_ASAP7_75t_R _24078_ (.A(_01952_),
    .Y(_06219_));
 INVx1_ASAP7_75t_R _24079_ (.A(_01953_),
    .Y(_06220_));
 AO22x1_ASAP7_75t_R _24080_ (.A1(net132),
    .A2(_06219_),
    .B1(_06220_),
    .B2(net131),
    .Y(_06221_));
 OR4x2_ASAP7_75t_R _24081_ (.A(_06213_),
    .B(_06215_),
    .C(_06218_),
    .D(_06221_),
    .Y(_06222_));
 NOR3x2_ASAP7_75t_R _24082_ (.B(_06210_),
    .C(_06222_),
    .Y(_06223_),
    .A(_06205_));
 OR2x6_ASAP7_75t_R _24083_ (.A(_06192_),
    .B(_06223_),
    .Y(_06224_));
 OA211x2_ASAP7_75t_R _24084_ (.A1(_06178_),
    .A2(_06179_),
    .B(_06187_),
    .C(_06224_),
    .Y(_06225_));
 OA21x2_ASAP7_75t_R _24085_ (.A1(_06164_),
    .A2(_06166_),
    .B(_06225_),
    .Y(_06226_));
 BUFx2_ASAP7_75t_R input99 (.A(instr_rdata_i[12]),
    .Y(net99));
 BUFx2_ASAP7_75t_R input98 (.A(instr_rdata_i[11]),
    .Y(net98));
 BUFx3_ASAP7_75t_R input97 (.A(instr_rdata_i[10]),
    .Y(net97));
 BUFx3_ASAP7_75t_R input96 (.A(instr_rdata_i[0]),
    .Y(net96));
 NOR2x1_ASAP7_75t_R _24090_ (.A(_06218_),
    .B(_06221_),
    .Y(_06231_));
 NOR2x1_ASAP7_75t_R _24091_ (.A(_06205_),
    .B(_06210_),
    .Y(_06232_));
 AND2x2_ASAP7_75t_R _24092_ (.A(_06231_),
    .B(_06232_),
    .Y(_06233_));
 AO21x1_ASAP7_75t_R _24093_ (.A1(net145),
    .A2(_01718_),
    .B(_06233_),
    .Y(_06234_));
 AND2x2_ASAP7_75t_R _24094_ (.A(net132),
    .B(_06219_),
    .Y(_06235_));
 INVx1_ASAP7_75t_R _24095_ (.A(net131),
    .Y(_06236_));
 NAND2x1_ASAP7_75t_R _24096_ (.A(net143),
    .B(_06217_),
    .Y(_06237_));
 NAND2x1_ASAP7_75t_R _24097_ (.A(net141),
    .B(_06200_),
    .Y(_06238_));
 INVx1_ASAP7_75t_R _24098_ (.A(net139),
    .Y(_06239_));
 NAND2x1_ASAP7_75t_R _24099_ (.A(net137),
    .B(_06194_),
    .Y(_06240_));
 AO32x1_ASAP7_75t_R _24100_ (.A1(net136),
    .A2(_06196_),
    .A3(_06240_),
    .B1(net138),
    .B2(_06193_),
    .Y(_06241_));
 OA21x2_ASAP7_75t_R _24101_ (.A1(_06239_),
    .A2(_01959_),
    .B(_06241_),
    .Y(_06242_));
 AO21x1_ASAP7_75t_R _24102_ (.A1(net140),
    .A2(_06202_),
    .B(_06242_),
    .Y(_06243_));
 AO22x1_ASAP7_75t_R _24103_ (.A1(net142),
    .A2(_06199_),
    .B1(_06238_),
    .B2(_06243_),
    .Y(_06244_));
 AO22x1_ASAP7_75t_R _24104_ (.A1(net144),
    .A2(_06216_),
    .B1(_06237_),
    .B2(_06244_),
    .Y(_06245_));
 OA21x2_ASAP7_75t_R _24105_ (.A1(_06236_),
    .A2(_01953_),
    .B(_06245_),
    .Y(_06246_));
 NAND2x1_ASAP7_75t_R _24106_ (.A(net133),
    .B(_06207_),
    .Y(_06247_));
 OA21x2_ASAP7_75t_R _24107_ (.A1(_06235_),
    .A2(_06246_),
    .B(_06247_),
    .Y(_06248_));
 NAND2x1_ASAP7_75t_R _24108_ (.A(net135),
    .B(_06206_),
    .Y(_06249_));
 OA21x2_ASAP7_75t_R _24109_ (.A1(_06209_),
    .A2(_06248_),
    .B(_06249_),
    .Y(_06250_));
 NOR2x2_ASAP7_75t_R _24110_ (.A(_06192_),
    .B(_06223_),
    .Y(_06251_));
 OA21x2_ASAP7_75t_R _24111_ (.A1(_06234_),
    .A2(_06250_),
    .B(_06251_),
    .Y(_06252_));
 INVx1_ASAP7_75t_R _24112_ (.A(_06252_),
    .Y(_06253_));
 OAI21x1_ASAP7_75t_R _24113_ (.A1(_06164_),
    .A2(_06166_),
    .B(_06225_),
    .Y(_06254_));
 BUFx2_ASAP7_75t_R input95 (.A(instr_gnt_i),
    .Y(net95));
 BUFx2_ASAP7_75t_R input94 (.A(instr_err_i),
    .Y(net94));
 NAND2x2_ASAP7_75t_R _24116_ (.A(_05527_),
    .B(_06167_),
    .Y(_06257_));
 OR2x6_ASAP7_75t_R _24117_ (.A(_05705_),
    .B(_06257_),
    .Y(_06258_));
 BUFx2_ASAP7_75t_R input93 (.A(hart_id_i[9]),
    .Y(net93));
 BUFx2_ASAP7_75t_R input92 (.A(hart_id_i[8]),
    .Y(net92));
 BUFx2_ASAP7_75t_R input91 (.A(hart_id_i[7]),
    .Y(net91));
 OR2x6_ASAP7_75t_R _24121_ (.A(_05712_),
    .B(_06257_),
    .Y(_06262_));
 BUFx2_ASAP7_75t_R input90 (.A(hart_id_i[6]),
    .Y(net90));
 BUFx2_ASAP7_75t_R input89 (.A(hart_id_i[5]),
    .Y(net89));
 BUFx2_ASAP7_75t_R input88 (.A(hart_id_i[4]),
    .Y(net88));
 NAND2x2_ASAP7_75t_R _24125_ (.A(_14580_),
    .B(_14583_),
    .Y(_06266_));
 BUFx2_ASAP7_75t_R input87 (.A(hart_id_i[3]),
    .Y(net87));
 BUFx2_ASAP7_75t_R input86 (.A(hart_id_i[31]),
    .Y(net86));
 BUFx2_ASAP7_75t_R input85 (.A(hart_id_i[30]),
    .Y(net85));
 OA222x2_ASAP7_75t_R _24129_ (.A1(_01575_),
    .A2(_06258_),
    .B1(_06262_),
    .B2(_01943_),
    .C1(_06266_),
    .C2(_05767_),
    .Y(_06270_));
 AND3x4_ASAP7_75t_R _24130_ (.A(_06253_),
    .B(_06254_),
    .C(_06270_),
    .Y(_06271_));
 AOI21x1_ASAP7_75t_R _24131_ (.A1(_01549_),
    .A2(net287),
    .B(_06271_),
    .Y(_18387_));
 BUFx2_ASAP7_75t_R input84 (.A(hart_id_i[2]),
    .Y(net84));
 BUFx2_ASAP7_75t_R input83 (.A(hart_id_i[29]),
    .Y(net83));
 BUFx2_ASAP7_75t_R input82 (.A(hart_id_i[28]),
    .Y(net82));
 NOR2x1_ASAP7_75t_R _24135_ (.A(_00237_),
    .B(_02201_),
    .Y(_06275_));
 AO21x1_ASAP7_75t_R _24136_ (.A1(_00237_),
    .A2(_18387_),
    .B(_06275_),
    .Y(net239));
 BUFx2_ASAP7_75t_R input81 (.A(hart_id_i[27]),
    .Y(net81));
 INVx5_ASAP7_75t_R _24138_ (.A(net275),
    .Y(_06277_));
 NAND3x2_ASAP7_75t_R _24139_ (.B(_01724_),
    .C(_01725_),
    .Y(_06278_),
    .A(_01719_));
 NAND2x2_ASAP7_75t_R _24140_ (.A(_05527_),
    .B(_06278_),
    .Y(_06279_));
 OA222x2_ASAP7_75t_R _24141_ (.A1(_06277_),
    .A2(_06266_),
    .B1(_06262_),
    .B2(_01942_),
    .C1(_06279_),
    .C2(_01311_),
    .Y(_06280_));
 INVx1_ASAP7_75t_R _24142_ (.A(net134),
    .Y(_06281_));
 INVx1_ASAP7_75t_R _24143_ (.A(_06218_),
    .Y(_06282_));
 AOI22x1_ASAP7_75t_R _24144_ (.A1(net140),
    .A2(_06202_),
    .B1(_06203_),
    .B2(net139),
    .Y(_06283_));
 AO21x1_ASAP7_75t_R _24145_ (.A1(_06195_),
    .A2(_06283_),
    .B(_06201_),
    .Y(_06284_));
 AO21x1_ASAP7_75t_R _24146_ (.A1(_06282_),
    .A2(_06284_),
    .B(_06221_),
    .Y(_06285_));
 OA211x2_ASAP7_75t_R _24147_ (.A1(_06281_),
    .A2(_01950_),
    .B(_06247_),
    .C(_06285_),
    .Y(_06286_));
 AO21x1_ASAP7_75t_R _24148_ (.A1(net135),
    .A2(_06206_),
    .B(_06234_),
    .Y(_06287_));
 OA21x2_ASAP7_75t_R _24149_ (.A1(_06286_),
    .A2(_06287_),
    .B(_06251_),
    .Y(_06288_));
 INVx1_ASAP7_75t_R _24150_ (.A(_06288_),
    .Y(_06289_));
 OR3x1_ASAP7_75t_R _24151_ (.A(_00081_),
    .B(_05705_),
    .C(_06257_),
    .Y(_06290_));
 AND4x2_ASAP7_75t_R _24152_ (.A(_06254_),
    .B(_06280_),
    .C(_06289_),
    .D(_06290_),
    .Y(_06291_));
 AOI21x1_ASAP7_75t_R _24153_ (.A1(_01548_),
    .A2(net287),
    .B(_06291_),
    .Y(_18357_));
 BUFx2_ASAP7_75t_R input80 (.A(hart_id_i[26]),
    .Y(net80));
 NOR2x1_ASAP7_75t_R _24155_ (.A(_00237_),
    .B(_02200_),
    .Y(_06293_));
 AO21x1_ASAP7_75t_R _24156_ (.A1(_00237_),
    .A2(_18357_),
    .B(_06293_),
    .Y(net242));
 OA22x2_ASAP7_75t_R _24157_ (.A1(_00084_),
    .A2(_05705_),
    .B1(_05712_),
    .B2(_01941_),
    .Y(_06294_));
 NOR3x1_ASAP7_75t_R _24158_ (.A(_06213_),
    .B(_06195_),
    .C(_06198_),
    .Y(_06295_));
 OR3x1_ASAP7_75t_R _24159_ (.A(_06201_),
    .B(_06204_),
    .C(_06295_),
    .Y(_06296_));
 NAND2x1_ASAP7_75t_R _24160_ (.A(_06231_),
    .B(_06296_),
    .Y(_06297_));
 AOI21x1_ASAP7_75t_R _24161_ (.A1(net145),
    .A2(_01718_),
    .B(_06210_),
    .Y(_06298_));
 AO21x2_ASAP7_75t_R _24162_ (.A1(_06297_),
    .A2(_06298_),
    .B(_06224_),
    .Y(_06299_));
 NAND2x1_ASAP7_75t_R _24163_ (.A(_14584_),
    .B(net175),
    .Y(_06300_));
 OA211x2_ASAP7_75t_R _24164_ (.A1(_06257_),
    .A2(_06294_),
    .B(_06299_),
    .C(_06300_),
    .Y(_06301_));
 AND2x2_ASAP7_75t_R _24165_ (.A(_06254_),
    .B(_06301_),
    .Y(_06302_));
 AOI21x1_ASAP7_75t_R _24166_ (.A1(_01547_),
    .A2(net287),
    .B(_06302_),
    .Y(_18359_));
 NOR2x1_ASAP7_75t_R _24167_ (.A(_00237_),
    .B(_02199_),
    .Y(_06303_));
 AO21x1_ASAP7_75t_R _24168_ (.A1(_00237_),
    .A2(_18359_),
    .B(_06303_),
    .Y(net243));
 AND2x4_ASAP7_75t_R _24169_ (.A(_05527_),
    .B(_06167_),
    .Y(_06304_));
 OAI22x1_ASAP7_75t_R _24170_ (.A1(_00087_),
    .A2(_05705_),
    .B1(_05712_),
    .B2(_01940_),
    .Y(_06305_));
 NAND2x1_ASAP7_75t_R _24171_ (.A(net129),
    .B(_06212_),
    .Y(_06306_));
 OA211x2_ASAP7_75t_R _24172_ (.A1(_06306_),
    .A2(_06205_),
    .B(_06231_),
    .C(_06298_),
    .Y(_06307_));
 NOR2x2_ASAP7_75t_R _24173_ (.A(_06224_),
    .B(_06307_),
    .Y(_06308_));
 AO221x2_ASAP7_75t_R _24174_ (.A1(net176),
    .A2(_14584_),
    .B1(_06304_),
    .B2(_06305_),
    .C(_06308_),
    .Y(_06309_));
 NOR2x2_ASAP7_75t_R _24175_ (.A(net287),
    .B(_06309_),
    .Y(_06310_));
 AO21x1_ASAP7_75t_R _24176_ (.A1(_01546_),
    .A2(net287),
    .B(_06310_),
    .Y(_06311_));
 CKINVDCx5p33_ASAP7_75t_R _24177_ (.A(_00237_),
    .Y(_06312_));
 BUFx2_ASAP7_75t_R input79 (.A(hart_id_i[25]),
    .Y(net79));
 AND2x2_ASAP7_75t_R _24179_ (.A(_06312_),
    .B(_02198_),
    .Y(_06314_));
 AOI21x1_ASAP7_75t_R _24180_ (.A1(_00237_),
    .A2(_06311_),
    .B(_06314_),
    .Y(net244));
 OAI22x1_ASAP7_75t_R _24181_ (.A1(_00090_),
    .A2(_05705_),
    .B1(_05712_),
    .B2(_01939_),
    .Y(_06315_));
 NAND2x1_ASAP7_75t_R _24182_ (.A(_06304_),
    .B(_06315_),
    .Y(_06316_));
 INVx1_ASAP7_75t_R _24183_ (.A(net145),
    .Y(_06317_));
 AO21x2_ASAP7_75t_R _24184_ (.A1(_06317_),
    .A2(_06233_),
    .B(_06192_),
    .Y(_06318_));
 OA211x2_ASAP7_75t_R _24185_ (.A1(_06266_),
    .A2(_05768_),
    .B(_06316_),
    .C(_06318_),
    .Y(_06319_));
 AND2x2_ASAP7_75t_R _24186_ (.A(_06254_),
    .B(_06319_),
    .Y(_06320_));
 AOI21x1_ASAP7_75t_R _24187_ (.A1(_01545_),
    .A2(net287),
    .B(_06320_),
    .Y(_18361_));
 BUFx2_ASAP7_75t_R input78 (.A(hart_id_i[24]),
    .Y(net78));
 NOR2x1_ASAP7_75t_R _24189_ (.A(_00237_),
    .B(_02197_),
    .Y(_06322_));
 AO21x1_ASAP7_75t_R _24190_ (.A1(_00237_),
    .A2(_18361_),
    .B(_06322_),
    .Y(net245));
 NOR2x2_ASAP7_75t_R _24191_ (.A(_14601_),
    .B(_05704_),
    .Y(_06323_));
 AND2x2_ASAP7_75t_R _24192_ (.A(_01714_),
    .B(_14581_),
    .Y(_06324_));
 AO21x1_ASAP7_75t_R _24193_ (.A1(_05526_),
    .A2(_06278_),
    .B(_14580_),
    .Y(_06325_));
 BUFx2_ASAP7_75t_R input77 (.A(hart_id_i[23]),
    .Y(net77));
 NOR2x2_ASAP7_75t_R _24195_ (.A(_01714_),
    .B(_06181_),
    .Y(_06327_));
 AO21x1_ASAP7_75t_R _24196_ (.A1(_06324_),
    .A2(_06325_),
    .B(_06327_),
    .Y(_06328_));
 AO21x2_ASAP7_75t_R _24197_ (.A1(_06304_),
    .A2(_06323_),
    .B(_06328_),
    .Y(_06329_));
 BUFx2_ASAP7_75t_R input76 (.A(hart_id_i[22]),
    .Y(net76));
 OA22x2_ASAP7_75t_R _24199_ (.A1(_01574_),
    .A2(_06258_),
    .B1(_06262_),
    .B2(_01938_),
    .Y(_06331_));
 OA211x2_ASAP7_75t_R _24200_ (.A1(_00676_),
    .A2(_06266_),
    .B(_06329_),
    .C(_06331_),
    .Y(_06332_));
 AND2x2_ASAP7_75t_R _24201_ (.A(_06254_),
    .B(_06332_),
    .Y(_06333_));
 AO21x1_ASAP7_75t_R _24202_ (.A1(_01544_),
    .A2(net287),
    .B(_06333_),
    .Y(_06334_));
 AND2x2_ASAP7_75t_R _24203_ (.A(_06312_),
    .B(_02196_),
    .Y(_06335_));
 AOI21x1_ASAP7_75t_R _24204_ (.A1(_00237_),
    .A2(_06334_),
    .B(_06335_),
    .Y(net246));
 INVx1_ASAP7_75t_R _24205_ (.A(_01543_),
    .Y(_06336_));
 BUFx2_ASAP7_75t_R input75 (.A(hart_id_i[21]),
    .Y(net75));
 INVx1_ASAP7_75t_R _24207_ (.A(net23),
    .Y(_06338_));
 AOI21x1_ASAP7_75t_R _24208_ (.A1(_06304_),
    .A2(_06323_),
    .B(_06328_),
    .Y(_06339_));
 AND2x6_ASAP7_75t_R _24209_ (.A(_05527_),
    .B(_06278_),
    .Y(_06340_));
 AOI21x1_ASAP7_75t_R _24210_ (.A1(_01311_),
    .A2(_06340_),
    .B(_06189_),
    .Y(_06341_));
 OA22x2_ASAP7_75t_R _24211_ (.A1(_06266_),
    .A2(_05773_),
    .B1(_06341_),
    .B2(_00095_),
    .Y(_06342_));
 OA22x2_ASAP7_75t_R _24212_ (.A1(_01937_),
    .A2(_14596_),
    .B1(_14599_),
    .B2(_01573_),
    .Y(_06343_));
 OR4x1_ASAP7_75t_R _24213_ (.A(_14600_),
    .B(_05704_),
    .C(_06257_),
    .D(_06343_),
    .Y(_06344_));
 AND3x1_ASAP7_75t_R _24214_ (.A(_06329_),
    .B(_06342_),
    .C(_06344_),
    .Y(_06345_));
 AO21x1_ASAP7_75t_R _24215_ (.A1(_06338_),
    .A2(_06339_),
    .B(_06345_),
    .Y(_06346_));
 NOR2x1_ASAP7_75t_R _24216_ (.A(net287),
    .B(_06346_),
    .Y(_06347_));
 AO21x1_ASAP7_75t_R _24217_ (.A1(_06336_),
    .A2(net287),
    .B(_06347_),
    .Y(_18363_));
 NAND2x1_ASAP7_75t_R _24218_ (.A(_06312_),
    .B(_02195_),
    .Y(_06348_));
 OA21x2_ASAP7_75t_R _24219_ (.A1(_06312_),
    .A2(_18363_),
    .B(_06348_),
    .Y(net247));
 INVx1_ASAP7_75t_R _24220_ (.A(_02194_),
    .Y(_06349_));
 INVx4_ASAP7_75t_R _24221_ (.A(net180),
    .Y(_06350_));
 OA22x2_ASAP7_75t_R _24222_ (.A1(_01572_),
    .A2(_05705_),
    .B1(_05712_),
    .B2(_01936_),
    .Y(_06351_));
 OA222x2_ASAP7_75t_R _24223_ (.A1(_06350_),
    .A2(_06266_),
    .B1(_06257_),
    .B2(_06351_),
    .C1(_06341_),
    .C2(_00098_),
    .Y(_06352_));
 NOR2x1_ASAP7_75t_R _24224_ (.A(net24),
    .B(_06329_),
    .Y(_06353_));
 AO21x2_ASAP7_75t_R _24225_ (.A1(_06329_),
    .A2(_06352_),
    .B(_06353_),
    .Y(_06354_));
 NOR2x1_ASAP7_75t_R _24226_ (.A(net287),
    .B(_06354_),
    .Y(_06355_));
 BUFx2_ASAP7_75t_R input74 (.A(hart_id_i[20]),
    .Y(net74));
 NOR2x1_ASAP7_75t_R _24228_ (.A(_01542_),
    .B(_06254_),
    .Y(_06357_));
 OR3x1_ASAP7_75t_R _24229_ (.A(_06312_),
    .B(_06355_),
    .C(_06357_),
    .Y(_06358_));
 OA21x2_ASAP7_75t_R _24230_ (.A1(_00237_),
    .A2(_06349_),
    .B(_06358_),
    .Y(net248));
 OAI22x1_ASAP7_75t_R _24231_ (.A1(_01571_),
    .A2(_05705_),
    .B1(_05712_),
    .B2(_01935_),
    .Y(_06359_));
 OAI22x1_ASAP7_75t_R _24232_ (.A1(_06266_),
    .A2(_05772_),
    .B1(_06341_),
    .B2(_00101_),
    .Y(_06360_));
 AO21x1_ASAP7_75t_R _24233_ (.A1(_06304_),
    .A2(_06359_),
    .B(_06360_),
    .Y(_06361_));
 AOI211x1_ASAP7_75t_R _24234_ (.A1(net1),
    .A2(_06339_),
    .B(_06361_),
    .C(net287),
    .Y(_06362_));
 AOI21x1_ASAP7_75t_R _24235_ (.A1(_01541_),
    .A2(net287),
    .B(_06362_),
    .Y(_18365_));
 NOR2x1_ASAP7_75t_R _24236_ (.A(_00237_),
    .B(_02193_),
    .Y(_06363_));
 AO21x1_ASAP7_75t_R _24237_ (.A1(_00237_),
    .A2(_18365_),
    .B(_06363_),
    .Y(net219));
 BUFx2_ASAP7_75t_R input73 (.A(hart_id_i[1]),
    .Y(net73));
 NOR2x1_ASAP7_75t_R _24239_ (.A(net2),
    .B(_06329_),
    .Y(_06365_));
 OAI22x1_ASAP7_75t_R _24240_ (.A1(_01570_),
    .A2(_05705_),
    .B1(_05712_),
    .B2(_01934_),
    .Y(_06366_));
 NAND2x1_ASAP7_75t_R _24241_ (.A(_06304_),
    .B(_06366_),
    .Y(_06367_));
 INVx4_ASAP7_75t_R _24242_ (.A(net152),
    .Y(_06368_));
 OR4x1_ASAP7_75t_R _24243_ (.A(_06368_),
    .B(_06180_),
    .C(_01715_),
    .D(_01717_),
    .Y(_06369_));
 OA21x2_ASAP7_75t_R _24244_ (.A1(_01714_),
    .A2(_14581_),
    .B(_06369_),
    .Y(_06370_));
 NOR2x1_ASAP7_75t_R _24245_ (.A(_06189_),
    .B(_06340_),
    .Y(_06371_));
 OA21x2_ASAP7_75t_R _24246_ (.A1(_01311_),
    .A2(_06279_),
    .B(_00657_),
    .Y(_06372_));
 OA22x2_ASAP7_75t_R _24247_ (.A1(_05526_),
    .A2(_06370_),
    .B1(_06371_),
    .B2(_06372_),
    .Y(_06373_));
 AND3x1_ASAP7_75t_R _24248_ (.A(_06329_),
    .B(_06367_),
    .C(_06373_),
    .Y(_06374_));
 OR3x2_ASAP7_75t_R _24249_ (.A(net287),
    .B(_06365_),
    .C(_06374_),
    .Y(_06375_));
 OA21x2_ASAP7_75t_R _24250_ (.A1(_01540_),
    .A2(_06254_),
    .B(_06375_),
    .Y(_06376_));
 AND2x2_ASAP7_75t_R _24251_ (.A(_06312_),
    .B(_02192_),
    .Y(_06377_));
 AOI21x1_ASAP7_75t_R _24252_ (.A1(_00237_),
    .A2(_06376_),
    .B(_06377_),
    .Y(net220));
 NAND2x1_ASAP7_75t_R _24253_ (.A(net3),
    .B(_06339_),
    .Y(_06378_));
 OA222x2_ASAP7_75t_R _24254_ (.A1(_06266_),
    .A2(_05771_),
    .B1(_06262_),
    .B2(_01933_),
    .C1(_00656_),
    .C2(_06341_),
    .Y(_06379_));
 OA211x2_ASAP7_75t_R _24255_ (.A1(_01569_),
    .A2(_06258_),
    .B(_06378_),
    .C(_06379_),
    .Y(_06380_));
 AND2x2_ASAP7_75t_R _24256_ (.A(_06254_),
    .B(_06380_),
    .Y(_06381_));
 AOI21x1_ASAP7_75t_R _24257_ (.A1(_01539_),
    .A2(net287),
    .B(_06381_),
    .Y(_18366_));
 NOR2x1_ASAP7_75t_R _24258_ (.A(net415),
    .B(_02191_),
    .Y(_06382_));
 AO21x1_ASAP7_75t_R _24259_ (.A1(_00237_),
    .A2(_18366_),
    .B(_06382_),
    .Y(net221));
 INVx1_ASAP7_75t_R _24260_ (.A(_02190_),
    .Y(_06383_));
 INVx5_ASAP7_75t_R _24261_ (.A(net154),
    .Y(_06384_));
 OA22x2_ASAP7_75t_R _24262_ (.A1(_01568_),
    .A2(_05705_),
    .B1(_05712_),
    .B2(_01932_),
    .Y(_06385_));
 OA222x2_ASAP7_75t_R _24263_ (.A1(_06384_),
    .A2(_06266_),
    .B1(_06257_),
    .B2(_06385_),
    .C1(_06341_),
    .C2(_00108_),
    .Y(_06386_));
 NOR2x1_ASAP7_75t_R _24264_ (.A(net4),
    .B(_06329_),
    .Y(_06387_));
 AO21x2_ASAP7_75t_R _24265_ (.A1(_06329_),
    .A2(_06386_),
    .B(_06387_),
    .Y(_06388_));
 NOR2x1_ASAP7_75t_R _24266_ (.A(net287),
    .B(_06388_),
    .Y(_06389_));
 NOR2x1_ASAP7_75t_R _24267_ (.A(_01538_),
    .B(_06254_),
    .Y(_06390_));
 OR3x1_ASAP7_75t_R _24268_ (.A(_06312_),
    .B(_06389_),
    .C(_06390_),
    .Y(_06391_));
 OA21x2_ASAP7_75t_R _24269_ (.A1(net415),
    .A2(_06383_),
    .B(_06391_),
    .Y(net222));
 OA222x2_ASAP7_75t_R _24270_ (.A1(_06266_),
    .A2(_15557_),
    .B1(_06262_),
    .B2(_01931_),
    .C1(_00111_),
    .C2(_06341_),
    .Y(_06392_));
 OAI21x1_ASAP7_75t_R _24271_ (.A1(_01567_),
    .A2(_06258_),
    .B(_06392_),
    .Y(_06393_));
 AO21x2_ASAP7_75t_R _24272_ (.A1(net5),
    .A2(_06339_),
    .B(_06393_),
    .Y(_06394_));
 NOR2x2_ASAP7_75t_R _24273_ (.A(net287),
    .B(_06394_),
    .Y(_06395_));
 AOI21x1_ASAP7_75t_R _24274_ (.A1(_01537_),
    .A2(net287),
    .B(_06395_),
    .Y(_18368_));
 NOR2x1_ASAP7_75t_R _24275_ (.A(net415),
    .B(_02189_),
    .Y(_06396_));
 AO21x1_ASAP7_75t_R _24276_ (.A1(net415),
    .A2(_18368_),
    .B(_06396_),
    .Y(net223));
 OA222x2_ASAP7_75t_R _24277_ (.A1(net256),
    .A2(_06266_),
    .B1(_06262_),
    .B2(_01930_),
    .C1(_06341_),
    .C2(_00114_),
    .Y(_06397_));
 OAI21x1_ASAP7_75t_R _24278_ (.A1(_01566_),
    .A2(_06258_),
    .B(_06397_),
    .Y(_06398_));
 AO21x1_ASAP7_75t_R _24279_ (.A1(net6),
    .A2(_06339_),
    .B(_06398_),
    .Y(_06399_));
 NOR2x1_ASAP7_75t_R _24280_ (.A(net286),
    .B(_06399_),
    .Y(_06400_));
 AO21x1_ASAP7_75t_R _24281_ (.A1(_01536_),
    .A2(net286),
    .B(_06400_),
    .Y(_06401_));
 AND2x2_ASAP7_75t_R _24282_ (.A(_06312_),
    .B(_02188_),
    .Y(_06402_));
 AOI21x1_ASAP7_75t_R _24283_ (.A1(net415),
    .A2(_06401_),
    .B(_06402_),
    .Y(net224));
 INVx1_ASAP7_75t_R _24284_ (.A(net7),
    .Y(_06403_));
 AND2x4_ASAP7_75t_R _24285_ (.A(_06185_),
    .B(_06371_),
    .Y(_06404_));
 OA21x2_ASAP7_75t_R _24286_ (.A1(_01311_),
    .A2(_06279_),
    .B(_06185_),
    .Y(_06405_));
 AND2x2_ASAP7_75t_R _24287_ (.A(_00117_),
    .B(_06405_),
    .Y(_06406_));
 OA222x2_ASAP7_75t_R _24288_ (.A1(_06266_),
    .A2(_05770_),
    .B1(_06404_),
    .B2(_06406_),
    .C1(_06258_),
    .C2(_01565_),
    .Y(_06407_));
 OA21x2_ASAP7_75t_R _24289_ (.A1(_01929_),
    .A2(_06262_),
    .B(_06407_),
    .Y(_06408_));
 OA211x2_ASAP7_75t_R _24290_ (.A1(_06403_),
    .A2(_06329_),
    .B(_06408_),
    .C(_06254_),
    .Y(_06409_));
 AOI21x1_ASAP7_75t_R _24291_ (.A1(_01535_),
    .A2(net286),
    .B(_06409_),
    .Y(_18370_));
 NOR2x1_ASAP7_75t_R _24292_ (.A(net415),
    .B(_02187_),
    .Y(_06410_));
 AO21x1_ASAP7_75t_R _24293_ (.A1(net415),
    .A2(_18370_),
    .B(_06410_),
    .Y(net225));
 INVx1_ASAP7_75t_R _24294_ (.A(net8),
    .Y(_06411_));
 CKINVDCx5p33_ASAP7_75t_R _24295_ (.A(net158),
    .Y(_06412_));
 OA222x2_ASAP7_75t_R _24296_ (.A1(_06412_),
    .A2(_06266_),
    .B1(_06262_),
    .B2(_01928_),
    .C1(_06341_),
    .C2(_00120_),
    .Y(_06413_));
 OA21x2_ASAP7_75t_R _24297_ (.A1(_01564_),
    .A2(_06258_),
    .B(_06413_),
    .Y(_06414_));
 OA211x2_ASAP7_75t_R _24298_ (.A1(_06411_),
    .A2(_06329_),
    .B(_06414_),
    .C(_06254_),
    .Y(_06415_));
 AO21x1_ASAP7_75t_R _24299_ (.A1(_01534_),
    .A2(net286),
    .B(_06415_),
    .Y(_06416_));
 INVx1_ASAP7_75t_R _24300_ (.A(_06416_),
    .Y(_06417_));
 NOR2x1_ASAP7_75t_R _24301_ (.A(net415),
    .B(_02186_),
    .Y(_06418_));
 AO21x1_ASAP7_75t_R _24302_ (.A1(net415),
    .A2(_06417_),
    .B(_06418_),
    .Y(net226));
 BUFx2_ASAP7_75t_R input72 (.A(hart_id_i[19]),
    .Y(net72));
 OA222x2_ASAP7_75t_R _24304_ (.A1(_06266_),
    .A2(_16020_),
    .B1(_06262_),
    .B2(_01927_),
    .C1(_00123_),
    .C2(_06341_),
    .Y(_06420_));
 OAI21x1_ASAP7_75t_R _24305_ (.A1(_01563_),
    .A2(_06258_),
    .B(_06420_),
    .Y(_06421_));
 AO21x1_ASAP7_75t_R _24306_ (.A1(net9),
    .A2(_06339_),
    .B(_06421_),
    .Y(_06422_));
 NAND2x1_ASAP7_75t_R _24307_ (.A(_01533_),
    .B(net286),
    .Y(_06423_));
 OA21x2_ASAP7_75t_R _24308_ (.A1(net286),
    .A2(_06422_),
    .B(_06423_),
    .Y(_18372_));
 NOR2x1_ASAP7_75t_R _24309_ (.A(net415),
    .B(_02185_),
    .Y(_06424_));
 AO21x1_ASAP7_75t_R _24310_ (.A1(net415),
    .A2(_18372_),
    .B(_06424_),
    .Y(net227));
 INVx1_ASAP7_75t_R _24311_ (.A(net10),
    .Y(_06425_));
 INVx4_ASAP7_75t_R _24312_ (.A(net160),
    .Y(_06426_));
 OA222x2_ASAP7_75t_R _24313_ (.A1(_06426_),
    .A2(_06266_),
    .B1(_06262_),
    .B2(_01926_),
    .C1(_06341_),
    .C2(_00126_),
    .Y(_06427_));
 OA21x2_ASAP7_75t_R _24314_ (.A1(_01562_),
    .A2(_06258_),
    .B(_06427_),
    .Y(_06428_));
 OA211x2_ASAP7_75t_R _24315_ (.A1(_06425_),
    .A2(_06329_),
    .B(_06428_),
    .C(_06254_),
    .Y(_06429_));
 AOI21x1_ASAP7_75t_R _24316_ (.A1(_01532_),
    .A2(net286),
    .B(_06429_),
    .Y(_06430_));
 NOR2x1_ASAP7_75t_R _24317_ (.A(net415),
    .B(_02184_),
    .Y(_06431_));
 AO21x1_ASAP7_75t_R _24318_ (.A1(net415),
    .A2(_06430_),
    .B(_06431_),
    .Y(net228));
 INVx1_ASAP7_75t_R _24319_ (.A(net11),
    .Y(_06432_));
 AND2x2_ASAP7_75t_R _24320_ (.A(_00129_),
    .B(_06405_),
    .Y(_06433_));
 OA222x2_ASAP7_75t_R _24321_ (.A1(_06266_),
    .A2(_16260_),
    .B1(_06404_),
    .B2(_06433_),
    .C1(_06258_),
    .C2(_01561_),
    .Y(_06434_));
 OA21x2_ASAP7_75t_R _24322_ (.A1(_01925_),
    .A2(_06262_),
    .B(_06434_),
    .Y(_06435_));
 OA211x2_ASAP7_75t_R _24323_ (.A1(_06432_),
    .A2(_06329_),
    .B(_06435_),
    .C(_06254_),
    .Y(_06436_));
 AOI21x1_ASAP7_75t_R _24324_ (.A1(_01531_),
    .A2(net286),
    .B(_06436_),
    .Y(_18374_));
 BUFx2_ASAP7_75t_R input71 (.A(hart_id_i[18]),
    .Y(net71));
 NOR2x1_ASAP7_75t_R _24326_ (.A(net415),
    .B(_02183_),
    .Y(_06438_));
 AO21x1_ASAP7_75t_R _24327_ (.A1(net415),
    .A2(_18374_),
    .B(_06438_),
    .Y(net229));
 INVx1_ASAP7_75t_R _24328_ (.A(net12),
    .Y(_06439_));
 INVx4_ASAP7_75t_R _24329_ (.A(net162),
    .Y(_06440_));
 OA222x2_ASAP7_75t_R _24330_ (.A1(_06440_),
    .A2(_06266_),
    .B1(_06262_),
    .B2(_01924_),
    .C1(_06341_),
    .C2(_00132_),
    .Y(_06441_));
 OA21x2_ASAP7_75t_R _24331_ (.A1(_01560_),
    .A2(_06258_),
    .B(_06441_),
    .Y(_06442_));
 OA211x2_ASAP7_75t_R _24332_ (.A1(_06439_),
    .A2(_06329_),
    .B(_06442_),
    .C(_06254_),
    .Y(_06443_));
 AOI21x1_ASAP7_75t_R _24333_ (.A1(_01530_),
    .A2(net286),
    .B(_06443_),
    .Y(_06444_));
 NOR2x1_ASAP7_75t_R _24334_ (.A(net415),
    .B(_02182_),
    .Y(_06445_));
 AO21x1_ASAP7_75t_R _24335_ (.A1(net415),
    .A2(_06444_),
    .B(_06445_),
    .Y(net230));
 INVx1_ASAP7_75t_R _24336_ (.A(net13),
    .Y(_06446_));
 OA222x2_ASAP7_75t_R _24337_ (.A1(_06266_),
    .A2(_05760_),
    .B1(_06262_),
    .B2(_01923_),
    .C1(_00135_),
    .C2(_06341_),
    .Y(_06447_));
 OA21x2_ASAP7_75t_R _24338_ (.A1(_01559_),
    .A2(_06258_),
    .B(_06447_),
    .Y(_06448_));
 OA211x2_ASAP7_75t_R _24339_ (.A1(_06446_),
    .A2(_06329_),
    .B(_06448_),
    .C(_06254_),
    .Y(_06449_));
 AOI21x1_ASAP7_75t_R _24340_ (.A1(_01529_),
    .A2(net286),
    .B(_06449_),
    .Y(_18376_));
 NOR2x1_ASAP7_75t_R _24341_ (.A(net415),
    .B(_02181_),
    .Y(_06450_));
 AO21x1_ASAP7_75t_R _24342_ (.A1(net415),
    .A2(_18376_),
    .B(_06450_),
    .Y(net231));
 INVx1_ASAP7_75t_R _24343_ (.A(net14),
    .Y(_06451_));
 INVx4_ASAP7_75t_R _24344_ (.A(net164),
    .Y(_06452_));
 OA222x2_ASAP7_75t_R _24345_ (.A1(_06452_),
    .A2(_06266_),
    .B1(_06262_),
    .B2(_01922_),
    .C1(_06341_),
    .C2(_00138_),
    .Y(_06453_));
 OA21x2_ASAP7_75t_R _24346_ (.A1(_01558_),
    .A2(_06258_),
    .B(_06453_),
    .Y(_06454_));
 OA211x2_ASAP7_75t_R _24347_ (.A1(_06451_),
    .A2(_06329_),
    .B(_06454_),
    .C(_06254_),
    .Y(_06455_));
 AOI21x1_ASAP7_75t_R _24348_ (.A1(_01528_),
    .A2(net286),
    .B(_06455_),
    .Y(_06456_));
 NOR2x1_ASAP7_75t_R _24349_ (.A(net415),
    .B(_02180_),
    .Y(_06457_));
 AO21x1_ASAP7_75t_R _24350_ (.A1(net415),
    .A2(_06456_),
    .B(_06457_),
    .Y(net232));
 INVx1_ASAP7_75t_R _24351_ (.A(net15),
    .Y(_06458_));
 OA222x2_ASAP7_75t_R _24352_ (.A1(_06266_),
    .A2(_04719_),
    .B1(_06262_),
    .B2(_01921_),
    .C1(_00141_),
    .C2(_06341_),
    .Y(_06459_));
 OA21x2_ASAP7_75t_R _24353_ (.A1(_01557_),
    .A2(_06258_),
    .B(_06459_),
    .Y(_06460_));
 OA211x2_ASAP7_75t_R _24354_ (.A1(_06458_),
    .A2(_06329_),
    .B(_06460_),
    .C(_06254_),
    .Y(_06461_));
 AOI21x1_ASAP7_75t_R _24355_ (.A1(_01527_),
    .A2(net286),
    .B(_06461_),
    .Y(_18378_));
 NOR2x1_ASAP7_75t_R _24356_ (.A(net415),
    .B(_02179_),
    .Y(_06462_));
 AO21x1_ASAP7_75t_R _24357_ (.A1(net415),
    .A2(_18378_),
    .B(_06462_),
    .Y(net233));
 INVx1_ASAP7_75t_R _24358_ (.A(net16),
    .Y(_06463_));
 INVx4_ASAP7_75t_R _24359_ (.A(net166),
    .Y(_06464_));
 AND2x2_ASAP7_75t_R _24360_ (.A(_00144_),
    .B(_06405_),
    .Y(_06465_));
 OA222x2_ASAP7_75t_R _24361_ (.A1(_06464_),
    .A2(_06266_),
    .B1(_06404_),
    .B2(_06465_),
    .C1(_06258_),
    .C2(_01556_),
    .Y(_06466_));
 OA21x2_ASAP7_75t_R _24362_ (.A1(_01920_),
    .A2(_06262_),
    .B(_06466_),
    .Y(_06467_));
 OA211x2_ASAP7_75t_R _24363_ (.A1(_06463_),
    .A2(_06329_),
    .B(_06467_),
    .C(_06254_),
    .Y(_06468_));
 AOI21x1_ASAP7_75t_R _24364_ (.A1(_01526_),
    .A2(net286),
    .B(_06468_),
    .Y(_06469_));
 NOR2x1_ASAP7_75t_R _24365_ (.A(net415),
    .B(_02178_),
    .Y(_06470_));
 AO21x1_ASAP7_75t_R _24366_ (.A1(net415),
    .A2(_06469_),
    .B(_06470_),
    .Y(net234));
 INVx1_ASAP7_75t_R _24367_ (.A(net17),
    .Y(_06471_));
 OA222x2_ASAP7_75t_R _24368_ (.A1(_06266_),
    .A2(_04937_),
    .B1(_06262_),
    .B2(_01919_),
    .C1(_00147_),
    .C2(_06341_),
    .Y(_06472_));
 OA21x2_ASAP7_75t_R _24369_ (.A1(_01555_),
    .A2(_06258_),
    .B(_06472_),
    .Y(_06473_));
 OA211x2_ASAP7_75t_R _24370_ (.A1(_06471_),
    .A2(_06329_),
    .B(_06473_),
    .C(_06254_),
    .Y(_06474_));
 AOI21x1_ASAP7_75t_R _24371_ (.A1(_01525_),
    .A2(net286),
    .B(_06474_),
    .Y(_18380_));
 NOR2x1_ASAP7_75t_R _24372_ (.A(net415),
    .B(_02177_),
    .Y(_06475_));
 AO21x1_ASAP7_75t_R _24373_ (.A1(net415),
    .A2(_18380_),
    .B(_06475_),
    .Y(net235));
 INVx1_ASAP7_75t_R _24374_ (.A(net18),
    .Y(_06476_));
 INVx4_ASAP7_75t_R _24375_ (.A(net168),
    .Y(_06477_));
 AND2x2_ASAP7_75t_R _24376_ (.A(_00150_),
    .B(_06405_),
    .Y(_06478_));
 OA222x2_ASAP7_75t_R _24377_ (.A1(_06477_),
    .A2(_06266_),
    .B1(_06404_),
    .B2(_06478_),
    .C1(_06258_),
    .C2(_01554_),
    .Y(_06479_));
 OA21x2_ASAP7_75t_R _24378_ (.A1(_01918_),
    .A2(_06262_),
    .B(_06479_),
    .Y(_06480_));
 OA211x2_ASAP7_75t_R _24379_ (.A1(_06476_),
    .A2(_06329_),
    .B(_06480_),
    .C(_06254_),
    .Y(_06481_));
 AOI21x1_ASAP7_75t_R _24380_ (.A1(_01524_),
    .A2(net286),
    .B(_06481_),
    .Y(_06482_));
 NOR2x1_ASAP7_75t_R _24381_ (.A(net415),
    .B(_02176_),
    .Y(_06483_));
 AO21x1_ASAP7_75t_R _24382_ (.A1(net415),
    .A2(_06482_),
    .B(_06483_),
    .Y(net236));
 INVx1_ASAP7_75t_R _24383_ (.A(net19),
    .Y(_06484_));
 AND2x2_ASAP7_75t_R _24384_ (.A(_00153_),
    .B(_06405_),
    .Y(_06485_));
 OA222x2_ASAP7_75t_R _24385_ (.A1(_06266_),
    .A2(_05154_),
    .B1(_06404_),
    .B2(_06485_),
    .C1(_06258_),
    .C2(_01553_),
    .Y(_06486_));
 OA21x2_ASAP7_75t_R _24386_ (.A1(_01917_),
    .A2(_06262_),
    .B(_06486_),
    .Y(_06487_));
 OA211x2_ASAP7_75t_R _24387_ (.A1(_06484_),
    .A2(_06329_),
    .B(_06487_),
    .C(_06254_),
    .Y(_06488_));
 AOI21x1_ASAP7_75t_R _24388_ (.A1(_01523_),
    .A2(net286),
    .B(_06488_),
    .Y(_18382_));
 NOR2x1_ASAP7_75t_R _24389_ (.A(net415),
    .B(_02175_),
    .Y(_06489_));
 AO21x1_ASAP7_75t_R _24390_ (.A1(net415),
    .A2(_18382_),
    .B(_06489_),
    .Y(net237));
 INVx1_ASAP7_75t_R _24391_ (.A(net20),
    .Y(_06490_));
 INVx4_ASAP7_75t_R _24392_ (.A(net2118),
    .Y(_06491_));
 OA222x2_ASAP7_75t_R _24393_ (.A1(_06491_),
    .A2(_06266_),
    .B1(_06262_),
    .B2(_01916_),
    .C1(_06341_),
    .C2(_00156_),
    .Y(_06492_));
 OA21x2_ASAP7_75t_R _24394_ (.A1(_01552_),
    .A2(_06258_),
    .B(_06492_),
    .Y(_06493_));
 OA211x2_ASAP7_75t_R _24395_ (.A1(_06490_),
    .A2(_06329_),
    .B(_06493_),
    .C(_06254_),
    .Y(_06494_));
 AOI21x1_ASAP7_75t_R _24396_ (.A1(_01522_),
    .A2(net286),
    .B(_06494_),
    .Y(_06495_));
 NOR2x1_ASAP7_75t_R _24397_ (.A(net415),
    .B(_02174_),
    .Y(_06496_));
 AO21x1_ASAP7_75t_R _24398_ (.A1(net415),
    .A2(_06495_),
    .B(_06496_),
    .Y(net238));
 INVx1_ASAP7_75t_R _24399_ (.A(net21),
    .Y(_06497_));
 OA222x2_ASAP7_75t_R _24400_ (.A1(_06266_),
    .A2(_05372_),
    .B1(_06262_),
    .B2(_01915_),
    .C1(_00159_),
    .C2(_06341_),
    .Y(_06498_));
 OA21x2_ASAP7_75t_R _24401_ (.A1(_01551_),
    .A2(_06258_),
    .B(_06498_),
    .Y(_06499_));
 OA211x2_ASAP7_75t_R _24402_ (.A1(_06497_),
    .A2(_06329_),
    .B(_06499_),
    .C(_06254_),
    .Y(_06500_));
 AOI21x1_ASAP7_75t_R _24403_ (.A1(_01521_),
    .A2(net286),
    .B(_06500_),
    .Y(_18384_));
 NOR2x1_ASAP7_75t_R _24404_ (.A(net415),
    .B(_02173_),
    .Y(_06501_));
 AO21x1_ASAP7_75t_R _24405_ (.A1(net415),
    .A2(_18384_),
    .B(_06501_),
    .Y(net240));
 NAND2x1_ASAP7_75t_R _24406_ (.A(net22),
    .B(_06339_),
    .Y(_06502_));
 OA222x2_ASAP7_75t_R _24407_ (.A1(_01550_),
    .A2(_06258_),
    .B1(_06262_),
    .B2(_01914_),
    .C1(_06341_),
    .C2(_00161_),
    .Y(_06503_));
 OA21x2_ASAP7_75t_R _24408_ (.A1(_06266_),
    .A2(_05512_),
    .B(_06503_),
    .Y(_06504_));
 AO21x1_ASAP7_75t_R _24409_ (.A1(_06502_),
    .A2(_06504_),
    .B(net286),
    .Y(_06505_));
 OA21x2_ASAP7_75t_R _24410_ (.A1(_01520_),
    .A2(_06254_),
    .B(_06505_),
    .Y(_06506_));
 AND2x2_ASAP7_75t_R _24411_ (.A(_06312_),
    .B(_01729_),
    .Y(_06507_));
 AOI21x1_ASAP7_75t_R _24412_ (.A1(net415),
    .A2(_06506_),
    .B(_06507_),
    .Y(net241));
 INVx2_ASAP7_75t_R _24413_ (.A(net95),
    .Y(_06508_));
 INVx2_ASAP7_75t_R _24414_ (.A(_01815_),
    .Y(_06509_));
 INVx2_ASAP7_75t_R _24415_ (.A(_01736_),
    .Y(_06510_));
 CKINVDCx20_ASAP7_75t_R _24416_ (.A(_00239_),
    .Y(_06511_));
 BUFx2_ASAP7_75t_R input70 (.A(hart_id_i[17]),
    .Y(net70));
 OA21x2_ASAP7_75t_R _24418_ (.A1(_06509_),
    .A2(_06510_),
    .B(_06511_),
    .Y(_06513_));
 AOI21x1_ASAP7_75t_R _24419_ (.A1(_01714_),
    .A2(_01717_),
    .B(_06181_),
    .Y(_06514_));
 OAI21x1_ASAP7_75t_R _24420_ (.A1(_06324_),
    .A2(_06514_),
    .B(_00238_),
    .Y(_06515_));
 AO21x2_ASAP7_75t_R _24421_ (.A1(net287),
    .A2(_06513_),
    .B(_06515_),
    .Y(_06516_));
 AND2x4_ASAP7_75t_R _24422_ (.A(_00237_),
    .B(_06516_),
    .Y(_06517_));
 AO21x1_ASAP7_75t_R _24423_ (.A1(_00238_),
    .A2(net128),
    .B(_01736_),
    .Y(_06518_));
 OAI21x1_ASAP7_75t_R _24424_ (.A1(_06508_),
    .A2(_06517_),
    .B(_06518_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ));
 OR3x1_ASAP7_75t_R _24425_ (.A(_06508_),
    .B(_01736_),
    .C(_06517_),
    .Y(_06519_));
 AND2x4_ASAP7_75t_R _24426_ (.A(net128),
    .B(_06510_),
    .Y(_06520_));
 AOI21x1_ASAP7_75t_R _24427_ (.A1(_00238_),
    .A2(_06519_),
    .B(_06520_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ));
 AO21x1_ASAP7_75t_R _24428_ (.A1(_01735_),
    .A2(net287),
    .B(_00237_),
    .Y(_06521_));
 INVx1_ASAP7_75t_R _24429_ (.A(_06521_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ));
 OR3x1_ASAP7_75t_R _24430_ (.A(_06508_),
    .B(_01736_),
    .C(_06521_),
    .Y(_06522_));
 OA211x2_ASAP7_75t_R _24431_ (.A1(_00238_),
    .A2(net287),
    .B(_06522_),
    .C(_01848_),
    .Y(_06523_));
 OAI21x1_ASAP7_75t_R _24432_ (.A1(net128),
    .A2(_06254_),
    .B(_06510_),
    .Y(_06524_));
 OA211x2_ASAP7_75t_R _24433_ (.A1(_06508_),
    .A2(_06521_),
    .B(_06524_),
    .C(_01737_),
    .Y(_06525_));
 AO21x1_ASAP7_75t_R _24434_ (.A1(_06520_),
    .A2(_06523_),
    .B(_06525_),
    .Y(_06526_));
 INVx1_ASAP7_75t_R _24435_ (.A(_06526_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ));
 NOR2x1_ASAP7_75t_R _24436_ (.A(_06520_),
    .B(_06523_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ));
 BUFx2_ASAP7_75t_R input69 (.A(hart_id_i[16]),
    .Y(net69));
 CKINVDCx14_ASAP7_75t_R _24438_ (.A(net416),
    .Y(_06528_));
 BUFx2_ASAP7_75t_R input68 (.A(hart_id_i[15]),
    .Y(net68));
 BUFx2_ASAP7_75t_R input67 (.A(hart_id_i[14]),
    .Y(net67));
 BUFx2_ASAP7_75t_R input66 (.A(hart_id_i[13]),
    .Y(net66));
 INVx1_ASAP7_75t_R _24442_ (.A(net103),
    .Y(_06532_));
 BUFx2_ASAP7_75t_R input65 (.A(hart_id_i[12]),
    .Y(net65));
 NAND2x1_ASAP7_75t_R _24444_ (.A(_00240_),
    .B(net104),
    .Y(_06534_));
 OR3x1_ASAP7_75t_R _24445_ (.A(_00240_),
    .B(_01829_),
    .C(_01830_),
    .Y(_06535_));
 OA21x2_ASAP7_75t_R _24446_ (.A1(_06532_),
    .A2(_06534_),
    .B(_06535_),
    .Y(_06536_));
 CKINVDCx20_ASAP7_75t_R _24447_ (.A(net414),
    .Y(_06537_));
 INVx2_ASAP7_75t_R _24448_ (.A(net94),
    .Y(_06538_));
 AND2x2_ASAP7_75t_R _24449_ (.A(_00240_),
    .B(_06538_),
    .Y(_06539_));
 AO21x2_ASAP7_75t_R _24450_ (.A1(_06537_),
    .A2(_01814_),
    .B(_06539_),
    .Y(_06540_));
 AND3x2_ASAP7_75t_R _24451_ (.A(_06528_),
    .B(_06536_),
    .C(_06540_),
    .Y(_17534_));
 OR3x1_ASAP7_75t_R _24452_ (.A(_00242_),
    .B(_01605_),
    .C(_01606_),
    .Y(_06541_));
 INVx1_ASAP7_75t_R _24453_ (.A(_06541_),
    .Y(_18343_));
 OR5x2_ASAP7_75t_R _24454_ (.A(_00242_),
    .B(_01603_),
    .C(_01604_),
    .D(_01605_),
    .E(_01606_),
    .Y(_06542_));
 INVx1_ASAP7_75t_R _24455_ (.A(_06542_),
    .Y(_18344_));
 OR3x1_ASAP7_75t_R _24456_ (.A(_01601_),
    .B(_01602_),
    .C(_06542_),
    .Y(_06543_));
 INVx1_ASAP7_75t_R _24457_ (.A(_06543_),
    .Y(_18345_));
 OR3x1_ASAP7_75t_R _24458_ (.A(_01599_),
    .B(_01600_),
    .C(_06543_),
    .Y(_06544_));
 INVx1_ASAP7_75t_R _24459_ (.A(_06544_),
    .Y(_18346_));
 OR3x1_ASAP7_75t_R _24460_ (.A(_01597_),
    .B(_01598_),
    .C(_06544_),
    .Y(_06545_));
 INVx1_ASAP7_75t_R _24461_ (.A(_06545_),
    .Y(_18347_));
 OR3x1_ASAP7_75t_R _24462_ (.A(_01595_),
    .B(_01596_),
    .C(_06545_),
    .Y(_06546_));
 INVx1_ASAP7_75t_R _24463_ (.A(_06546_),
    .Y(_18348_));
 OR3x1_ASAP7_75t_R _24464_ (.A(_01593_),
    .B(_01594_),
    .C(_06546_),
    .Y(_06547_));
 INVx1_ASAP7_75t_R _24465_ (.A(_06547_),
    .Y(_18349_));
 OR3x1_ASAP7_75t_R _24466_ (.A(_01591_),
    .B(_01592_),
    .C(_06547_),
    .Y(_06548_));
 INVx1_ASAP7_75t_R _24467_ (.A(_06548_),
    .Y(_18350_));
 OR3x1_ASAP7_75t_R _24468_ (.A(_01589_),
    .B(_01590_),
    .C(_06548_),
    .Y(_06549_));
 INVx1_ASAP7_75t_R _24469_ (.A(_06549_),
    .Y(_18351_));
 OR3x1_ASAP7_75t_R _24470_ (.A(_01587_),
    .B(_01588_),
    .C(_06549_),
    .Y(_06550_));
 INVx1_ASAP7_75t_R _24471_ (.A(_06550_),
    .Y(_18352_));
 OR3x1_ASAP7_75t_R _24472_ (.A(_01585_),
    .B(_01586_),
    .C(_06550_),
    .Y(_06551_));
 INVx1_ASAP7_75t_R _24473_ (.A(_06551_),
    .Y(_18353_));
 OR3x1_ASAP7_75t_R _24474_ (.A(_01583_),
    .B(_01584_),
    .C(_06551_),
    .Y(_06552_));
 INVx1_ASAP7_75t_R _24475_ (.A(_06552_),
    .Y(_18354_));
 OR3x1_ASAP7_75t_R _24476_ (.A(_01581_),
    .B(_01582_),
    .C(_06552_),
    .Y(_06553_));
 INVx1_ASAP7_75t_R _24477_ (.A(_06553_),
    .Y(_18355_));
 AND2x2_ASAP7_75t_R _24478_ (.A(_06183_),
    .B(_01734_),
    .Y(_06554_));
 AO21x2_ASAP7_75t_R _24479_ (.A1(_06223_),
    .A2(_06554_),
    .B(_01747_),
    .Y(net150));
 AND3x2_ASAP7_75t_R _24480_ (.A(_01714_),
    .B(_01715_),
    .C(_05526_),
    .Y(_06555_));
 INVx1_ASAP7_75t_R _24481_ (.A(_06555_),
    .Y(_06556_));
 AND4x1_ASAP7_75t_R _24482_ (.A(_13227_),
    .B(_06178_),
    .C(_06186_),
    .D(_06556_),
    .Y(_06557_));
 OR3x2_ASAP7_75t_R _24483_ (.A(_06266_),
    .B(_05591_),
    .C(_05696_),
    .Y(_06558_));
 AOI211x1_ASAP7_75t_R _24484_ (.A1(_00282_),
    .A2(_13359_),
    .B(_14492_),
    .C(_13228_),
    .Y(_06559_));
 OR3x2_ASAP7_75t_R _24485_ (.A(_13384_),
    .B(_13336_),
    .C(_06559_),
    .Y(_06560_));
 NOR3x2_ASAP7_75t_R _24486_ (.B(_13380_),
    .C(_06560_),
    .Y(_06561_),
    .A(_13349_));
 OR3x1_ASAP7_75t_R _24487_ (.A(_13364_),
    .B(_13376_),
    .C(_06561_),
    .Y(_06562_));
 NAND3x2_ASAP7_75t_R _24488_ (.B(_13366_),
    .C(_06561_),
    .Y(_06563_),
    .A(_13329_));
 AO21x1_ASAP7_75t_R _24489_ (.A1(_06562_),
    .A2(_06563_),
    .B(_05478_),
    .Y(_06564_));
 NAND3x1_ASAP7_75t_R _24490_ (.A(_05478_),
    .B(_06562_),
    .C(_06563_),
    .Y(_06565_));
 AOI21x1_ASAP7_75t_R _24491_ (.A1(_06564_),
    .A2(_06565_),
    .B(_01310_),
    .Y(_06566_));
 AND5x1_ASAP7_75t_R _24492_ (.A(_01310_),
    .B(_05479_),
    .C(_05485_),
    .D(_05508_),
    .E(_05509_),
    .Y(_06567_));
 AOI211x1_ASAP7_75t_R _24493_ (.A1(_01310_),
    .A2(_05510_),
    .B(_06566_),
    .C(_06567_),
    .Y(_06568_));
 NAND3x1_ASAP7_75t_R _24494_ (.A(_13328_),
    .B(_13235_),
    .C(_13252_),
    .Y(_06569_));
 OR2x2_ASAP7_75t_R _24495_ (.A(_13382_),
    .B(_06569_),
    .Y(_06570_));
 OR2x2_ASAP7_75t_R _24496_ (.A(_05907_),
    .B(_06569_),
    .Y(_06571_));
 OA22x2_ASAP7_75t_R _24497_ (.A1(_06568_),
    .A2(_06570_),
    .B1(_06571_),
    .B2(_05777_),
    .Y(_06572_));
 NOR3x2_ASAP7_75t_R _24498_ (.B(_13356_),
    .C(_13363_),
    .Y(_06573_),
    .A(_13349_));
 OR3x4_ASAP7_75t_R _24499_ (.A(_13349_),
    .B(_13380_),
    .C(_06560_),
    .Y(_06574_));
 BUFx2_ASAP7_75t_R input64 (.A(hart_id_i[11]),
    .Y(net64));
 NAND2x2_ASAP7_75t_R _24501_ (.A(_13376_),
    .B(_06574_),
    .Y(_06576_));
 OA21x2_ASAP7_75t_R _24502_ (.A1(_13376_),
    .A2(_06574_),
    .B(_13364_),
    .Y(_06577_));
 AO21x1_ASAP7_75t_R _24503_ (.A1(_06573_),
    .A2(_06576_),
    .B(_06577_),
    .Y(_06578_));
 OA21x2_ASAP7_75t_R _24504_ (.A1(_13325_),
    .A2(_00282_),
    .B(_13329_),
    .Y(_06579_));
 AO21x1_ASAP7_75t_R _24505_ (.A1(_06578_),
    .A2(_06579_),
    .B(_13386_),
    .Y(_06580_));
 OR3x1_ASAP7_75t_R _24506_ (.A(_00281_),
    .B(_13381_),
    .C(_06569_),
    .Y(_06581_));
 AND4x1_ASAP7_75t_R _24507_ (.A(_13253_),
    .B(_05776_),
    .C(_06580_),
    .D(_06581_),
    .Y(_06582_));
 AOI21x1_ASAP7_75t_R _24508_ (.A1(_06578_),
    .A2(_06579_),
    .B(_13386_),
    .Y(_06583_));
 AND2x2_ASAP7_75t_R _24509_ (.A(_13253_),
    .B(_06583_),
    .Y(_06584_));
 AND4x2_ASAP7_75t_R _24510_ (.A(_01314_),
    .B(_01728_),
    .C(_13576_),
    .D(_05790_),
    .Y(_06585_));
 INVx1_ASAP7_75t_R _24511_ (.A(_05522_),
    .Y(_06586_));
 OA211x2_ASAP7_75t_R _24512_ (.A1(_01713_),
    .A2(_06586_),
    .B(_14615_),
    .C(_13227_),
    .Y(_06587_));
 AO21x1_ASAP7_75t_R _24513_ (.A1(_14585_),
    .A2(_06585_),
    .B(_06587_),
    .Y(_06588_));
 AO21x1_ASAP7_75t_R _24514_ (.A1(_14625_),
    .A2(_06588_),
    .B(_06162_),
    .Y(_06589_));
 AOI221x1_ASAP7_75t_R _24515_ (.A1(_05512_),
    .A2(_06582_),
    .B1(_06584_),
    .B2(_06568_),
    .C(_06589_),
    .Y(_06590_));
 AO21x1_ASAP7_75t_R _24516_ (.A1(_01713_),
    .A2(_05735_),
    .B(_06585_),
    .Y(_06591_));
 AO21x1_ASAP7_75t_R _24517_ (.A1(_14585_),
    .A2(_06591_),
    .B(_06587_),
    .Y(_06592_));
 NAND2x1_ASAP7_75t_R _24518_ (.A(_14625_),
    .B(_06592_),
    .Y(_06593_));
 AO21x2_ASAP7_75t_R _24519_ (.A1(_06572_),
    .A2(_06590_),
    .B(_06593_),
    .Y(_06594_));
 INVx1_ASAP7_75t_R _24520_ (.A(_06323_),
    .Y(_06595_));
 INVx1_ASAP7_75t_R _24521_ (.A(_14599_),
    .Y(_06596_));
 INVx1_ASAP7_75t_R _24522_ (.A(_02287_),
    .Y(_06597_));
 AND2x2_ASAP7_75t_R _24523_ (.A(_01744_),
    .B(_00245_),
    .Y(_06598_));
 AND4x1_ASAP7_75t_R _24524_ (.A(_02288_),
    .B(_06597_),
    .C(_06598_),
    .D(_05534_),
    .Y(_06599_));
 AND5x1_ASAP7_75t_R _24525_ (.A(_00245_),
    .B(_02287_),
    .C(_14155_),
    .D(_05720_),
    .E(_05534_),
    .Y(_06600_));
 AO21x1_ASAP7_75t_R _24526_ (.A1(_06596_),
    .A2(_06599_),
    .B(_06600_),
    .Y(_06601_));
 AND3x1_ASAP7_75t_R _24527_ (.A(_14585_),
    .B(_05535_),
    .C(_06601_),
    .Y(_06602_));
 INVx1_ASAP7_75t_R _24528_ (.A(_06602_),
    .Y(_06603_));
 AND4x1_ASAP7_75t_R _24529_ (.A(_05525_),
    .B(_05711_),
    .C(_06595_),
    .D(_06603_),
    .Y(_06604_));
 AO21x1_ASAP7_75t_R _24530_ (.A1(_05725_),
    .A2(_06604_),
    .B(_06266_),
    .Y(_06605_));
 AND2x2_ASAP7_75t_R _24531_ (.A(_06594_),
    .B(_06605_),
    .Y(_06606_));
 AND2x2_ASAP7_75t_R _24532_ (.A(_06558_),
    .B(_06606_),
    .Y(_06607_));
 INVx1_ASAP7_75t_R _24533_ (.A(_06607_),
    .Y(_06608_));
 INVx2_ASAP7_75t_R _24534_ (.A(_06191_),
    .Y(_06609_));
 NOR2x2_ASAP7_75t_R _24535_ (.A(_06609_),
    .B(_06223_),
    .Y(_06610_));
 NOR2x1_ASAP7_75t_R _24536_ (.A(_01317_),
    .B(_02034_),
    .Y(_06611_));
 OA21x2_ASAP7_75t_R _24537_ (.A1(net60),
    .A2(_06611_),
    .B(_01311_),
    .Y(_06612_));
 OA21x2_ASAP7_75t_R _24538_ (.A1(_06610_),
    .A2(_06612_),
    .B(_14583_),
    .Y(_06613_));
 BUFx2_ASAP7_75t_R input63 (.A(hart_id_i[10]),
    .Y(net63));
 BUFx2_ASAP7_75t_R input62 (.A(hart_id_i[0]),
    .Y(net62));
 AO21x1_ASAP7_75t_R _24541_ (.A1(_06536_),
    .A2(_06540_),
    .B(_00662_),
    .Y(_06616_));
 AND3x4_ASAP7_75t_R _24542_ (.A(net128),
    .B(_06510_),
    .C(_01737_),
    .Y(_06617_));
 BUFx2_ASAP7_75t_R input61 (.A(fetch_enable_i),
    .Y(net61));
 NAND2x1_ASAP7_75t_R _24544_ (.A(_06616_),
    .B(_06617_),
    .Y(_06619_));
 BUFx3_ASAP7_75t_R input60 (.A(debug_req_i),
    .Y(net60));
 OA211x2_ASAP7_75t_R _24546_ (.A1(_00239_),
    .A2(_06616_),
    .B(_06619_),
    .C(_00240_),
    .Y(_06621_));
 OR2x2_ASAP7_75t_R _24547_ (.A(_06511_),
    .B(_06617_),
    .Y(_06622_));
 NOR2x1_ASAP7_75t_R _24548_ (.A(_06616_),
    .B(_06622_),
    .Y(_06623_));
 OR5x2_ASAP7_75t_R _24549_ (.A(_05527_),
    .B(_06555_),
    .C(_06613_),
    .D(_06621_),
    .E(_06623_),
    .Y(_06624_));
 INVx1_ASAP7_75t_R _24550_ (.A(_06624_),
    .Y(_06625_));
 AND3x1_ASAP7_75t_R _24551_ (.A(_06226_),
    .B(_06607_),
    .C(_06625_),
    .Y(_06626_));
 AO21x1_ASAP7_75t_R _24552_ (.A1(_06557_),
    .A2(_06608_),
    .B(_06626_),
    .Y(\if_stage_i.instr_valid_id_d ));
 AND2x2_ASAP7_75t_R _24553_ (.A(_06580_),
    .B(_06581_),
    .Y(_06627_));
 AO22x1_ASAP7_75t_R _24554_ (.A1(_06568_),
    .A2(_06583_),
    .B1(_06627_),
    .B2(_05777_),
    .Y(_06628_));
 INVx1_ASAP7_75t_R _24555_ (.A(_06628_),
    .Y(_06629_));
 NAND2x1_ASAP7_75t_R _24556_ (.A(_06629_),
    .B(_06572_),
    .Y(_06630_));
 AND2x2_ASAP7_75t_R _24557_ (.A(_13253_),
    .B(_06630_),
    .Y(_06631_));
 AND4x1_ASAP7_75t_R _24558_ (.A(_01713_),
    .B(_05735_),
    .C(_05729_),
    .D(_06631_),
    .Y(\id_stage_i.branch_set_d ));
 INVx1_ASAP7_75t_R _24559_ (.A(_02566_),
    .Y(_18358_));
 AOI211x1_ASAP7_75t_R _24560_ (.A1(_01546_),
    .A2(net287),
    .B(_06310_),
    .C(_02566_),
    .Y(_06632_));
 AND2x2_ASAP7_75t_R _24561_ (.A(_18359_),
    .B(_06632_),
    .Y(_18360_));
 OR3x1_ASAP7_75t_R _24562_ (.A(_01544_),
    .B(_01545_),
    .C(_01547_),
    .Y(_06633_));
 OR4x1_ASAP7_75t_R _24563_ (.A(net287),
    .B(_06301_),
    .C(_06319_),
    .D(_06332_),
    .Y(_06634_));
 OAI21x1_ASAP7_75t_R _24564_ (.A1(_06254_),
    .A2(_06633_),
    .B(_06634_),
    .Y(_06635_));
 AND2x2_ASAP7_75t_R _24565_ (.A(_06632_),
    .B(_06635_),
    .Y(_18362_));
 OR2x2_ASAP7_75t_R _24566_ (.A(_01542_),
    .B(_01543_),
    .Y(_06636_));
 OR3x1_ASAP7_75t_R _24567_ (.A(net287),
    .B(_06346_),
    .C(_06354_),
    .Y(_06637_));
 OAI21x1_ASAP7_75t_R _24568_ (.A1(_06254_),
    .A2(_06636_),
    .B(_06637_),
    .Y(_06638_));
 AND3x1_ASAP7_75t_R _24569_ (.A(_06632_),
    .B(_06635_),
    .C(_06638_),
    .Y(_18364_));
 NOR2x1_ASAP7_75t_R _24570_ (.A(_01540_),
    .B(_01541_),
    .Y(_06639_));
 NAND2x1_ASAP7_75t_R _24571_ (.A(_06367_),
    .B(_06373_),
    .Y(_06640_));
 AO32x1_ASAP7_75t_R _24572_ (.A1(net1),
    .A2(net2),
    .A3(_06339_),
    .B1(_06361_),
    .B2(_06640_),
    .Y(_06641_));
 AND2x2_ASAP7_75t_R _24573_ (.A(_06254_),
    .B(_06641_),
    .Y(_06642_));
 AO21x1_ASAP7_75t_R _24574_ (.A1(net287),
    .A2(_06639_),
    .B(_06642_),
    .Y(_06643_));
 AND2x2_ASAP7_75t_R _24575_ (.A(_18364_),
    .B(_06643_),
    .Y(_18367_));
 OR3x1_ASAP7_75t_R _24576_ (.A(_01538_),
    .B(_01539_),
    .C(_06254_),
    .Y(_06644_));
 OR3x1_ASAP7_75t_R _24577_ (.A(net287),
    .B(_06380_),
    .C(_06388_),
    .Y(_06645_));
 NAND2x1_ASAP7_75t_R _24578_ (.A(_06644_),
    .B(_06645_),
    .Y(_06646_));
 AND5x2_ASAP7_75t_R _24579_ (.A(_06632_),
    .B(_06635_),
    .C(_06638_),
    .D(_06643_),
    .E(_06646_),
    .Y(_18369_));
 NOR2x1_ASAP7_75t_R _24580_ (.A(_01536_),
    .B(_01537_),
    .Y(_06647_));
 AND3x1_ASAP7_75t_R _24581_ (.A(_06254_),
    .B(_06394_),
    .C(_06399_),
    .Y(_06648_));
 AO21x1_ASAP7_75t_R _24582_ (.A1(net286),
    .A2(_06647_),
    .B(_06648_),
    .Y(_06649_));
 AND2x2_ASAP7_75t_R _24583_ (.A(_18369_),
    .B(_06649_),
    .Y(_18371_));
 AND4x1_ASAP7_75t_R _24584_ (.A(_18370_),
    .B(_06417_),
    .C(_18369_),
    .D(_06649_),
    .Y(_18373_));
 AND3x1_ASAP7_75t_R _24585_ (.A(_18372_),
    .B(_06430_),
    .C(_18373_),
    .Y(_18375_));
 AND3x2_ASAP7_75t_R _24586_ (.A(_18374_),
    .B(_06444_),
    .C(_18375_),
    .Y(_18377_));
 AND2x2_ASAP7_75t_R _24587_ (.A(_18376_),
    .B(_06456_),
    .Y(_06650_));
 AND2x2_ASAP7_75t_R _24588_ (.A(_18377_),
    .B(_06650_),
    .Y(_18379_));
 AND4x1_ASAP7_75t_R _24589_ (.A(_18378_),
    .B(_06469_),
    .C(_18377_),
    .D(_06650_),
    .Y(_18381_));
 AND3x1_ASAP7_75t_R _24590_ (.A(_18380_),
    .B(_06482_),
    .C(_18381_),
    .Y(_18383_));
 AND3x1_ASAP7_75t_R _24591_ (.A(_18382_),
    .B(_06495_),
    .C(_18383_),
    .Y(_18385_));
 AND3x1_ASAP7_75t_R _24592_ (.A(_01311_),
    .B(_06223_),
    .C(_06184_),
    .Y(_06651_));
 AND5x1_ASAP7_75t_R _24593_ (.A(_00238_),
    .B(_01608_),
    .C(_01609_),
    .D(_01736_),
    .E(_06555_),
    .Y(_06652_));
 OA211x2_ASAP7_75t_R _24594_ (.A1(_01717_),
    .A2(_06651_),
    .B(_06652_),
    .C(_00277_),
    .Y(_06653_));
 NAND2x1_ASAP7_75t_R _24595_ (.A(_06517_),
    .B(_06653_),
    .Y(core_busy_d));
 AND2x2_ASAP7_75t_R _24596_ (.A(clknet_leaf_24_clk_i),
    .B(\core_clock_gate_i.en_latch ),
    .Y(\core_clock_gate_i.clk_o ));
 INVx1_ASAP7_75t_R _24597_ (.A(net149),
    .Y(_06654_));
 NAND2x1_ASAP7_75t_R _24598_ (.A(_06654_),
    .B(net150),
    .Y(_00008_));
 INVx1_ASAP7_75t_R _24599_ (.A(_06517_),
    .Y(net249));
 NOR2x1_ASAP7_75t_R _24600_ (.A(net95),
    .B(_06517_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ));
 NOR3x2_ASAP7_75t_R _24601_ (.B(_05591_),
    .C(_05696_),
    .Y(_06655_),
    .A(_06266_));
 NAND2x1_ASAP7_75t_R _24602_ (.A(_06594_),
    .B(_06605_),
    .Y(_06656_));
 BUFx3_ASAP7_75t_R input59 (.A(data_rvalid_i),
    .Y(net59));
 BUFx3_ASAP7_75t_R input58 (.A(data_rdata_i[9]),
    .Y(net58));
 OA211x2_ASAP7_75t_R _24605_ (.A1(_01845_),
    .A2(_01846_),
    .B(_06537_),
    .C(_01814_),
    .Y(_06659_));
 AND3x1_ASAP7_75t_R _24606_ (.A(_00240_),
    .B(net107),
    .C(net96),
    .Y(_06660_));
 INVx1_ASAP7_75t_R _24607_ (.A(_06660_),
    .Y(_06661_));
 BUFx3_ASAP7_75t_R input57 (.A(data_rdata_i[8]),
    .Y(net57));
 BUFx3_ASAP7_75t_R input56 (.A(data_rdata_i[7]),
    .Y(net56));
 OA211x2_ASAP7_75t_R _24610_ (.A1(_06539_),
    .A2(_06659_),
    .B(_06661_),
    .C(_00662_),
    .Y(_06664_));
 OR2x2_ASAP7_75t_R _24611_ (.A(_06624_),
    .B(_06664_),
    .Y(_06665_));
 OR3x4_ASAP7_75t_R _24612_ (.A(_06655_),
    .B(_06656_),
    .C(_06665_),
    .Y(_06666_));
 BUFx3_ASAP7_75t_R input55 (.A(data_rdata_i[6]),
    .Y(net55));
 BUFx3_ASAP7_75t_R input54 (.A(data_rdata_i[5]),
    .Y(net54));
 OA21x2_ASAP7_75t_R _24615_ (.A1(_06617_),
    .A2(_06666_),
    .B(_06511_),
    .Y(_06669_));
 NAND2x2_ASAP7_75t_R _24616_ (.A(_01737_),
    .B(_06520_),
    .Y(_06670_));
 BUFx2_ASAP7_75t_R input53 (.A(data_rdata_i[4]),
    .Y(net53));
 BUFx3_ASAP7_75t_R input52 (.A(data_rdata_i[3]),
    .Y(net52));
 NAND2x1_ASAP7_75t_R _24619_ (.A(_06537_),
    .B(_06666_),
    .Y(_06673_));
 OR2x6_ASAP7_75t_R _24620_ (.A(_01815_),
    .B(_06666_),
    .Y(_06674_));
 BUFx3_ASAP7_75t_R input51 (.A(data_rdata_i[31]),
    .Y(net51));
 BUFx2_ASAP7_75t_R input50 (.A(data_rdata_i[30]),
    .Y(net50));
 OAI21x1_ASAP7_75t_R _24623_ (.A1(_06670_),
    .A2(_06673_),
    .B(_06674_),
    .Y(_06677_));
 BUFx2_ASAP7_75t_R input49 (.A(data_rdata_i[2]),
    .Y(net49));
 OA21x2_ASAP7_75t_R _24625_ (.A1(_06669_),
    .A2(_06677_),
    .B(net287),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ));
 BUFx3_ASAP7_75t_R input48 (.A(data_rdata_i[29]),
    .Y(net48));
 NOR2x2_ASAP7_75t_R _24627_ (.A(_00239_),
    .B(_06666_),
    .Y(_06680_));
 AO21x1_ASAP7_75t_R _24628_ (.A1(_06617_),
    .A2(_06666_),
    .B(_06680_),
    .Y(_06681_));
 BUFx2_ASAP7_75t_R input47 (.A(data_rdata_i[28]),
    .Y(net47));
 OA21x2_ASAP7_75t_R _24630_ (.A1(_06622_),
    .A2(_06666_),
    .B(net287),
    .Y(_06683_));
 OA21x2_ASAP7_75t_R _24631_ (.A1(_06537_),
    .A2(_06681_),
    .B(_06683_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ));
 AO21x1_ASAP7_75t_R _24632_ (.A1(_06511_),
    .A2(_06617_),
    .B(_06509_),
    .Y(_06684_));
 AND3x1_ASAP7_75t_R _24633_ (.A(net287),
    .B(_06666_),
    .C(_06684_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ));
 INVx1_ASAP7_75t_R _24634_ (.A(_00660_),
    .Y(\cs_registers_i.mhpmcounter[2][0] ));
 INVx1_ASAP7_75t_R _24635_ (.A(_00659_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[0] ));
 INVx1_ASAP7_75t_R _24636_ (.A(_17536_),
    .Y(\cs_registers_i.pc_if_i[2] ));
 INVx1_ASAP7_75t_R _24637_ (.A(_17601_),
    .Y(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ));
 NAND2x1_ASAP7_75t_R _24638_ (.A(_05835_),
    .B(_05855_),
    .Y(_16776_));
 BUFx3_ASAP7_75t_R input46 (.A(data_rdata_i[27]),
    .Y(net46));
 NAND2x1_ASAP7_75t_R _24640_ (.A(_05832_),
    .B(_05858_),
    .Y(_16784_));
 BUFx2_ASAP7_75t_R input45 (.A(data_rdata_i[26]),
    .Y(net45));
 NAND2x1_ASAP7_75t_R _24642_ (.A(_05893_),
    .B(_05928_),
    .Y(_16798_));
 BUFx2_ASAP7_75t_R input44 (.A(data_rdata_i[25]),
    .Y(net44));
 NAND2x1_ASAP7_75t_R _24644_ (.A(_05835_),
    .B(_05936_),
    .Y(_16816_));
 NAND2x1_ASAP7_75t_R _24645_ (.A(_05832_),
    .B(_05863_),
    .Y(_16826_));
 NAND2x1_ASAP7_75t_R _24646_ (.A(_05904_),
    .B(_05928_),
    .Y(_16843_));
 NAND2x1_ASAP7_75t_R _24647_ (.A(_05843_),
    .B(_05936_),
    .Y(_16864_));
 BUFx3_ASAP7_75t_R input43 (.A(data_rdata_i[24]),
    .Y(net43));
 NAND2x1_ASAP7_75t_R _24649_ (.A(_05840_),
    .B(_05863_),
    .Y(_16873_));
 BUFx4f_ASAP7_75t_R input42 (.A(data_rdata_i[23]),
    .Y(net42));
 NAND2x1_ASAP7_75t_R _24651_ (.A(_05796_),
    .B(_05924_),
    .Y(_16889_));
 NAND2x2_ASAP7_75t_R _24652_ (.A(_05898_),
    .B(_05916_),
    .Y(_17494_));
 NAND2x1_ASAP7_75t_R _24653_ (.A(_05815_),
    .B(_05928_),
    .Y(_16547_));
 NAND2x1_ASAP7_75t_R _24654_ (.A(_05819_),
    .B(_05928_),
    .Y(_16550_));
 NAND2x1_ASAP7_75t_R _24655_ (.A(_05828_),
    .B(_05928_),
    .Y(_16557_));
 NAND2x1_ASAP7_75t_R _24656_ (.A(_05835_),
    .B(_05928_),
    .Y(_16571_));
 NAND2x1_ASAP7_75t_R _24657_ (.A(_05843_),
    .B(_05928_),
    .Y(_16592_));
 NAND2x1_ASAP7_75t_R _24658_ (.A(_05851_),
    .B(_05928_),
    .Y(_16611_));
 NAND2x1_ASAP7_75t_R _24659_ (.A(_05815_),
    .B(_05840_),
    .Y(_16625_));
 NAND2x1_ASAP7_75t_R _24660_ (.A(_05858_),
    .B(_05928_),
    .Y(_16637_));
 NAND2x1_ASAP7_75t_R _24661_ (.A(_05819_),
    .B(_05840_),
    .Y(_16655_));
 NAND2x1_ASAP7_75t_R _24662_ (.A(_05863_),
    .B(_05928_),
    .Y(_16664_));
 NAND2x1_ASAP7_75t_R _24663_ (.A(_05828_),
    .B(_05840_),
    .Y(_16679_));
 NAND2x1_ASAP7_75t_R _24664_ (.A(_05871_),
    .B(_05928_),
    .Y(_16692_));
 NAND2x1_ASAP7_75t_R _24665_ (.A(_05815_),
    .B(_05936_),
    .Y(_16709_));
 NAND2x1_ASAP7_75t_R _24666_ (.A(_05835_),
    .B(_05840_),
    .Y(_16712_));
 NAND2x1_ASAP7_75t_R _24667_ (.A(_05878_),
    .B(_05928_),
    .Y(_16725_));
 NAND2x1_ASAP7_75t_R _24668_ (.A(_05819_),
    .B(_05936_),
    .Y(_16741_));
 NAND2x1_ASAP7_75t_R _24669_ (.A(_05840_),
    .B(_05843_),
    .Y(_16744_));
 NAND2x1_ASAP7_75t_R _24670_ (.A(_05883_),
    .B(_05928_),
    .Y(_16759_));
 NAND2x1_ASAP7_75t_R _24671_ (.A(_05819_),
    .B(_05875_),
    .Y(_16813_));
 NAND2x1_ASAP7_75t_R _24672_ (.A(_05843_),
    .B(_05855_),
    .Y(_16817_));
 NAND2x1_ASAP7_75t_R _24673_ (.A(_05840_),
    .B(_05858_),
    .Y(_16827_));
 NAND2x1_ASAP7_75t_R _24674_ (.A(_05796_),
    .B(_05920_),
    .Y(_16844_));
 NAND2x1_ASAP7_75t_R _24675_ (.A(_05851_),
    .B(_05855_),
    .Y(_16865_));
 NAND2x1_ASAP7_75t_R _24676_ (.A(_05832_),
    .B(_05871_),
    .Y(_16874_));
 OA22x2_ASAP7_75t_R _24677_ (.A1(_01314_),
    .A2(_01677_),
    .B1(_05519_),
    .B2(_00816_),
    .Y(_16904_));
 NAND2x1_ASAP7_75t_R _24678_ (.A(_05843_),
    .B(_05867_),
    .Y(_16915_));
 NAND2x1_ASAP7_75t_R _24679_ (.A(_05846_),
    .B(_05863_),
    .Y(_16924_));
 NAND2x1_ASAP7_75t_R _24680_ (.A(_05807_),
    .B(_05920_),
    .Y(_16941_));
 OR2x2_ASAP7_75t_R _24681_ (.A(_05815_),
    .B(_05911_),
    .Y(_16959_));
 NAND2x1_ASAP7_75t_R _24682_ (.A(_05858_),
    .B(_05936_),
    .Y(_16970_));
 NAND2x1_ASAP7_75t_R _24683_ (.A(_05840_),
    .B(_05878_),
    .Y(_16981_));
 OR2x2_ASAP7_75t_R _24684_ (.A(_05819_),
    .B(_05911_),
    .Y(_17009_));
 NAND2x1_ASAP7_75t_R _24685_ (.A(_05863_),
    .B(_05936_),
    .Y(_17020_));
 NAND2x1_ASAP7_75t_R _24686_ (.A(_05840_),
    .B(_05883_),
    .Y(_17030_));
 NAND2x1_ASAP7_75t_R _24687_ (.A(_05825_),
    .B(_05920_),
    .Y(_17035_));
 OR2x2_ASAP7_75t_R _24688_ (.A(_05828_),
    .B(_05911_),
    .Y(_17060_));
 NAND2x1_ASAP7_75t_R _24689_ (.A(_05871_),
    .B(_05936_),
    .Y(_17071_));
 NAND2x1_ASAP7_75t_R _24690_ (.A(_05840_),
    .B(_05893_),
    .Y(_17081_));
 NAND2x1_ASAP7_75t_R _24691_ (.A(_05825_),
    .B(_05924_),
    .Y(_17086_));
 OR2x2_ASAP7_75t_R _24692_ (.A(_05835_),
    .B(_05911_),
    .Y(_17104_));
 NAND2x1_ASAP7_75t_R _24693_ (.A(_05878_),
    .B(_05936_),
    .Y(_17115_));
 NAND2x1_ASAP7_75t_R _24694_ (.A(_05840_),
    .B(_05904_),
    .Y(_17125_));
 OR2x2_ASAP7_75t_R _24695_ (.A(_05843_),
    .B(_05911_),
    .Y(_17148_));
 NAND2x1_ASAP7_75t_R _24696_ (.A(_05863_),
    .B(_05901_),
    .Y(_17153_));
 NAND2x1_ASAP7_75t_R _24697_ (.A(_05883_),
    .B(_05936_),
    .Y(_17160_));
 NAND2x1_ASAP7_75t_R _24698_ (.A(_05840_),
    .B(_05920_),
    .Y(_17170_));
 OR2x2_ASAP7_75t_R _24699_ (.A(_05851_),
    .B(_05911_),
    .Y(_17196_));
 NAND2x1_ASAP7_75t_R _24700_ (.A(_05871_),
    .B(_05901_),
    .Y(_17201_));
 NAND2x1_ASAP7_75t_R _24701_ (.A(_05893_),
    .B(_05936_),
    .Y(_17208_));
 NAND2x1_ASAP7_75t_R _24702_ (.A(_05840_),
    .B(_05924_),
    .Y(_17217_));
 OR2x2_ASAP7_75t_R _24703_ (.A(_05858_),
    .B(_05911_),
    .Y(_17239_));
 NAND2x1_ASAP7_75t_R _24704_ (.A(_05878_),
    .B(_05901_),
    .Y(_17244_));
 NAND2x1_ASAP7_75t_R _24705_ (.A(_05904_),
    .B(_05936_),
    .Y(_17251_));
 OR2x2_ASAP7_75t_R _24706_ (.A(_05863_),
    .B(_05911_),
    .Y(_17275_));
 NAND2x1_ASAP7_75t_R _24707_ (.A(_05883_),
    .B(_05901_),
    .Y(_17280_));
 NAND2x1_ASAP7_75t_R _24708_ (.A(_05920_),
    .B(_05936_),
    .Y(_17287_));
 OR2x2_ASAP7_75t_R _24709_ (.A(_05871_),
    .B(_05911_),
    .Y(_17317_));
 NAND2x1_ASAP7_75t_R _24710_ (.A(_05893_),
    .B(_05901_),
    .Y(_17322_));
 NAND2x1_ASAP7_75t_R _24711_ (.A(_05924_),
    .B(_05936_),
    .Y(_17329_));
 OR2x2_ASAP7_75t_R _24712_ (.A(_05878_),
    .B(_05911_),
    .Y(_17351_));
 NAND2x1_ASAP7_75t_R _24713_ (.A(_05901_),
    .B(_05904_),
    .Y(_17356_));
 OR2x2_ASAP7_75t_R _24714_ (.A(_05883_),
    .B(_05911_),
    .Y(_17383_));
 NAND2x1_ASAP7_75t_R _24715_ (.A(_05901_),
    .B(_05920_),
    .Y(_17388_));
 OR2x2_ASAP7_75t_R _24716_ (.A(_05893_),
    .B(_05911_),
    .Y(_17413_));
 NAND2x1_ASAP7_75t_R _24717_ (.A(_05901_),
    .B(_05924_),
    .Y(_17418_));
 OR2x2_ASAP7_75t_R _24718_ (.A(_05904_),
    .B(_05911_),
    .Y(_17441_));
 OR2x2_ASAP7_75t_R _24719_ (.A(_05911_),
    .B(_05920_),
    .Y(_17463_));
 OR2x2_ASAP7_75t_R _24720_ (.A(_05911_),
    .B(_05924_),
    .Y(_17493_));
 NAND2x1_ASAP7_75t_R _24721_ (.A(_05796_),
    .B(_05819_),
    .Y(_16548_));
 NAND2x1_ASAP7_75t_R _24722_ (.A(_05796_),
    .B(_05828_),
    .Y(_16551_));
 NAND2x1_ASAP7_75t_R _24723_ (.A(_05796_),
    .B(_05835_),
    .Y(_16558_));
 NAND2x1_ASAP7_75t_R _24724_ (.A(_05796_),
    .B(_05843_),
    .Y(_16572_));
 NAND2x1_ASAP7_75t_R _24725_ (.A(_05796_),
    .B(_05851_),
    .Y(_16593_));
 NAND2x1_ASAP7_75t_R _24726_ (.A(_05796_),
    .B(_05858_),
    .Y(_16612_));
 NAND2x1_ASAP7_75t_R _24727_ (.A(_05819_),
    .B(_05832_),
    .Y(_16626_));
 NAND2x1_ASAP7_75t_R _24728_ (.A(_05796_),
    .B(_05863_),
    .Y(_16638_));
 NAND2x1_ASAP7_75t_R _24729_ (.A(_05828_),
    .B(_05832_),
    .Y(_16656_));
 NAND2x1_ASAP7_75t_R _24730_ (.A(_05796_),
    .B(_05871_),
    .Y(_16665_));
 NAND2x1_ASAP7_75t_R _24731_ (.A(_05832_),
    .B(_05835_),
    .Y(_16680_));
 NAND2x1_ASAP7_75t_R _24732_ (.A(_05796_),
    .B(_05878_),
    .Y(_16693_));
 NAND2x1_ASAP7_75t_R _24733_ (.A(_05819_),
    .B(_05855_),
    .Y(_16710_));
 NAND2x1_ASAP7_75t_R _24734_ (.A(_05832_),
    .B(_05843_),
    .Y(_16713_));
 NAND2x1_ASAP7_75t_R _24735_ (.A(_05796_),
    .B(_05883_),
    .Y(_16726_));
 NAND2x1_ASAP7_75t_R _24736_ (.A(_05828_),
    .B(_05855_),
    .Y(_16742_));
 NAND2x1_ASAP7_75t_R _24737_ (.A(_05832_),
    .B(_05851_),
    .Y(_16745_));
 NAND2x1_ASAP7_75t_R _24738_ (.A(_05796_),
    .B(_05893_),
    .Y(_16760_));
 NAND2x1_ASAP7_75t_R _24739_ (.A(_05828_),
    .B(_05936_),
    .Y(_16778_));
 NAND2x1_ASAP7_75t_R _24740_ (.A(_05840_),
    .B(_05851_),
    .Y(_16786_));
 NAND2x1_ASAP7_75t_R _24741_ (.A(_05796_),
    .B(_05904_),
    .Y(_16800_));
 NAND2x1_ASAP7_75t_R _24742_ (.A(_05815_),
    .B(_05901_),
    .Y(_16814_));
 NAND2x1_ASAP7_75t_R _24743_ (.A(_05920_),
    .B(_05928_),
    .Y(_16891_));
 OR2x2_ASAP7_75t_R _24744_ (.A(_05803_),
    .B(_05911_),
    .Y(_16905_));
 NAND2x1_ASAP7_75t_R _24745_ (.A(_05851_),
    .B(_05936_),
    .Y(_16916_));
 NAND2x1_ASAP7_75t_R _24746_ (.A(_05840_),
    .B(_05871_),
    .Y(_16925_));
 NAND2x1_ASAP7_75t_R _24747_ (.A(_05924_),
    .B(_05928_),
    .Y(_16942_));
 OA211x2_ASAP7_75t_R _24748_ (.A1(_05946_),
    .A2(_05947_),
    .B(_05949_),
    .C(_00025_),
    .Y(_06690_));
 OA21x2_ASAP7_75t_R _24749_ (.A1(_00024_),
    .A2(_06690_),
    .B(_02342_),
    .Y(_16957_));
 BUFx3_ASAP7_75t_R input41 (.A(data_rdata_i[22]),
    .Y(net41));
 NAND2x1_ASAP7_75t_R _24751_ (.A(_05819_),
    .B(_05898_),
    .Y(_16960_));
 NAND2x1_ASAP7_75t_R _24752_ (.A(_05855_),
    .B(_05863_),
    .Y(_16971_));
 NAND2x1_ASAP7_75t_R _24753_ (.A(_05832_),
    .B(_05883_),
    .Y(_16982_));
 NAND2x1_ASAP7_75t_R _24754_ (.A(_05828_),
    .B(_05898_),
    .Y(_17010_));
 NAND2x1_ASAP7_75t_R _24755_ (.A(_05855_),
    .B(_05871_),
    .Y(_17021_));
 NAND2x1_ASAP7_75t_R _24756_ (.A(_05832_),
    .B(_05893_),
    .Y(_17031_));
 NAND2x1_ASAP7_75t_R _24757_ (.A(_05812_),
    .B(_05924_),
    .Y(_17036_));
 NAND2x1_ASAP7_75t_R _24758_ (.A(_05835_),
    .B(_05898_),
    .Y(_17061_));
 NAND2x1_ASAP7_75t_R _24759_ (.A(_05855_),
    .B(_05878_),
    .Y(_17072_));
 NAND2x1_ASAP7_75t_R _24760_ (.A(_05832_),
    .B(_05904_),
    .Y(_17082_));
 NAND2x1_ASAP7_75t_R _24761_ (.A(_05843_),
    .B(_05898_),
    .Y(_17105_));
 NAND2x1_ASAP7_75t_R _24762_ (.A(_05855_),
    .B(_05883_),
    .Y(_17116_));
 NAND2x1_ASAP7_75t_R _24763_ (.A(_05832_),
    .B(_05920_),
    .Y(_17126_));
 NAND2x1_ASAP7_75t_R _24764_ (.A(_05851_),
    .B(_05898_),
    .Y(_17149_));
 NAND2x1_ASAP7_75t_R _24765_ (.A(_05871_),
    .B(_05875_),
    .Y(_17154_));
 NAND2x1_ASAP7_75t_R _24766_ (.A(_05855_),
    .B(_05893_),
    .Y(_17161_));
 NAND2x1_ASAP7_75t_R _24767_ (.A(_05832_),
    .B(_05924_),
    .Y(_17171_));
 NAND2x1_ASAP7_75t_R _24768_ (.A(_05858_),
    .B(_05898_),
    .Y(_17197_));
 NAND2x1_ASAP7_75t_R _24769_ (.A(_05875_),
    .B(_05878_),
    .Y(_17202_));
 NAND2x1_ASAP7_75t_R _24770_ (.A(_05855_),
    .B(_05904_),
    .Y(_17209_));
 NAND2x1_ASAP7_75t_R _24771_ (.A(_05863_),
    .B(_05898_),
    .Y(_17240_));
 NAND2x1_ASAP7_75t_R _24772_ (.A(_05875_),
    .B(_05883_),
    .Y(_17245_));
 NAND2x1_ASAP7_75t_R _24773_ (.A(_05855_),
    .B(_05920_),
    .Y(_17252_));
 NAND2x1_ASAP7_75t_R _24774_ (.A(_05871_),
    .B(_05898_),
    .Y(_17276_));
 NAND2x1_ASAP7_75t_R _24775_ (.A(_05875_),
    .B(_05893_),
    .Y(_17281_));
 NAND2x1_ASAP7_75t_R _24776_ (.A(_05855_),
    .B(_05924_),
    .Y(_17288_));
 NAND2x1_ASAP7_75t_R _24777_ (.A(_05878_),
    .B(_05898_),
    .Y(_17318_));
 NAND2x1_ASAP7_75t_R _24778_ (.A(_05875_),
    .B(_05904_),
    .Y(_17323_));
 NAND2x1_ASAP7_75t_R _24779_ (.A(_05883_),
    .B(_05898_),
    .Y(_17352_));
 NAND2x1_ASAP7_75t_R _24780_ (.A(_05875_),
    .B(_05920_),
    .Y(_17357_));
 NAND2x1_ASAP7_75t_R _24781_ (.A(_05893_),
    .B(_05898_),
    .Y(_17384_));
 NAND2x1_ASAP7_75t_R _24782_ (.A(_05875_),
    .B(_05924_),
    .Y(_17389_));
 NAND2x1_ASAP7_75t_R _24783_ (.A(_05898_),
    .B(_05904_),
    .Y(_17414_));
 NAND2x1_ASAP7_75t_R _24784_ (.A(_05898_),
    .B(_05920_),
    .Y(_17442_));
 NAND2x1_ASAP7_75t_R _24785_ (.A(_05898_),
    .B(_05924_),
    .Y(_17464_));
 OR3x2_ASAP7_75t_R _24786_ (.A(_05788_),
    .B(_05910_),
    .C(_05916_),
    .Y(_17518_));
 BUFx3_ASAP7_75t_R input40 (.A(data_rdata_i[21]),
    .Y(net40));
 BUFx3_ASAP7_75t_R input39 (.A(data_rdata_i[20]),
    .Y(net39));
 BUFx3_ASAP7_75t_R input38 (.A(data_rdata_i[1]),
    .Y(net38));
 OR3x1_ASAP7_75t_R _24790_ (.A(_00663_),
    .B(net294),
    .C(_13574_),
    .Y(_06695_));
 OAI21x1_ASAP7_75t_R _24791_ (.A1(_13576_),
    .A2(_14688_),
    .B(_06695_),
    .Y(_17540_));
 BUFx3_ASAP7_75t_R input37 (.A(data_rdata_i[19]),
    .Y(net37));
 XNOR2x1_ASAP7_75t_R _24793_ (.B(_14083_),
    .Y(_06697_),
    .A(_13387_));
 BUFx3_ASAP7_75t_R input36 (.A(data_rdata_i[18]),
    .Y(net36));
 INVx1_ASAP7_75t_R _24795_ (.A(_00668_),
    .Y(_06699_));
 INVx1_ASAP7_75t_R _24796_ (.A(_01448_),
    .Y(_06700_));
 OA222x2_ASAP7_75t_R _24797_ (.A1(_00285_),
    .A2(_06699_),
    .B1(_06700_),
    .B2(_13574_),
    .C1(_13763_),
    .C2(_14080_),
    .Y(_06701_));
 OA211x2_ASAP7_75t_R _24798_ (.A1(_00284_),
    .A2(_14820_),
    .B(_06701_),
    .C(_13576_),
    .Y(_06702_));
 AOI21x1_ASAP7_75t_R _24799_ (.A1(net294),
    .A2(_06697_),
    .B(_06702_),
    .Y(_17544_));
 XNOR2x1_ASAP7_75t_R _24800_ (.B(_18135_),
    .Y(_06703_),
    .A(_13387_));
 INVx1_ASAP7_75t_R _24801_ (.A(_14936_),
    .Y(_06704_));
 INVx6_ASAP7_75t_R _24802_ (.A(_00284_),
    .Y(_06705_));
 BUFx3_ASAP7_75t_R input35 (.A(data_rdata_i[17]),
    .Y(net35));
 BUFx4f_ASAP7_75t_R input34 (.A(data_rdata_i[16]),
    .Y(net34));
 AO221x1_ASAP7_75t_R _24805_ (.A1(_13530_),
    .A2(_00672_),
    .B1(_01446_),
    .B2(_13533_),
    .C(net295),
    .Y(_06708_));
 AO221x1_ASAP7_75t_R _24806_ (.A1(_13528_),
    .A2(_05605_),
    .B1(_06704_),
    .B2(_06705_),
    .C(_06708_),
    .Y(_06709_));
 OA21x2_ASAP7_75t_R _24807_ (.A1(_13576_),
    .A2(_06703_),
    .B(_06709_),
    .Y(_17548_));
 NAND2x2_ASAP7_75t_R _24808_ (.A(_14961_),
    .B(_14989_),
    .Y(_06710_));
 BUFx3_ASAP7_75t_R input33 (.A(data_rdata_i[15]),
    .Y(net33));
 AO221x1_ASAP7_75t_R _24810_ (.A1(_13530_),
    .A2(_00674_),
    .B1(_01445_),
    .B2(_13533_),
    .C(net295),
    .Y(_06712_));
 AO221x1_ASAP7_75t_R _24811_ (.A1(_13528_),
    .A2(_05653_),
    .B1(_06710_),
    .B2(_06705_),
    .C(_06712_),
    .Y(_06713_));
 OAI21x1_ASAP7_75t_R _24812_ (.A1(_13387_),
    .A2(_14256_),
    .B(net294),
    .Y(_06714_));
 AO22x2_ASAP7_75t_R _24813_ (.A1(_13781_),
    .A2(_14256_),
    .B1(_06713_),
    .B2(_06714_),
    .Y(_16510_));
 BUFx2_ASAP7_75t_R input32 (.A(data_rdata_i[14]),
    .Y(net32));
 NAND2x1_ASAP7_75t_R _24815_ (.A(_13781_),
    .B(_18147_),
    .Y(_06716_));
 AO22x1_ASAP7_75t_R _24816_ (.A1(_13530_),
    .A2(_00677_),
    .B1(_01444_),
    .B2(_13533_),
    .Y(_06717_));
 OAI22x1_ASAP7_75t_R _24817_ (.A1(_13763_),
    .A2(_14316_),
    .B1(_15042_),
    .B2(_00284_),
    .Y(_06718_));
 OR3x1_ASAP7_75t_R _24818_ (.A(net295),
    .B(_06717_),
    .C(_06718_),
    .Y(_06719_));
 OA211x2_ASAP7_75t_R _24819_ (.A1(_13387_),
    .A2(_18147_),
    .B(_06716_),
    .C(_06719_),
    .Y(_17550_));
 OR3x1_ASAP7_75t_R _24820_ (.A(_00682_),
    .B(net295),
    .C(_13574_),
    .Y(_06720_));
 OAI21x1_ASAP7_75t_R _24821_ (.A1(_13576_),
    .A2(_18158_),
    .B(_06720_),
    .Y(_17554_));
 AO221x1_ASAP7_75t_R _24822_ (.A1(_13530_),
    .A2(_00686_),
    .B1(_02221_),
    .B2(_13533_),
    .C(net295),
    .Y(_06721_));
 AO221x1_ASAP7_75t_R _24823_ (.A1(_06705_),
    .A2(_13878_),
    .B1(_15266_),
    .B2(_13528_),
    .C(_06721_),
    .Y(_06722_));
 OAI21x1_ASAP7_75t_R _24824_ (.A1(_13387_),
    .A2(_18166_),
    .B(net294),
    .Y(_06723_));
 AO22x1_ASAP7_75t_R _24825_ (.A1(_13781_),
    .A2(_18166_),
    .B1(_06722_),
    .B2(_06723_),
    .Y(_17558_));
 AO221x1_ASAP7_75t_R _24826_ (.A1(_13530_),
    .A2(_00750_),
    .B1(_02219_),
    .B2(_13533_),
    .C(net295),
    .Y(_06724_));
 AO221x1_ASAP7_75t_R _24827_ (.A1(_13528_),
    .A2(_15507_),
    .B1(_15555_),
    .B2(_06705_),
    .C(_06724_),
    .Y(_06725_));
 OAI21x1_ASAP7_75t_R _24828_ (.A1(_13387_),
    .A2(_18177_),
    .B(net294),
    .Y(_06726_));
 AO22x1_ASAP7_75t_R _24829_ (.A1(_13781_),
    .A2(_18177_),
    .B1(_06725_),
    .B2(_06726_),
    .Y(_17562_));
 AOI22x1_ASAP7_75t_R _24830_ (.A1(_13530_),
    .A2(_00783_),
    .B1(_02218_),
    .B2(_13533_),
    .Y(_06727_));
 OA211x2_ASAP7_75t_R _24831_ (.A1(_00284_),
    .A2(_15665_),
    .B(_06727_),
    .C(_13763_),
    .Y(_06728_));
 AO21x1_ASAP7_75t_R _24832_ (.A1(_13528_),
    .A2(_15617_),
    .B(_06728_),
    .Y(_06729_));
 AOI22x1_ASAP7_75t_R _24833_ (.A1(_13781_),
    .A2(_15620_),
    .B1(_06729_),
    .B2(_13576_),
    .Y(_06730_));
 OA21x2_ASAP7_75t_R _24834_ (.A1(_13387_),
    .A2(_15620_),
    .B(_06730_),
    .Y(_16522_));
 OR3x1_ASAP7_75t_R _24835_ (.A(_00816_),
    .B(net294),
    .C(_13574_),
    .Y(_06731_));
 OAI21x1_ASAP7_75t_R _24836_ (.A1(_13576_),
    .A2(_18186_),
    .B(_06731_),
    .Y(_17564_));
 XNOR2x1_ASAP7_75t_R _24837_ (.B(_18197_),
    .Y(_06732_),
    .A(_13387_));
 AO222x2_ASAP7_75t_R _24838_ (.A1(_13530_),
    .A2(_00881_),
    .B1(_02215_),
    .B2(_13533_),
    .C1(_16018_),
    .C2(_06705_),
    .Y(_06733_));
 AO21x1_ASAP7_75t_R _24839_ (.A1(_13528_),
    .A2(_15971_),
    .B(_06733_),
    .Y(_06734_));
 AND2x2_ASAP7_75t_R _24840_ (.A(_13576_),
    .B(_06734_),
    .Y(_06735_));
 AO21x1_ASAP7_75t_R _24841_ (.A1(net295),
    .A2(_06732_),
    .B(_06735_),
    .Y(_17568_));
 OR3x1_ASAP7_75t_R _24842_ (.A(_00946_),
    .B(net295),
    .C(_13574_),
    .Y(_06736_));
 OAI21x1_ASAP7_75t_R _24843_ (.A1(_13576_),
    .A2(_18206_),
    .B(_06736_),
    .Y(_17572_));
 INVx1_ASAP7_75t_R _24844_ (.A(_18211_),
    .Y(_18213_));
 INVx1_ASAP7_75t_R _24845_ (.A(_00979_),
    .Y(_06737_));
 BUFx3_ASAP7_75t_R input31 (.A(data_rdata_i[13]),
    .Y(net31));
 AND3x1_ASAP7_75t_R _24847_ (.A(_06737_),
    .B(_13576_),
    .C(_13533_),
    .Y(_06739_));
 AO21x2_ASAP7_75t_R _24848_ (.A1(net295),
    .A2(_18213_),
    .B(_06739_),
    .Y(_16532_));
 OA21x2_ASAP7_75t_R _24849_ (.A1(_00915_),
    .A2(_16529_),
    .B(_00948_),
    .Y(_06740_));
 OAI21x1_ASAP7_75t_R _24850_ (.A1(_00947_),
    .A2(_06740_),
    .B(_02277_),
    .Y(_16531_));
 XOR2x1_ASAP7_75t_R _24851_ (.A(_13387_),
    .Y(_06741_),
    .B(_18218_));
 AOI22x1_ASAP7_75t_R _24852_ (.A1(_13530_),
    .A2(_01011_),
    .B1(_02211_),
    .B2(_13533_),
    .Y(_06742_));
 OA211x2_ASAP7_75t_R _24853_ (.A1(_00284_),
    .A2(_05849_),
    .B(_06742_),
    .C(_13576_),
    .Y(_06743_));
 INVx1_ASAP7_75t_R _24854_ (.A(_06743_),
    .Y(_06744_));
 AO21x1_ASAP7_75t_R _24855_ (.A1(_13528_),
    .A2(_16433_),
    .B(_06744_),
    .Y(_06745_));
 OA21x2_ASAP7_75t_R _24856_ (.A1(_13576_),
    .A2(_06741_),
    .B(_06745_),
    .Y(_17574_));
 AO221x1_ASAP7_75t_R _24857_ (.A1(_13530_),
    .A2(_01077_),
    .B1(_02209_),
    .B2(_13533_),
    .C(net295),
    .Y(_06746_));
 OAI22x1_ASAP7_75t_R _24858_ (.A1(_13763_),
    .A2(_04667_),
    .B1(_04715_),
    .B2(_00284_),
    .Y(_06747_));
 NOR2x1_ASAP7_75t_R _24859_ (.A(_13781_),
    .B(_18227_),
    .Y(_06748_));
 AO21x1_ASAP7_75t_R _24860_ (.A1(_13387_),
    .A2(_18227_),
    .B(_06748_),
    .Y(_06749_));
 OA21x2_ASAP7_75t_R _24861_ (.A1(_06746_),
    .A2(_06747_),
    .B(_06749_),
    .Y(_17578_));
 INVx1_ASAP7_75t_R _24862_ (.A(_01110_),
    .Y(_06750_));
 AND3x1_ASAP7_75t_R _24863_ (.A(_06750_),
    .B(_13576_),
    .C(_13533_),
    .Y(_06751_));
 AO21x2_ASAP7_75t_R _24864_ (.A1(net295),
    .A2(_04829_),
    .B(_06751_),
    .Y(_16538_));
 OR3x1_ASAP7_75t_R _24865_ (.A(_01078_),
    .B(_01046_),
    .C(_16534_),
    .Y(_06752_));
 NAND2x1_ASAP7_75t_R _24866_ (.A(_05486_),
    .B(_06752_),
    .Y(_16537_));
 AO221x1_ASAP7_75t_R _24867_ (.A1(_13530_),
    .A2(_01142_),
    .B1(_02207_),
    .B2(_13533_),
    .C(net295),
    .Y(_06753_));
 AO221x1_ASAP7_75t_R _24868_ (.A1(_13528_),
    .A2(_04888_),
    .B1(_04935_),
    .B2(_06705_),
    .C(_06753_),
    .Y(_06754_));
 OAI21x1_ASAP7_75t_R _24869_ (.A1(_13387_),
    .A2(_18236_),
    .B(net295),
    .Y(_06755_));
 AO22x1_ASAP7_75t_R _24870_ (.A1(_13781_),
    .A2(_18236_),
    .B1(_06754_),
    .B2(_06755_),
    .Y(_17580_));
 AO221x1_ASAP7_75t_R _24871_ (.A1(_13530_),
    .A2(_01176_),
    .B1(_02206_),
    .B2(_13533_),
    .C(net295),
    .Y(_06756_));
 AOI21x1_ASAP7_75t_R _24872_ (.A1(_13528_),
    .A2(_04996_),
    .B(_06756_),
    .Y(_06757_));
 OA21x2_ASAP7_75t_R _24873_ (.A1(_00284_),
    .A2(_05044_),
    .B(_06757_),
    .Y(_06758_));
 AOI21x1_ASAP7_75t_R _24874_ (.A1(_13781_),
    .A2(_04998_),
    .B(_06758_),
    .Y(_06759_));
 OA21x2_ASAP7_75t_R _24875_ (.A1(_13387_),
    .A2(_04998_),
    .B(_06759_),
    .Y(_16540_));
 NOR2x1_ASAP7_75t_R _24876_ (.A(_00284_),
    .B(_05891_),
    .Y(_06760_));
 AO221x1_ASAP7_75t_R _24877_ (.A1(_13530_),
    .A2(_01208_),
    .B1(_02205_),
    .B2(_13533_),
    .C(_13528_),
    .Y(_06761_));
 OAI22x1_ASAP7_75t_R _24878_ (.A1(_13763_),
    .A2(_05105_),
    .B1(_06760_),
    .B2(_06761_),
    .Y(_06762_));
 AOI22x1_ASAP7_75t_R _24879_ (.A1(_13781_),
    .A2(_05107_),
    .B1(_06762_),
    .B2(_13576_),
    .Y(_06763_));
 OA21x2_ASAP7_75t_R _24880_ (.A1(_13387_),
    .A2(_05107_),
    .B(_06763_),
    .Y(_17582_));
 AO221x1_ASAP7_75t_R _24881_ (.A1(_13530_),
    .A2(_01242_),
    .B1(_02204_),
    .B2(_13533_),
    .C(net295),
    .Y(_06764_));
 AO221x1_ASAP7_75t_R _24882_ (.A1(_13528_),
    .A2(_05213_),
    .B1(_05261_),
    .B2(_06705_),
    .C(_06764_),
    .Y(_06765_));
 NAND2x1_ASAP7_75t_R _24883_ (.A(_13781_),
    .B(_05215_),
    .Y(_06766_));
 OA211x2_ASAP7_75t_R _24884_ (.A1(_13387_),
    .A2(_05215_),
    .B(_06765_),
    .C(_06766_),
    .Y(_16543_));
 NOR2x1_ASAP7_75t_R _24885_ (.A(_00284_),
    .B(_05369_),
    .Y(_06767_));
 AO221x1_ASAP7_75t_R _24886_ (.A1(_13530_),
    .A2(_01274_),
    .B1(_02203_),
    .B2(_13533_),
    .C(_13528_),
    .Y(_06768_));
 OA22x2_ASAP7_75t_R _24887_ (.A1(_13763_),
    .A2(_05323_),
    .B1(_06767_),
    .B2(_06768_),
    .Y(_06769_));
 OAI22x1_ASAP7_75t_R _24888_ (.A1(_13387_),
    .A2(_05325_),
    .B1(_06769_),
    .B2(net295),
    .Y(_06770_));
 AOI21x1_ASAP7_75t_R _24889_ (.A1(_13781_),
    .A2(_05325_),
    .B(_06770_),
    .Y(_17584_));
 AND2x2_ASAP7_75t_R _24890_ (.A(_14376_),
    .B(_05535_),
    .Y(_17591_));
 NAND2x1_ASAP7_75t_R _24891_ (.A(_14319_),
    .B(_05535_),
    .Y(_17593_));
 AND2x2_ASAP7_75t_R _24892_ (.A(_05803_),
    .B(_05928_),
    .Y(_17611_));
 AND2x2_ASAP7_75t_R _24893_ (.A(_05803_),
    .B(_05825_),
    .Y(_17638_));
 INVx1_ASAP7_75t_R _24894_ (.A(_01379_),
    .Y(_16578_));
 INVx1_ASAP7_75t_R _24895_ (.A(_01382_),
    .Y(_16583_));
 AND2x2_ASAP7_75t_R _24896_ (.A(_05803_),
    .B(_05936_),
    .Y(_17694_));
 INVx1_ASAP7_75t_R _24897_ (.A(_01438_),
    .Y(_17726_));
 INVx1_ASAP7_75t_R _24898_ (.A(_05946_),
    .Y(_16774_));
 AND2x2_ASAP7_75t_R _24899_ (.A(_05803_),
    .B(_05901_),
    .Y(_17742_));
 INVx1_ASAP7_75t_R _24900_ (.A(_00020_),
    .Y(_17779_));
 INVx1_ASAP7_75t_R _24901_ (.A(_00042_),
    .Y(_17187_));
 INVx2_ASAP7_75t_R _24902_ (.A(_17049_),
    .Y(_17047_));
 INVx2_ASAP7_75t_R _24903_ (.A(_17095_),
    .Y(_17046_));
 INVx1_ASAP7_75t_R _24904_ (.A(_00046_),
    .Y(_17226_));
 INVx3_ASAP7_75t_R _24905_ (.A(_17179_),
    .Y(_17178_));
 INVx2_ASAP7_75t_R _24906_ (.A(_17399_),
    .Y(_17398_));
 INVx2_ASAP7_75t_R _24907_ (.A(_17424_),
    .Y(_17397_));
 INVx2_ASAP7_75t_R _24908_ (.A(_17471_),
    .Y(_17470_));
 INVx1_ASAP7_75t_R _24909_ (.A(_15407_),
    .Y(_18170_));
 INVx1_ASAP7_75t_R _24910_ (.A(_18177_),
    .Y(_18175_));
 INVx1_ASAP7_75t_R _24911_ (.A(_18187_),
    .Y(_18185_));
 INVx1_ASAP7_75t_R _24912_ (.A(_18197_),
    .Y(_18195_));
 INVx1_ASAP7_75t_R _24913_ (.A(_16137_),
    .Y(_18200_));
 INVx1_ASAP7_75t_R _24914_ (.A(_16480_),
    .Y(_18215_));
 NOR2x1_ASAP7_75t_R _24915_ (.A(_17534_),
    .B(_06664_),
    .Y(_17533_));
 INVx1_ASAP7_75t_R _24916_ (.A(_00243_),
    .Y(_18356_));
 OR2x6_ASAP7_75t_R _24917_ (.A(_06312_),
    .B(_06516_),
    .Y(_06771_));
 BUFx3_ASAP7_75t_R input30 (.A(data_rdata_i[12]),
    .Y(net30));
 BUFx3_ASAP7_75t_R input29 (.A(data_rdata_i[11]),
    .Y(net29));
 INVx1_ASAP7_75t_R _24920_ (.A(_06771_),
    .Y(_18386_));
 XNOR2x1_ASAP7_75t_R _24921_ (.B(_13954_),
    .Y(_06774_),
    .A(_13387_));
 AO22x1_ASAP7_75t_R _24922_ (.A1(_13530_),
    .A2(_00663_),
    .B1(_01450_),
    .B2(_13533_),
    .Y(_06775_));
 OAI22x1_ASAP7_75t_R _24923_ (.A1(_13763_),
    .A2(_13943_),
    .B1(_14684_),
    .B2(_00284_),
    .Y(_06776_));
 OA21x2_ASAP7_75t_R _24924_ (.A1(_06775_),
    .A2(_06776_),
    .B(_13576_),
    .Y(_06777_));
 AO21x1_ASAP7_75t_R _24925_ (.A1(net294),
    .A2(_06774_),
    .B(_06777_),
    .Y(_17541_));
 INVx1_ASAP7_75t_R _24926_ (.A(_14822_),
    .Y(_18128_));
 AND3x1_ASAP7_75t_R _24927_ (.A(_06699_),
    .B(_13576_),
    .C(_13533_),
    .Y(_06778_));
 AO21x1_ASAP7_75t_R _24928_ (.A1(net294),
    .A2(_18128_),
    .B(_06778_),
    .Y(_17545_));
 OR3x1_ASAP7_75t_R _24929_ (.A(_00672_),
    .B(net294),
    .C(_13574_),
    .Y(_06779_));
 OAI21x1_ASAP7_75t_R _24930_ (.A1(_13576_),
    .A2(_18138_),
    .B(_06779_),
    .Y(_17549_));
 OR3x1_ASAP7_75t_R _24931_ (.A(_00674_),
    .B(net294),
    .C(_13574_),
    .Y(_06780_));
 OAI21x1_ASAP7_75t_R _24932_ (.A1(_13576_),
    .A2(_18143_),
    .B(_06780_),
    .Y(_16511_));
 OR3x1_ASAP7_75t_R _24933_ (.A(_00677_),
    .B(net294),
    .C(_13574_),
    .Y(_06781_));
 OAI21x1_ASAP7_75t_R _24934_ (.A1(_13576_),
    .A2(_18148_),
    .B(_06781_),
    .Y(_17551_));
 AO221x1_ASAP7_75t_R _24935_ (.A1(_13530_),
    .A2(_00682_),
    .B1(_01442_),
    .B2(_13533_),
    .C(net295),
    .Y(_06782_));
 AOI21x1_ASAP7_75t_R _24936_ (.A1(_13528_),
    .A2(_05672_),
    .B(_06782_),
    .Y(_06783_));
 OAI21x1_ASAP7_75t_R _24937_ (.A1(_00284_),
    .A2(_15157_),
    .B(_06783_),
    .Y(_06784_));
 NAND2x1_ASAP7_75t_R _24938_ (.A(_13781_),
    .B(_18157_),
    .Y(_06785_));
 OA211x2_ASAP7_75t_R _24939_ (.A1(_13387_),
    .A2(_18157_),
    .B(_06784_),
    .C(_06785_),
    .Y(_17555_));
 OR3x1_ASAP7_75t_R _24940_ (.A(_00686_),
    .B(net295),
    .C(_13574_),
    .Y(_06786_));
 OAI21x1_ASAP7_75t_R _24941_ (.A1(_13576_),
    .A2(_18167_),
    .B(_06786_),
    .Y(_17559_));
 INVx2_ASAP7_75t_R _24942_ (.A(_15556_),
    .Y(_18178_));
 INVx2_ASAP7_75t_R _24943_ (.A(_00750_),
    .Y(_06787_));
 AND3x1_ASAP7_75t_R _24944_ (.A(_06787_),
    .B(_13576_),
    .C(_13533_),
    .Y(_06788_));
 AO21x1_ASAP7_75t_R _24945_ (.A1(net294),
    .A2(_18178_),
    .B(_06788_),
    .Y(_17563_));
 INVx1_ASAP7_75t_R _24946_ (.A(_00783_),
    .Y(_06789_));
 AND3x1_ASAP7_75t_R _24947_ (.A(_06789_),
    .B(_13576_),
    .C(_13533_),
    .Y(_06790_));
 AO21x1_ASAP7_75t_R _24948_ (.A1(net294),
    .A2(_15668_),
    .B(_06790_),
    .Y(_16524_));
 XNOR2x1_ASAP7_75t_R _24949_ (.B(_18187_),
    .Y(_06791_),
    .A(_13387_));
 AND2x2_ASAP7_75t_R _24950_ (.A(_15754_),
    .B(_15777_),
    .Y(_06792_));
 NOR2x1_ASAP7_75t_R _24951_ (.A(_00284_),
    .B(_06792_),
    .Y(_06793_));
 AO22x1_ASAP7_75t_R _24952_ (.A1(_13530_),
    .A2(_00816_),
    .B1(_02217_),
    .B2(_13533_),
    .Y(_06794_));
 OR3x1_ASAP7_75t_R _24953_ (.A(_13528_),
    .B(_06793_),
    .C(_06794_),
    .Y(_06795_));
 OA211x2_ASAP7_75t_R _24954_ (.A1(_13763_),
    .A2(_15731_),
    .B(_06795_),
    .C(_13576_),
    .Y(_06796_));
 AO21x1_ASAP7_75t_R _24955_ (.A1(net295),
    .A2(_06791_),
    .B(_06796_),
    .Y(_17565_));
 OR3x1_ASAP7_75t_R _24956_ (.A(_00881_),
    .B(net295),
    .C(_13574_),
    .Y(_06797_));
 OAI21x1_ASAP7_75t_R _24957_ (.A1(_13576_),
    .A2(_18196_),
    .B(_06797_),
    .Y(_17569_));
 XOR2x1_ASAP7_75t_R _24958_ (.A(_13387_),
    .Y(_06798_),
    .B(_18205_));
 INVx1_ASAP7_75t_R _24959_ (.A(_16256_),
    .Y(_06799_));
 AO22x1_ASAP7_75t_R _24960_ (.A1(_13528_),
    .A2(_16205_),
    .B1(_06799_),
    .B2(_06705_),
    .Y(_06800_));
 AO221x1_ASAP7_75t_R _24961_ (.A1(_13530_),
    .A2(_00946_),
    .B1(_02213_),
    .B2(_13533_),
    .C(net295),
    .Y(_06801_));
 OA22x2_ASAP7_75t_R _24962_ (.A1(_13576_),
    .A2(_06798_),
    .B1(_06800_),
    .B2(_06801_),
    .Y(_17573_));
 AO221x1_ASAP7_75t_R _24963_ (.A1(_13530_),
    .A2(_00979_),
    .B1(_02212_),
    .B2(_13533_),
    .C(net295),
    .Y(_06802_));
 NOR2x1_ASAP7_75t_R _24964_ (.A(_00284_),
    .B(_16372_),
    .Y(_06803_));
 AO21x1_ASAP7_75t_R _24965_ (.A1(_13528_),
    .A2(_16324_),
    .B(_06803_),
    .Y(_06804_));
 OAI22x1_ASAP7_75t_R _24966_ (.A1(_13387_),
    .A2(_16326_),
    .B1(_06802_),
    .B2(_06804_),
    .Y(_06805_));
 AOI21x1_ASAP7_75t_R _24967_ (.A1(_13781_),
    .A2(_16326_),
    .B(_06805_),
    .Y(_16533_));
 INVx1_ASAP7_75t_R _24968_ (.A(_01011_),
    .Y(_06806_));
 AND3x1_ASAP7_75t_R _24969_ (.A(_06806_),
    .B(_13576_),
    .C(_13533_),
    .Y(_06807_));
 AO21x1_ASAP7_75t_R _24970_ (.A1(net295),
    .A2(_18215_),
    .B(_06807_),
    .Y(_17575_));
 OR3x1_ASAP7_75t_R _24971_ (.A(_01077_),
    .B(net295),
    .C(_13574_),
    .Y(_06808_));
 OAI21x1_ASAP7_75t_R _24972_ (.A1(_13576_),
    .A2(_18226_),
    .B(_06808_),
    .Y(_17579_));
 NOR2x1_ASAP7_75t_R _24973_ (.A(_00284_),
    .B(_04828_),
    .Y(_06809_));
 AO221x1_ASAP7_75t_R _24974_ (.A1(_13530_),
    .A2(_01110_),
    .B1(_02208_),
    .B2(_13533_),
    .C(_13528_),
    .Y(_06810_));
 OA22x2_ASAP7_75t_R _24975_ (.A1(_13763_),
    .A2(_04780_),
    .B1(_06809_),
    .B2(_06810_),
    .Y(_06811_));
 OAI22x1_ASAP7_75t_R _24976_ (.A1(_13387_),
    .A2(_04782_),
    .B1(_06811_),
    .B2(net295),
    .Y(_06812_));
 AOI21x1_ASAP7_75t_R _24977_ (.A1(_13781_),
    .A2(_04782_),
    .B(_06812_),
    .Y(_16539_));
 INVx1_ASAP7_75t_R _24978_ (.A(_01142_),
    .Y(_06813_));
 AND3x1_ASAP7_75t_R _24979_ (.A(_06813_),
    .B(_13576_),
    .C(_13533_),
    .Y(_06814_));
 AO21x1_ASAP7_75t_R _24980_ (.A1(net295),
    .A2(_18235_),
    .B(_06814_),
    .Y(_17581_));
 INVx1_ASAP7_75t_R _24981_ (.A(_01176_),
    .Y(_06815_));
 AND3x1_ASAP7_75t_R _24982_ (.A(_06815_),
    .B(_13576_),
    .C(_13533_),
    .Y(_06816_));
 AO21x1_ASAP7_75t_R _24983_ (.A1(net295),
    .A2(_05045_),
    .B(_06816_),
    .Y(_16542_));
 OA21x2_ASAP7_75t_R _24984_ (.A1(_16534_),
    .A2(_05495_),
    .B(_05489_),
    .Y(_06817_));
 INVx1_ASAP7_75t_R _24985_ (.A(_06817_),
    .Y(_16541_));
 OR3x1_ASAP7_75t_R _24986_ (.A(_01208_),
    .B(net294),
    .C(_13574_),
    .Y(_06818_));
 OAI21x1_ASAP7_75t_R _24987_ (.A1(_13576_),
    .A2(_18246_),
    .B(_06818_),
    .Y(_17583_));
 OR3x1_ASAP7_75t_R _24988_ (.A(_01242_),
    .B(net295),
    .C(_13574_),
    .Y(_06819_));
 OAI21x1_ASAP7_75t_R _24989_ (.A1(_13576_),
    .A2(_18251_),
    .B(_06819_),
    .Y(_16544_));
 OA21x2_ASAP7_75t_R _24990_ (.A1(_01177_),
    .A2(_06817_),
    .B(_01210_),
    .Y(_06820_));
 OAI21x1_ASAP7_75t_R _24991_ (.A1(_01209_),
    .A2(_06820_),
    .B(_02281_),
    .Y(_16545_));
 OR3x1_ASAP7_75t_R _24992_ (.A(_01274_),
    .B(net295),
    .C(_13574_),
    .Y(_06821_));
 OAI21x1_ASAP7_75t_R _24993_ (.A1(_13576_),
    .A2(_18256_),
    .B(_06821_),
    .Y(_17585_));
 BUFx3_ASAP7_75t_R input28 (.A(data_rdata_i[10]),
    .Y(net28));
 BUFx2_ASAP7_75t_R input27 (.A(data_rdata_i[0]),
    .Y(net27));
 AND2x2_ASAP7_75t_R _24996_ (.A(_05796_),
    .B(_05815_),
    .Y(_17612_));
 AND2x2_ASAP7_75t_R _24997_ (.A(_05812_),
    .B(_05815_),
    .Y(_17639_));
 INVx1_ASAP7_75t_R _24998_ (.A(_01395_),
    .Y(_16582_));
 INVx1_ASAP7_75t_R _24999_ (.A(_05939_),
    .Y(_16605_));
 OA21x2_ASAP7_75t_R _25000_ (.A1(_01398_),
    .A2(_05939_),
    .B(_01411_),
    .Y(_06823_));
 OAI21x1_ASAP7_75t_R _25001_ (.A1(_01410_),
    .A2(_06823_),
    .B(_02322_),
    .Y(_16653_));
 AND2x2_ASAP7_75t_R _25002_ (.A(_05815_),
    .B(_05855_),
    .Y(_17695_));
 AOI21x1_ASAP7_75t_R _25003_ (.A1(_02326_),
    .A2(_05943_),
    .B(_05941_),
    .Y(_16707_));
 INVx1_ASAP7_75t_R _25004_ (.A(_01433_),
    .Y(_17709_));
 INVx1_ASAP7_75t_R _25005_ (.A(_01439_),
    .Y(_17729_));
 AND2x2_ASAP7_75t_R _25006_ (.A(_05815_),
    .B(_05875_),
    .Y(_17743_));
 OA21x2_ASAP7_75t_R _25007_ (.A1(_00009_),
    .A2(_05946_),
    .B(_00016_),
    .Y(_06824_));
 OAI21x1_ASAP7_75t_R _25008_ (.A1(_00015_),
    .A2(_06824_),
    .B(_02336_),
    .Y(_16857_));
 INVx1_ASAP7_75t_R _25009_ (.A(_00026_),
    .Y(_16910_));
 INVx1_ASAP7_75t_R _25010_ (.A(_00028_),
    .Y(_16949_));
 OR3x1_ASAP7_75t_R _25011_ (.A(_00031_),
    .B(_05951_),
    .C(_05953_),
    .Y(_06825_));
 NAND2x1_ASAP7_75t_R _25012_ (.A(_02344_),
    .B(_06825_),
    .Y(_17058_));
 NAND2x1_ASAP7_75t_R _25013_ (.A(_02347_),
    .B(_05957_),
    .Y(_17146_));
 INVx1_ASAP7_75t_R _25014_ (.A(_17227_),
    .Y(_17177_));
 INVx1_ASAP7_75t_R _25015_ (.A(_00047_),
    .Y(_17186_));
 INVx1_ASAP7_75t_R _25016_ (.A(_05961_),
    .Y(_17237_));
 INVx1_ASAP7_75t_R _25017_ (.A(_00050_),
    .Y(_17225_));
 OA21x2_ASAP7_75t_R _25018_ (.A1(_00049_),
    .A2(_05961_),
    .B(_00053_),
    .Y(_06826_));
 OAI21x1_ASAP7_75t_R _25019_ (.A1(_00052_),
    .A2(_06826_),
    .B(_02353_),
    .Y(_17315_));
 AO21x1_ASAP7_75t_R _25020_ (.A1(_00056_),
    .A2(_05965_),
    .B(_00055_),
    .Y(_06827_));
 NAND2x1_ASAP7_75t_R _25021_ (.A(_02354_),
    .B(_06827_),
    .Y(_17381_));
 INVx1_ASAP7_75t_R _25022_ (.A(_05969_),
    .Y(_17439_));
 INVx1_ASAP7_75t_R _25023_ (.A(_05971_),
    .Y(_17491_));
 INVx1_ASAP7_75t_R _25024_ (.A(_17500_),
    .Y(_17469_));
 INVx1_ASAP7_75t_R _25025_ (.A(_17507_),
    .Y(_17477_));
 INVx1_ASAP7_75t_R _25026_ (.A(_14688_),
    .Y(_18117_));
 INVx1_ASAP7_75t_R _25027_ (.A(_18133_),
    .Y(_18131_));
 INVx1_ASAP7_75t_R _25028_ (.A(_18143_),
    .Y(_18141_));
 INVx1_ASAP7_75t_R _25029_ (.A(_18148_),
    .Y(_18146_));
 INVx1_ASAP7_75t_R _25030_ (.A(_14576_),
    .Y(_18163_));
 INVx1_ASAP7_75t_R _25031_ (.A(_18166_),
    .Y(_18168_));
 INVx1_ASAP7_75t_R _25032_ (.A(_15897_),
    .Y(_18193_));
 INVx1_ASAP7_75t_R _25033_ (.A(_18236_),
    .Y(_18238_));
 INVx1_ASAP7_75t_R _25034_ (.A(_01718_),
    .Y(_06828_));
 AO32x1_ASAP7_75t_R _25035_ (.A1(net145),
    .A2(_06189_),
    .A3(_06191_),
    .B1(_06262_),
    .B2(_06828_),
    .Y(_02647_));
 NOR2x1_ASAP7_75t_R _25036_ (.A(_05709_),
    .B(_06170_),
    .Y(_06829_));
 AND5x1_ASAP7_75t_R _25037_ (.A(_13227_),
    .B(_01740_),
    .C(_01741_),
    .D(_05557_),
    .E(_06598_),
    .Y(_06830_));
 AND3x1_ASAP7_75t_R _25038_ (.A(_13772_),
    .B(_05720_),
    .C(_06830_),
    .Y(_06831_));
 AND3x2_ASAP7_75t_R _25039_ (.A(_01312_),
    .B(_01721_),
    .C(_06831_),
    .Y(_06832_));
 OAI21x1_ASAP7_75t_R _25040_ (.A1(net60),
    .A2(_06611_),
    .B(_01311_),
    .Y(_06833_));
 AO21x1_ASAP7_75t_R _25041_ (.A1(_06829_),
    .A2(_06832_),
    .B(_06833_),
    .Y(_06834_));
 OA211x2_ASAP7_75t_R _25042_ (.A1(_05711_),
    .A2(_06278_),
    .B(_06834_),
    .C(_05527_),
    .Y(_06835_));
 AND2x2_ASAP7_75t_R _25043_ (.A(_06180_),
    .B(_01716_),
    .Y(_06836_));
 AO21x1_ASAP7_75t_R _25044_ (.A1(_01714_),
    .A2(_01717_),
    .B(_06836_),
    .Y(_06837_));
 AND2x2_ASAP7_75t_R _25045_ (.A(_01717_),
    .B(_06833_),
    .Y(_06838_));
 AO22x1_ASAP7_75t_R _25046_ (.A1(_14581_),
    .A2(_06188_),
    .B1(_06838_),
    .B2(_01716_),
    .Y(_06839_));
 AND3x2_ASAP7_75t_R _25047_ (.A(_14580_),
    .B(_06555_),
    .C(_06651_),
    .Y(_06840_));
 AO221x1_ASAP7_75t_R _25048_ (.A1(_01715_),
    .A2(_06837_),
    .B1(_06839_),
    .B2(_01714_),
    .C(_06840_),
    .Y(_06841_));
 OA21x2_ASAP7_75t_R _25049_ (.A1(_05527_),
    .A2(_05726_),
    .B(_06604_),
    .Y(_06842_));
 AND2x2_ASAP7_75t_R _25050_ (.A(_06594_),
    .B(_06612_),
    .Y(_06843_));
 NOR2x1_ASAP7_75t_R _25051_ (.A(_06266_),
    .B(_06843_),
    .Y(_06844_));
 AND2x2_ASAP7_75t_R _25052_ (.A(_06842_),
    .B(_06844_),
    .Y(_06845_));
 OR4x2_ASAP7_75t_R _25053_ (.A(_06180_),
    .B(_01715_),
    .C(_01716_),
    .D(_14580_),
    .Y(_06846_));
 AND3x1_ASAP7_75t_R _25054_ (.A(_06846_),
    .B(_06556_),
    .C(_06607_),
    .Y(_06847_));
 NAND2x1_ASAP7_75t_R _25055_ (.A(_14583_),
    .B(_06838_),
    .Y(_06848_));
 OA33x2_ASAP7_75t_R _25056_ (.A1(_06835_),
    .A2(_06841_),
    .A3(_06845_),
    .B1(_06847_),
    .B2(_06848_),
    .B3(_06610_),
    .Y(_02648_));
 AOI21x1_ASAP7_75t_R _25057_ (.A1(_06594_),
    .A2(_06610_),
    .B(_05526_),
    .Y(_06849_));
 OAI21x1_ASAP7_75t_R _25058_ (.A1(_06843_),
    .A2(_06849_),
    .B(_06842_),
    .Y(_06850_));
 AND3x1_ASAP7_75t_R _25059_ (.A(_14583_),
    .B(_06610_),
    .C(_06833_),
    .Y(_06851_));
 OA21x2_ASAP7_75t_R _25060_ (.A1(_06555_),
    .A2(_06851_),
    .B(_01717_),
    .Y(_06852_));
 INVx1_ASAP7_75t_R _25061_ (.A(_05711_),
    .Y(_06853_));
 AO21x1_ASAP7_75t_R _25062_ (.A1(_06602_),
    .A2(_06610_),
    .B(_06853_),
    .Y(_06854_));
 AND3x1_ASAP7_75t_R _25063_ (.A(_06304_),
    .B(_06834_),
    .C(_06854_),
    .Y(_06855_));
 OR3x1_ASAP7_75t_R _25064_ (.A(_06840_),
    .B(_06852_),
    .C(_06855_),
    .Y(_06856_));
 AO21x1_ASAP7_75t_R _25065_ (.A1(_14584_),
    .A2(_06850_),
    .B(_06856_),
    .Y(_02649_));
 AO21x1_ASAP7_75t_R _25066_ (.A1(_01714_),
    .A2(_14580_),
    .B(_06836_),
    .Y(_06857_));
 AND3x1_ASAP7_75t_R _25067_ (.A(_14581_),
    .B(_01716_),
    .C(_06838_),
    .Y(_06858_));
 OA21x2_ASAP7_75t_R _25068_ (.A1(_06188_),
    .A2(_06858_),
    .B(_01714_),
    .Y(_06859_));
 AO221x1_ASAP7_75t_R _25069_ (.A1(_06177_),
    .A2(_06835_),
    .B1(_06857_),
    .B2(_01715_),
    .C(_06859_),
    .Y(_06860_));
 INVx1_ASAP7_75t_R _25070_ (.A(_06860_),
    .Y(_06861_));
 AO21x1_ASAP7_75t_R _25071_ (.A1(_06843_),
    .A2(_06842_),
    .B(_06266_),
    .Y(_06862_));
 AOI21x1_ASAP7_75t_R _25072_ (.A1(_06861_),
    .A2(_06862_),
    .B(_06840_),
    .Y(_02650_));
 AO21x1_ASAP7_75t_R _25073_ (.A1(_06594_),
    .A2(_06842_),
    .B(_01717_),
    .Y(_06863_));
 NAND2x1_ASAP7_75t_R _25074_ (.A(_06177_),
    .B(_06834_),
    .Y(_06864_));
 AO32x1_ASAP7_75t_R _25075_ (.A1(_14583_),
    .A2(_06612_),
    .A3(_06863_),
    .B1(_06864_),
    .B2(_05527_),
    .Y(_02651_));
 OR3x1_ASAP7_75t_R _25076_ (.A(_14615_),
    .B(_06162_),
    .C(_06631_),
    .Y(_06865_));
 AO21x1_ASAP7_75t_R _25077_ (.A1(_14615_),
    .A2(_06586_),
    .B(_06585_),
    .Y(_06866_));
 AO21x1_ASAP7_75t_R _25078_ (.A1(_01713_),
    .A2(_06865_),
    .B(_06866_),
    .Y(_06867_));
 INVx1_ASAP7_75t_R _25079_ (.A(_06585_),
    .Y(_06868_));
 AOI21x1_ASAP7_75t_R _25080_ (.A1(_14585_),
    .A2(_06868_),
    .B(_01713_),
    .Y(_06869_));
 AO21x1_ASAP7_75t_R _25081_ (.A1(_05729_),
    .A2(_06867_),
    .B(_06869_),
    .Y(_02652_));
 INVx2_ASAP7_75t_R _25082_ (.A(_02034_),
    .Y(_06870_));
 OR3x1_ASAP7_75t_R _25083_ (.A(_05677_),
    .B(_01717_),
    .C(_06170_),
    .Y(_06871_));
 OAI21x1_ASAP7_75t_R _25084_ (.A1(_14580_),
    .A2(_06184_),
    .B(_06871_),
    .Y(_06872_));
 NAND2x2_ASAP7_75t_R _25085_ (.A(_06327_),
    .B(_06872_),
    .Y(_06873_));
 BUFx4f_ASAP7_75t_R input26 (.A(data_gnt_i),
    .Y(net26));
 AO32x1_ASAP7_75t_R _25087_ (.A1(_01717_),
    .A2(_06870_),
    .A3(_06327_),
    .B1(_06873_),
    .B2(_01712_),
    .Y(_06875_));
 INVx1_ASAP7_75t_R _25088_ (.A(_06875_),
    .Y(_02653_));
 OR3x4_ASAP7_75t_R _25089_ (.A(_01714_),
    .B(_14580_),
    .C(_06181_),
    .Y(_06876_));
 INVx1_ASAP7_75t_R _25090_ (.A(_06876_),
    .Y(_06877_));
 BUFx2_ASAP7_75t_R input25 (.A(data_err_i),
    .Y(net25));
 INVx1_ASAP7_75t_R _25092_ (.A(_01711_),
    .Y(_06879_));
 AO32x1_ASAP7_75t_R _25093_ (.A1(net60),
    .A2(_02034_),
    .A3(_06877_),
    .B1(_06873_),
    .B2(_06879_),
    .Y(_02654_));
 INVx4_ASAP7_75t_R _25094_ (.A(_06873_),
    .Y(_06880_));
 OAI22x1_ASAP7_75t_R _25095_ (.A1(_02034_),
    .A2(_06876_),
    .B1(_06880_),
    .B2(_01726_),
    .Y(_02655_));
 AND2x4_ASAP7_75t_R _25096_ (.A(_00187_),
    .B(_00191_),
    .Y(_06881_));
 AND2x2_ASAP7_75t_R _25097_ (.A(_13652_),
    .B(_00184_),
    .Y(_06882_));
 AND4x1_ASAP7_75t_R _25098_ (.A(_05523_),
    .B(_01316_),
    .C(_01607_),
    .D(_05522_),
    .Y(_06883_));
 OA211x2_ASAP7_75t_R _25099_ (.A1(_14084_),
    .A2(_05588_),
    .B(_05601_),
    .C(_14140_),
    .Y(_06884_));
 BUFx2_ASAP7_75t_R input24 (.A(boot_addr_i[9]),
    .Y(net24));
 OA211x2_ASAP7_75t_R _25101_ (.A1(_14084_),
    .A2(_05588_),
    .B(_05661_),
    .C(_14140_),
    .Y(_06886_));
 BUFx2_ASAP7_75t_R input23 (.A(boot_addr_i[8]),
    .Y(net23));
 AND4x1_ASAP7_75t_R _25103_ (.A(_13369_),
    .B(_05531_),
    .C(_05534_),
    .D(_05535_),
    .Y(_06888_));
 AND4x2_ASAP7_75t_R _25104_ (.A(_13301_),
    .B(net289),
    .C(_13954_),
    .D(_05542_),
    .Y(_06889_));
 BUFx2_ASAP7_75t_R input22 (.A(boot_addr_i[31]),
    .Y(net22));
 AND4x2_ASAP7_75t_R _25106_ (.A(_18162_),
    .B(_05609_),
    .C(_06888_),
    .D(_06889_),
    .Y(_06891_));
 AND5x2_ASAP7_75t_R _25107_ (.A(_14084_),
    .B(_14497_),
    .C(_05571_),
    .D(_05606_),
    .E(_06888_),
    .Y(_06892_));
 AND5x1_ASAP7_75t_R _25108_ (.A(_13306_),
    .B(_14138_),
    .C(_14497_),
    .D(_05536_),
    .E(_05606_),
    .Y(_06893_));
 OAI21x1_ASAP7_75t_R _25109_ (.A1(_13954_),
    .A2(_14026_),
    .B(_05616_),
    .Y(_06894_));
 AO32x1_ASAP7_75t_R _25110_ (.A1(_05677_),
    .A2(_05624_),
    .A3(_06892_),
    .B1(_06893_),
    .B2(_06894_),
    .Y(_06895_));
 OR4x1_ASAP7_75t_R _25111_ (.A(_06884_),
    .B(_06886_),
    .C(_06891_),
    .D(_06895_),
    .Y(_06896_));
 AND3x1_ASAP7_75t_R _25112_ (.A(_14083_),
    .B(_14140_),
    .C(_18142_),
    .Y(_06897_));
 OA211x2_ASAP7_75t_R _25113_ (.A1(_05558_),
    .A2(_06897_),
    .B(_06889_),
    .C(_05576_),
    .Y(_06898_));
 OR3x1_ASAP7_75t_R _25114_ (.A(_13954_),
    .B(_14026_),
    .C(_14084_),
    .Y(_06899_));
 OA211x2_ASAP7_75t_R _25115_ (.A1(_05541_),
    .A2(_06899_),
    .B(_14139_),
    .C(_05538_),
    .Y(_06900_));
 NAND2x1_ASAP7_75t_R _25116_ (.A(_05542_),
    .B(_05611_),
    .Y(_06901_));
 NOR3x1_ASAP7_75t_R _25117_ (.A(_18162_),
    .B(_05655_),
    .C(_06901_),
    .Y(_06902_));
 NOR2x1_ASAP7_75t_R _25118_ (.A(_14084_),
    .B(_05571_),
    .Y(_06903_));
 AND4x1_ASAP7_75t_R _25119_ (.A(_13301_),
    .B(_13955_),
    .C(_06902_),
    .D(_06903_),
    .Y(_06904_));
 OR4x1_ASAP7_75t_R _25120_ (.A(_05628_),
    .B(_06898_),
    .C(_06900_),
    .D(_06904_),
    .Y(_06905_));
 AND4x2_ASAP7_75t_R _25121_ (.A(_13301_),
    .B(_13658_),
    .C(_13955_),
    .D(_05542_),
    .Y(_06906_));
 AO32x1_ASAP7_75t_R _25122_ (.A1(_14083_),
    .A2(_14139_),
    .A3(_05582_),
    .B1(_05631_),
    .B2(_06906_),
    .Y(_06907_));
 OA21x2_ASAP7_75t_R _25123_ (.A1(_13954_),
    .A2(_05581_),
    .B(_05535_),
    .Y(_06908_));
 OR4x1_ASAP7_75t_R _25124_ (.A(_13302_),
    .B(net289),
    .C(_13955_),
    .D(_05560_),
    .Y(_06909_));
 OA21x2_ASAP7_75t_R _25125_ (.A1(_14084_),
    .A2(_14139_),
    .B(_05535_),
    .Y(_06910_));
 NAND2x2_ASAP7_75t_R _25126_ (.A(_05579_),
    .B(_05576_),
    .Y(_06911_));
 AOI211x1_ASAP7_75t_R _25127_ (.A1(_06908_),
    .A2(_06909_),
    .B(_06910_),
    .C(_06911_),
    .Y(_06912_));
 AO21x1_ASAP7_75t_R _25128_ (.A1(_05538_),
    .A2(_06907_),
    .B(_06912_),
    .Y(_06913_));
 INVx1_ASAP7_75t_R _25129_ (.A(_05703_),
    .Y(_06914_));
 OA31x2_ASAP7_75t_R _25130_ (.A1(_06896_),
    .A2(_06905_),
    .A3(_06913_),
    .B1(_06914_),
    .Y(_06915_));
 INVx1_ASAP7_75t_R _25131_ (.A(_05729_),
    .Y(_06916_));
 OA211x2_ASAP7_75t_R _25132_ (.A1(_13547_),
    .A2(_05557_),
    .B(_13250_),
    .C(_13257_),
    .Y(_06917_));
 OR3x1_ASAP7_75t_R _25133_ (.A(_06916_),
    .B(_06585_),
    .C(_06917_),
    .Y(_06918_));
 INVx1_ASAP7_75t_R _25134_ (.A(_06918_),
    .Y(_06919_));
 OA21x2_ASAP7_75t_R _25135_ (.A1(_05558_),
    .A2(_06915_),
    .B(_06919_),
    .Y(_06920_));
 BUFx2_ASAP7_75t_R input21 (.A(boot_addr_i[30]),
    .Y(net21));
 OR2x4_ASAP7_75t_R _25137_ (.A(_06883_),
    .B(_06920_),
    .Y(_06922_));
 AND3x2_ASAP7_75t_R _25138_ (.A(_00194_),
    .B(_06882_),
    .C(_06922_),
    .Y(_06923_));
 AND2x6_ASAP7_75t_R _25139_ (.A(_06881_),
    .B(_06923_),
    .Y(_06924_));
 BUFx2_ASAP7_75t_R input20 (.A(boot_addr_i[29]),
    .Y(net20));
 BUFx2_ASAP7_75t_R input19 (.A(boot_addr_i[28]),
    .Y(net19));
 OA31x2_ASAP7_75t_R _25142_ (.A1(_02357_),
    .A2(_13954_),
    .A3(_14026_),
    .B1(_13228_),
    .Y(_06927_));
 XNOR2x2_ASAP7_75t_R _25143_ (.A(_14084_),
    .B(_06927_),
    .Y(_06928_));
 BUFx2_ASAP7_75t_R input18 (.A(boot_addr_i[27]),
    .Y(net18));
 BUFx2_ASAP7_75t_R input17 (.A(boot_addr_i[26]),
    .Y(net17));
 AND2x2_ASAP7_75t_R _25146_ (.A(_02358_),
    .B(_13228_),
    .Y(_06931_));
 XNOR2x2_ASAP7_75t_R _25147_ (.A(_14026_),
    .B(_06931_),
    .Y(_06932_));
 BUFx2_ASAP7_75t_R input16 (.A(boot_addr_i[25]),
    .Y(net16));
 NAND2x1_ASAP7_75t_R _25149_ (.A(_00073_),
    .B(_13228_),
    .Y(_06934_));
 OAI21x1_ASAP7_75t_R _25150_ (.A1(_13228_),
    .A2(_13954_),
    .B(_06934_),
    .Y(_06935_));
 BUFx2_ASAP7_75t_R input15 (.A(boot_addr_i[24]),
    .Y(net15));
 BUFx2_ASAP7_75t_R input14 (.A(boot_addr_i[23]),
    .Y(net14));
 AND2x2_ASAP7_75t_R _25153_ (.A(_00072_),
    .B(_13228_),
    .Y(_06938_));
 AO21x2_ASAP7_75t_R _25154_ (.A1(_13328_),
    .A2(_13301_),
    .B(_06938_),
    .Y(_06939_));
 BUFx2_ASAP7_75t_R input13 (.A(boot_addr_i[22]),
    .Y(net13));
 BUFx2_ASAP7_75t_R input12 (.A(boot_addr_i[21]),
    .Y(net12));
 AO21x2_ASAP7_75t_R _25157_ (.A1(_13264_),
    .A2(_13329_),
    .B(_13342_),
    .Y(_06942_));
 AND3x4_ASAP7_75t_R _25158_ (.A(_13364_),
    .B(_13376_),
    .C(_06942_),
    .Y(_06943_));
 BUFx2_ASAP7_75t_R input11 (.A(boot_addr_i[20]),
    .Y(net11));
 BUFx2_ASAP7_75t_R input10 (.A(boot_addr_i[19]),
    .Y(net10));
 NAND3x2_ASAP7_75t_R _25161_ (.B(_13376_),
    .C(_06942_),
    .Y(_06946_),
    .A(_13364_));
 BUFx2_ASAP7_75t_R input9 (.A(boot_addr_i[18]),
    .Y(net9));
 OR3x1_ASAP7_75t_R _25163_ (.A(_14990_),
    .B(_14992_),
    .C(_06946_),
    .Y(_06948_));
 OA21x2_ASAP7_75t_R _25164_ (.A1(_04718_),
    .A2(_06943_),
    .B(_06948_),
    .Y(_06949_));
 BUFx2_ASAP7_75t_R input8 (.A(boot_addr_i[17]),
    .Y(net8));
 BUFx2_ASAP7_75t_R input7 (.A(boot_addr_i[16]),
    .Y(net7));
 NAND2x1_ASAP7_75t_R _25167_ (.A(_18133_),
    .B(_06943_),
    .Y(_06952_));
 AOI21x1_ASAP7_75t_R _25168_ (.A1(_13328_),
    .A2(_13301_),
    .B(_06938_),
    .Y(_06953_));
 OA211x2_ASAP7_75t_R _25169_ (.A1(_18235_),
    .A2(_06943_),
    .B(_06952_),
    .C(net281),
    .Y(_06954_));
 AO21x1_ASAP7_75t_R _25170_ (.A1(_06939_),
    .A2(_06949_),
    .B(_06954_),
    .Y(_06955_));
 NAND2x1_ASAP7_75t_R _25171_ (.A(_14822_),
    .B(_06943_),
    .Y(_06956_));
 OA21x2_ASAP7_75t_R _25172_ (.A1(_05045_),
    .A2(_06943_),
    .B(_06956_),
    .Y(_06957_));
 AND2x2_ASAP7_75t_R _25173_ (.A(_14938_),
    .B(_06943_),
    .Y(_06958_));
 AND2x2_ASAP7_75t_R _25174_ (.A(_04829_),
    .B(_06946_),
    .Y(_06959_));
 OR3x1_ASAP7_75t_R _25175_ (.A(net281),
    .B(_06958_),
    .C(_06959_),
    .Y(_06960_));
 BUFx2_ASAP7_75t_R input6 (.A(boot_addr_i[15]),
    .Y(net6));
 OA211x2_ASAP7_75t_R _25177_ (.A1(_06939_),
    .A2(_06957_),
    .B(_06960_),
    .C(_13658_),
    .Y(_06962_));
 AO21x1_ASAP7_75t_R _25178_ (.A1(net290),
    .A2(_06955_),
    .B(_06962_),
    .Y(_06963_));
 AND2x2_ASAP7_75t_R _25179_ (.A(_06935_),
    .B(_06963_),
    .Y(_06964_));
 BUFx2_ASAP7_75t_R input5 (.A(boot_addr_i[14]),
    .Y(net5));
 BUFx2_ASAP7_75t_R input4 (.A(boot_addr_i[13]),
    .Y(net4));
 AND2x2_ASAP7_75t_R _25182_ (.A(_05478_),
    .B(_06946_),
    .Y(_06967_));
 AO21x1_ASAP7_75t_R _25183_ (.A1(_13777_),
    .A2(_06943_),
    .B(_06967_),
    .Y(_06968_));
 BUFx2_ASAP7_75t_R input3 (.A(boot_addr_i[12]),
    .Y(net3));
 OR2x2_ASAP7_75t_R _25185_ (.A(_05371_),
    .B(_06943_),
    .Y(_06970_));
 OA211x2_ASAP7_75t_R _25186_ (.A1(_13573_),
    .A2(_06946_),
    .B(_06970_),
    .C(net290),
    .Y(_06971_));
 AO21x2_ASAP7_75t_R _25187_ (.A1(_13658_),
    .A2(_06968_),
    .B(_06971_),
    .Y(_06972_));
 BUFx2_ASAP7_75t_R input2 (.A(boot_addr_i[11]),
    .Y(net2));
 BUFx2_ASAP7_75t_R input1 (.A(boot_addr_i[10]),
    .Y(net1));
 NAND2x1_ASAP7_75t_R _25190_ (.A(_18246_),
    .B(_06946_),
    .Y(_06975_));
 OA211x2_ASAP7_75t_R _25191_ (.A1(_14761_),
    .A2(_06946_),
    .B(_06975_),
    .C(net290),
    .Y(_06976_));
 NAND2x1_ASAP7_75t_R _25192_ (.A(_14688_),
    .B(_06943_),
    .Y(_06977_));
 OA211x2_ASAP7_75t_R _25193_ (.A1(_18253_),
    .A2(_06943_),
    .B(_06977_),
    .C(_13658_),
    .Y(_06978_));
 OR3x1_ASAP7_75t_R _25194_ (.A(_06953_),
    .B(_06976_),
    .C(_06978_),
    .Y(_06979_));
 OAI21x1_ASAP7_75t_R _25195_ (.A1(_06939_),
    .A2(_06972_),
    .B(_06979_),
    .Y(_06980_));
 NOR2x2_ASAP7_75t_R _25196_ (.A(_06935_),
    .B(_06980_),
    .Y(_06981_));
 XNOR2x2_ASAP7_75t_R _25197_ (.A(_14025_),
    .B(_06931_),
    .Y(_06982_));
 NAND2x1_ASAP7_75t_R _25198_ (.A(_18148_),
    .B(_06943_),
    .Y(_06983_));
 OR3x1_ASAP7_75t_R _25199_ (.A(_04601_),
    .B(_04602_),
    .C(_06943_),
    .Y(_06984_));
 NAND2x1_ASAP7_75t_R _25200_ (.A(_16480_),
    .B(_06946_),
    .Y(_06985_));
 OA21x2_ASAP7_75t_R _25201_ (.A1(_15104_),
    .A2(_06946_),
    .B(net288),
    .Y(_06986_));
 AO32x1_ASAP7_75t_R _25202_ (.A1(_13658_),
    .A2(_06983_),
    .A3(_06984_),
    .B1(_06985_),
    .B2(_06986_),
    .Y(_06987_));
 AND2x2_ASAP7_75t_R _25203_ (.A(net281),
    .B(_06987_),
    .Y(_06988_));
 NAND2x1_ASAP7_75t_R _25204_ (.A(_14576_),
    .B(_06943_),
    .Y(_06989_));
 OA21x2_ASAP7_75t_R _25205_ (.A1(_16259_),
    .A2(_06943_),
    .B(_06989_),
    .Y(_06990_));
 TAPCELL_ASAP7_75t_R TAP_826 ();
 AND2x2_ASAP7_75t_R _25207_ (.A(_15159_),
    .B(_06943_),
    .Y(_06992_));
 NOR2x1_ASAP7_75t_R _25208_ (.A(_18211_),
    .B(_06943_),
    .Y(_06993_));
 OR3x1_ASAP7_75t_R _25209_ (.A(net288),
    .B(_06992_),
    .C(_06993_),
    .Y(_06994_));
 OA211x2_ASAP7_75t_R _25210_ (.A1(_13658_),
    .A2(_06990_),
    .B(_06994_),
    .C(_06939_),
    .Y(_06995_));
 OA21x2_ASAP7_75t_R _25211_ (.A1(_13228_),
    .A2(_13954_),
    .B(_06934_),
    .Y(_06996_));
 OA21x2_ASAP7_75t_R _25212_ (.A1(_06988_),
    .A2(_06995_),
    .B(_06996_),
    .Y(_06997_));
 NAND2x2_ASAP7_75t_R _25213_ (.A(net288),
    .B(_06946_),
    .Y(_06998_));
 OR2x2_ASAP7_75t_R _25214_ (.A(_15781_),
    .B(_06998_),
    .Y(_06999_));
 NAND2x1_ASAP7_75t_R _25215_ (.A(net288),
    .B(_06943_),
    .Y(_07000_));
 NAND2x2_ASAP7_75t_R _25216_ (.A(_13658_),
    .B(_06946_),
    .Y(_07001_));
 NAND2x2_ASAP7_75t_R _25217_ (.A(_13658_),
    .B(_06943_),
    .Y(_07002_));
 OA222x2_ASAP7_75t_R _25218_ (.A1(_15668_),
    .A2(_07000_),
    .B1(_07001_),
    .B2(_18193_),
    .C1(_07002_),
    .C2(_18178_),
    .Y(_07003_));
 AO21x1_ASAP7_75t_R _25219_ (.A1(_06999_),
    .A2(_07003_),
    .B(net281),
    .Y(_07004_));
 NAND2x1_ASAP7_75t_R _25220_ (.A(_15407_),
    .B(_06943_),
    .Y(_07005_));
 OA211x2_ASAP7_75t_R _25221_ (.A1(_18198_),
    .A2(_06943_),
    .B(_07005_),
    .C(net288),
    .Y(_07006_));
 AND2x2_ASAP7_75t_R _25222_ (.A(_16137_),
    .B(_06946_),
    .Y(_07007_));
 AOI211x1_ASAP7_75t_R _25223_ (.A1(_18167_),
    .A2(_06943_),
    .B(_07007_),
    .C(net288),
    .Y(_07008_));
 OR3x1_ASAP7_75t_R _25224_ (.A(_06939_),
    .B(_07006_),
    .C(_07008_),
    .Y(_07009_));
 AND3x1_ASAP7_75t_R _25225_ (.A(_06935_),
    .B(_07004_),
    .C(_07009_),
    .Y(_07010_));
 OR3x1_ASAP7_75t_R _25226_ (.A(_06982_),
    .B(_06997_),
    .C(_07010_),
    .Y(_07011_));
 OA31x2_ASAP7_75t_R _25227_ (.A1(_06932_),
    .A2(_06964_),
    .A3(_06981_),
    .B1(_07011_),
    .Y(_07012_));
 TAPCELL_ASAP7_75t_R TAP_825 ();
 TAPCELL_ASAP7_75t_R TAP_824 ();
 TAPCELL_ASAP7_75t_R TAP_823 ();
 NAND2x1_ASAP7_75t_R _25231_ (.A(_06996_),
    .B(net281),
    .Y(_07016_));
 OA222x2_ASAP7_75t_R _25232_ (.A1(_18178_),
    .A2(_06998_),
    .B1(_07000_),
    .B2(_18193_),
    .C1(_07001_),
    .C2(_15668_),
    .Y(_07017_));
 OA21x2_ASAP7_75t_R _25233_ (.A1(_15781_),
    .A2(_07002_),
    .B(_07017_),
    .Y(_07018_));
 TAPCELL_ASAP7_75t_R TAP_822 ();
 AND2x2_ASAP7_75t_R _25235_ (.A(_16137_),
    .B(_06943_),
    .Y(_07020_));
 AOI211x1_ASAP7_75t_R _25236_ (.A1(_18167_),
    .A2(_06946_),
    .B(_07020_),
    .C(_13658_),
    .Y(_07021_));
 TAPCELL_ASAP7_75t_R TAP_821 ();
 NAND2x1_ASAP7_75t_R _25238_ (.A(_15407_),
    .B(_06946_),
    .Y(_07023_));
 OA211x2_ASAP7_75t_R _25239_ (.A1(_18198_),
    .A2(_06946_),
    .B(_07023_),
    .C(_13658_),
    .Y(_07024_));
 OR4x1_ASAP7_75t_R _25240_ (.A(_06935_),
    .B(net281),
    .C(_07021_),
    .D(_07024_),
    .Y(_07025_));
 NAND2x1_ASAP7_75t_R _25241_ (.A(_06935_),
    .B(_06939_),
    .Y(_07026_));
 NAND2x1_ASAP7_75t_R _25242_ (.A(_18148_),
    .B(_06946_),
    .Y(_07027_));
 OA211x2_ASAP7_75t_R _25243_ (.A1(_04603_),
    .A2(_06946_),
    .B(_07027_),
    .C(net288),
    .Y(_07028_));
 NAND2x1_ASAP7_75t_R _25244_ (.A(_16480_),
    .B(_06943_),
    .Y(_07029_));
 OA211x2_ASAP7_75t_R _25245_ (.A1(_15104_),
    .A2(_06943_),
    .B(_07029_),
    .C(_13658_),
    .Y(_07030_));
 NAND2x1_ASAP7_75t_R _25246_ (.A(_18211_),
    .B(_06943_),
    .Y(_07031_));
 OR2x2_ASAP7_75t_R _25247_ (.A(_15159_),
    .B(_06943_),
    .Y(_07032_));
 AND3x1_ASAP7_75t_R _25248_ (.A(net288),
    .B(_07031_),
    .C(_07032_),
    .Y(_07033_));
 NAND2x1_ASAP7_75t_R _25249_ (.A(_14576_),
    .B(_06946_),
    .Y(_07034_));
 OA211x2_ASAP7_75t_R _25250_ (.A1(_16259_),
    .A2(_06946_),
    .B(_07034_),
    .C(_13658_),
    .Y(_07035_));
 NAND2x1_ASAP7_75t_R _25251_ (.A(_06935_),
    .B(net281),
    .Y(_07036_));
 OA33x2_ASAP7_75t_R _25252_ (.A1(_07026_),
    .A2(_07028_),
    .A3(_07030_),
    .B1(_07033_),
    .B2(_07035_),
    .B3(_07036_),
    .Y(_07037_));
 OA211x2_ASAP7_75t_R _25253_ (.A1(_07016_),
    .A2(_07018_),
    .B(_07025_),
    .C(_07037_),
    .Y(_07038_));
 TAPCELL_ASAP7_75t_R TAP_820 ();
 TAPCELL_ASAP7_75t_R TAP_819 ();
 AND2x2_ASAP7_75t_R _25256_ (.A(_14938_),
    .B(_06946_),
    .Y(_07041_));
 AND2x2_ASAP7_75t_R _25257_ (.A(_04829_),
    .B(_06943_),
    .Y(_07042_));
 OA21x2_ASAP7_75t_R _25258_ (.A1(_07041_),
    .A2(_07042_),
    .B(net288),
    .Y(_07043_));
 OR3x1_ASAP7_75t_R _25259_ (.A(_14990_),
    .B(_14992_),
    .C(_06943_),
    .Y(_07044_));
 OA21x2_ASAP7_75t_R _25260_ (.A1(_04718_),
    .A2(_06946_),
    .B(_07044_),
    .Y(_07045_));
 AND2x2_ASAP7_75t_R _25261_ (.A(_13658_),
    .B(_07045_),
    .Y(_07046_));
 NAND2x1_ASAP7_75t_R _25262_ (.A(_14822_),
    .B(_06946_),
    .Y(_07047_));
 OA211x2_ASAP7_75t_R _25263_ (.A1(_05045_),
    .A2(_06946_),
    .B(_07047_),
    .C(net288),
    .Y(_07048_));
 NAND2x1_ASAP7_75t_R _25264_ (.A(_18133_),
    .B(_06946_),
    .Y(_07049_));
 OA211x2_ASAP7_75t_R _25265_ (.A1(_18235_),
    .A2(_06946_),
    .B(_07049_),
    .C(_13658_),
    .Y(_07050_));
 OR3x1_ASAP7_75t_R _25266_ (.A(net281),
    .B(_07048_),
    .C(_07050_),
    .Y(_07051_));
 OA31x2_ASAP7_75t_R _25267_ (.A1(_06939_),
    .A2(_07043_),
    .A3(_07046_),
    .B1(_07051_),
    .Y(_07052_));
 AND3x1_ASAP7_75t_R _25268_ (.A(_06932_),
    .B(_06996_),
    .C(_07052_),
    .Y(_07053_));
 AO21x1_ASAP7_75t_R _25269_ (.A1(_06982_),
    .A2(_07038_),
    .B(_07053_),
    .Y(_07054_));
 AND2x2_ASAP7_75t_R _25270_ (.A(_06932_),
    .B(_06935_),
    .Y(_07055_));
 TAPCELL_ASAP7_75t_R TAP_818 ();
 NAND2x1_ASAP7_75t_R _25272_ (.A(_14688_),
    .B(_06946_),
    .Y(_07057_));
 OA21x2_ASAP7_75t_R _25273_ (.A1(_18253_),
    .A2(_06946_),
    .B(_07057_),
    .Y(_07058_));
 OA222x2_ASAP7_75t_R _25274_ (.A1(_14761_),
    .A2(_07001_),
    .B1(_07002_),
    .B2(_18248_),
    .C1(_07058_),
    .C2(_13658_),
    .Y(_07059_));
 OR2x2_ASAP7_75t_R _25275_ (.A(_05371_),
    .B(_06946_),
    .Y(_07060_));
 OA21x2_ASAP7_75t_R _25276_ (.A1(_13573_),
    .A2(_06943_),
    .B(_07060_),
    .Y(_07061_));
 AO21x1_ASAP7_75t_R _25277_ (.A1(_05478_),
    .A2(_06943_),
    .B(_13658_),
    .Y(_07062_));
 AO21x1_ASAP7_75t_R _25278_ (.A1(_13777_),
    .A2(_06946_),
    .B(_07062_),
    .Y(_07063_));
 OA211x2_ASAP7_75t_R _25279_ (.A1(net290),
    .A2(_07061_),
    .B(_07063_),
    .C(_06939_),
    .Y(_07064_));
 AO21x1_ASAP7_75t_R _25280_ (.A1(_06953_),
    .A2(_07059_),
    .B(_07064_),
    .Y(_07065_));
 XNOR2x2_ASAP7_75t_R _25281_ (.A(_14083_),
    .B(_06927_),
    .Y(_07066_));
 TAPCELL_ASAP7_75t_R TAP_817 ();
 AO21x1_ASAP7_75t_R _25283_ (.A1(_07055_),
    .A2(_07065_),
    .B(_07066_),
    .Y(_07068_));
 OR2x2_ASAP7_75t_R _25284_ (.A(_07054_),
    .B(_07068_),
    .Y(_07069_));
 NAND2x1_ASAP7_75t_R _25285_ (.A(_13364_),
    .B(_13376_),
    .Y(_07070_));
 AND2x6_ASAP7_75t_R _25286_ (.A(_13342_),
    .B(_07070_),
    .Y(_07071_));
 TAPCELL_ASAP7_75t_R TAP_816 ();
 OA211x2_ASAP7_75t_R _25288_ (.A1(_06928_),
    .A2(_07012_),
    .B(_07069_),
    .C(_07071_),
    .Y(_07073_));
 OR3x1_ASAP7_75t_R _25289_ (.A(_13349_),
    .B(_13380_),
    .C(_13385_),
    .Y(_07074_));
 TAPCELL_ASAP7_75t_R TAP_815 ();
 NAND2x2_ASAP7_75t_R _25291_ (.A(_13317_),
    .B(_05743_),
    .Y(_07076_));
 OR3x4_ASAP7_75t_R _25292_ (.A(_05515_),
    .B(_14577_),
    .C(_05518_),
    .Y(_07077_));
 AND2x6_ASAP7_75t_R _25293_ (.A(_07076_),
    .B(_07077_),
    .Y(_07078_));
 NOR3x2_ASAP7_75t_R _25294_ (.B(_14577_),
    .C(_05518_),
    .Y(_07079_),
    .A(_05515_));
 OR2x6_ASAP7_75t_R _25295_ (.A(_05743_),
    .B(_07079_),
    .Y(_07080_));
 TAPCELL_ASAP7_75t_R TAP_814 ();
 AOI22x1_ASAP7_75t_R _25297_ (.A1(_01356_),
    .A2(_07078_),
    .B1(_07080_),
    .B2(_00324_),
    .Y(_07082_));
 AO21x1_ASAP7_75t_R _25298_ (.A1(_13576_),
    .A2(_07082_),
    .B(_06918_),
    .Y(_07083_));
 OR3x1_ASAP7_75t_R _25299_ (.A(_13376_),
    .B(_06574_),
    .C(_06942_),
    .Y(_07084_));
 NAND2x1_ASAP7_75t_R _25300_ (.A(_13386_),
    .B(_13364_),
    .Y(_07085_));
 AO21x2_ASAP7_75t_R _25301_ (.A1(_06576_),
    .A2(_07084_),
    .B(_07085_),
    .Y(_07086_));
 TAPCELL_ASAP7_75t_R TAP_813 ();
 TAPCELL_ASAP7_75t_R TAP_812 ();
 NAND2x1_ASAP7_75t_R _25304_ (.A(_13386_),
    .B(_06574_),
    .Y(_07089_));
 AND3x1_ASAP7_75t_R _25305_ (.A(_02360_),
    .B(_13386_),
    .C(_06574_),
    .Y(_07090_));
 AO21x1_ASAP7_75t_R _25306_ (.A1(_02359_),
    .A2(_07089_),
    .B(_07090_),
    .Y(_07091_));
 NAND2x1_ASAP7_75t_R _25307_ (.A(_07086_),
    .B(_07091_),
    .Y(_07092_));
 AOI21x1_ASAP7_75t_R _25308_ (.A1(_13264_),
    .A2(_13329_),
    .B(_13342_),
    .Y(_07093_));
 OA211x2_ASAP7_75t_R _25309_ (.A1(_13364_),
    .A2(_06574_),
    .B(_07093_),
    .C(_13386_),
    .Y(_07094_));
 TAPCELL_ASAP7_75t_R TAP_811 ();
 OA211x2_ASAP7_75t_R _25311_ (.A1(_00074_),
    .A2(_07086_),
    .B(_07092_),
    .C(_07094_),
    .Y(_07096_));
 AND3x4_ASAP7_75t_R _25312_ (.A(_06573_),
    .B(_06561_),
    .C(_07093_),
    .Y(_07097_));
 TAPCELL_ASAP7_75t_R TAP_810 ();
 AO21x1_ASAP7_75t_R _25314_ (.A1(\ex_block_i.alu_adder_result_ex_o[0] ),
    .A2(_07097_),
    .B(_13567_),
    .Y(_07099_));
 NAND2x2_ASAP7_75t_R _25315_ (.A(_06928_),
    .B(_06932_),
    .Y(_07100_));
 AND4x2_ASAP7_75t_R _25316_ (.A(_13342_),
    .B(_06573_),
    .C(_13376_),
    .D(_05478_),
    .Y(_07101_));
 TAPCELL_ASAP7_75t_R TAP_809 ();
 AND3x1_ASAP7_75t_R _25318_ (.A(_13342_),
    .B(_06573_),
    .C(_13376_),
    .Y(_07103_));
 AND2x2_ASAP7_75t_R _25319_ (.A(net290),
    .B(_06939_),
    .Y(_07104_));
 OA211x2_ASAP7_75t_R _25320_ (.A1(_07103_),
    .A2(_07104_),
    .B(_06935_),
    .C(_06968_),
    .Y(_07105_));
 AO21x2_ASAP7_75t_R _25321_ (.A1(_06996_),
    .A2(_07101_),
    .B(_07105_),
    .Y(_07106_));
 AND2x2_ASAP7_75t_R _25322_ (.A(_06928_),
    .B(_06932_),
    .Y(_07107_));
 TAPCELL_ASAP7_75t_R TAP_808 ();
 OA21x2_ASAP7_75t_R _25324_ (.A1(_07107_),
    .A2(_07101_),
    .B(_06943_),
    .Y(_07109_));
 OA21x2_ASAP7_75t_R _25325_ (.A1(_07100_),
    .A2(_07106_),
    .B(_07109_),
    .Y(_07110_));
 OR4x1_ASAP7_75t_R _25326_ (.A(_07083_),
    .B(_07096_),
    .C(_07099_),
    .D(_07110_),
    .Y(_07111_));
 AO21x1_ASAP7_75t_R _25327_ (.A1(_07074_),
    .A2(_06630_),
    .B(_07111_),
    .Y(_07112_));
 OAI21x1_ASAP7_75t_R _25328_ (.A1(_05558_),
    .A2(_06915_),
    .B(_06919_),
    .Y(_07113_));
 TAPCELL_ASAP7_75t_R TAP_807 ();
 NAND2x2_ASAP7_75t_R _25330_ (.A(_01730_),
    .B(_01731_),
    .Y(_07115_));
 INVx1_ASAP7_75t_R _25331_ (.A(_01863_),
    .Y(_07116_));
 AND2x6_ASAP7_75t_R _25332_ (.A(_01730_),
    .B(_01731_),
    .Y(_07117_));
 AND2x2_ASAP7_75t_R _25333_ (.A(_07116_),
    .B(_07117_),
    .Y(_07118_));
 AO21x1_ASAP7_75t_R _25334_ (.A1(net34),
    .A2(_07115_),
    .B(_07118_),
    .Y(_07119_));
 CKINVDCx8_ASAP7_75t_R _25335_ (.A(net418),
    .Y(_07120_));
 TAPCELL_ASAP7_75t_R TAP_806 ();
 AND2x6_ASAP7_75t_R _25337_ (.A(_07120_),
    .B(net419),
    .Y(_07122_));
 TAPCELL_ASAP7_75t_R TAP_805 ();
 TAPCELL_ASAP7_75t_R TAP_804 ();
 TAPCELL_ASAP7_75t_R TAP_803 ();
 TAPCELL_ASAP7_75t_R TAP_802 ();
 TAPCELL_ASAP7_75t_R TAP_801 ();
 NOR2x2_ASAP7_75t_R _25343_ (.A(net418),
    .B(net419),
    .Y(_07128_));
 AND2x6_ASAP7_75t_R _25344_ (.A(_05738_),
    .B(_01731_),
    .Y(_07129_));
 NOR2x1_ASAP7_75t_R _25345_ (.A(_01855_),
    .B(_07129_),
    .Y(_07130_));
 AO21x1_ASAP7_75t_R _25346_ (.A1(net43),
    .A2(_05738_),
    .B(_07130_),
    .Y(_07131_));
 TAPCELL_ASAP7_75t_R TAP_800 ();
 AND2x2_ASAP7_75t_R _25348_ (.A(net27),
    .B(net420),
    .Y(_07133_));
 NAND2x1_ASAP7_75t_R _25349_ (.A(_01871_),
    .B(_07117_),
    .Y(_07134_));
 INVx13_ASAP7_75t_R _25350_ (.A(net419),
    .Y(_07135_));
 OA211x2_ASAP7_75t_R _25351_ (.A1(net57),
    .A2(_07117_),
    .B(_07134_),
    .C(_07135_),
    .Y(_07136_));
 TAPCELL_ASAP7_75t_R TAP_799 ();
 OA21x2_ASAP7_75t_R _25353_ (.A1(_07133_),
    .A2(_07136_),
    .B(_01642_),
    .Y(_07138_));
 AO221x1_ASAP7_75t_R _25354_ (.A1(_07119_),
    .A2(_07122_),
    .B1(_07128_),
    .B2(_07131_),
    .C(_07138_),
    .Y(_07139_));
 NAND2x2_ASAP7_75t_R _25355_ (.A(_05625_),
    .B(_05629_),
    .Y(_07140_));
 TAPCELL_ASAP7_75t_R TAP_798 ();
 OR4x2_ASAP7_75t_R _25357_ (.A(_13301_),
    .B(_13658_),
    .C(_13954_),
    .D(_05560_),
    .Y(_07142_));
 OA22x2_ASAP7_75t_R _25358_ (.A1(_02139_),
    .A2(_06908_),
    .B1(_07142_),
    .B2(_01913_),
    .Y(_07143_));
 AND4x2_ASAP7_75t_R _25359_ (.A(_13302_),
    .B(_13658_),
    .C(_13955_),
    .D(_05542_),
    .Y(_07144_));
 NAND2x2_ASAP7_75t_R _25360_ (.A(_05679_),
    .B(_07144_),
    .Y(_07145_));
 NAND2x2_ASAP7_75t_R _25361_ (.A(_05630_),
    .B(_07144_),
    .Y(_07146_));
 OA22x2_ASAP7_75t_R _25362_ (.A1(_01995_),
    .A2(_07145_),
    .B1(_07146_),
    .B2(_02029_),
    .Y(_07147_));
 TAPCELL_ASAP7_75t_R TAP_797 ();
 NAND2x2_ASAP7_75t_R _25364_ (.A(_06906_),
    .B(_05630_),
    .Y(_07149_));
 OR4x2_ASAP7_75t_R _25365_ (.A(_13302_),
    .B(net289),
    .C(_13955_),
    .D(_05560_),
    .Y(_07150_));
 OR3x4_ASAP7_75t_R _25366_ (.A(_06911_),
    .B(_06910_),
    .C(_07150_),
    .Y(_07151_));
 TAPCELL_ASAP7_75t_R TAP_796 ();
 OA21x2_ASAP7_75t_R _25368_ (.A1(_01945_),
    .A2(_07149_),
    .B(_07151_),
    .Y(_07153_));
 OA211x2_ASAP7_75t_R _25369_ (.A1(_07140_),
    .A2(_07143_),
    .B(_07147_),
    .C(_07153_),
    .Y(_07154_));
 AND4x2_ASAP7_75t_R _25370_ (.A(_18162_),
    .B(_05609_),
    .C(_05611_),
    .D(_06889_),
    .Y(_07155_));
 TAPCELL_ASAP7_75t_R TAP_795 ();
 NAND2x1_ASAP7_75t_R _25372_ (.A(net62),
    .B(_07155_),
    .Y(_07157_));
 TAPCELL_ASAP7_75t_R TAP_794 ();
 OA31x2_ASAP7_75t_R _25374_ (.A1(_13954_),
    .A2(_14084_),
    .A3(_05581_),
    .B1(_05535_),
    .Y(_07159_));
 TAPCELL_ASAP7_75t_R TAP_793 ();
 TAPCELL_ASAP7_75t_R TAP_792 ();
 OR5x2_ASAP7_75t_R _25377_ (.A(_13301_),
    .B(_13658_),
    .C(_13954_),
    .D(_14084_),
    .E(_05560_),
    .Y(_07162_));
 TAPCELL_ASAP7_75t_R TAP_791 ();
 TAPCELL_ASAP7_75t_R TAP_790 ();
 OAI22x1_ASAP7_75t_R _25380_ (.A1(_02172_),
    .A2(net283),
    .B1(net282),
    .B2(_02066_),
    .Y(_07165_));
 NAND2x1_ASAP7_75t_R _25381_ (.A(_06886_),
    .B(_07165_),
    .Y(_07166_));
 TAPCELL_ASAP7_75t_R TAP_789 ();
 NAND2x2_ASAP7_75t_R _25383_ (.A(_05539_),
    .B(_05582_),
    .Y(_07168_));
 TAPCELL_ASAP7_75t_R TAP_788 ();
 AND4x2_ASAP7_75t_R _25385_ (.A(_13302_),
    .B(net289),
    .C(_13955_),
    .D(_05542_),
    .Y(_07170_));
 NAND2x2_ASAP7_75t_R _25386_ (.A(_05679_),
    .B(_07170_),
    .Y(_07171_));
 NAND2x2_ASAP7_75t_R _25387_ (.A(_05582_),
    .B(_05679_),
    .Y(_07172_));
 OA222x2_ASAP7_75t_R _25388_ (.A1(_00661_),
    .A2(_07168_),
    .B1(_07171_),
    .B2(_02098_),
    .C1(_07172_),
    .C2(_01577_),
    .Y(_07173_));
 OAI22x1_ASAP7_75t_R _25389_ (.A1(_00659_),
    .A2(net284),
    .B1(_07162_),
    .B2(_00660_),
    .Y(_07174_));
 NAND2x1_ASAP7_75t_R _25390_ (.A(_06884_),
    .B(_07174_),
    .Y(_07175_));
 AND5x2_ASAP7_75t_R _25391_ (.A(_07154_),
    .B(_07157_),
    .C(_07166_),
    .D(_07173_),
    .E(_07175_),
    .Y(_07176_));
 NAND2x1_ASAP7_75t_R _25392_ (.A(_13567_),
    .B(_07176_),
    .Y(_07177_));
 OA211x2_ASAP7_75t_R _25393_ (.A1(net294),
    .A2(_07083_),
    .B(_07177_),
    .C(_06920_),
    .Y(_07178_));
 AO21x1_ASAP7_75t_R _25394_ (.A1(_07113_),
    .A2(_07139_),
    .B(_07178_),
    .Y(_07179_));
 OA21x2_ASAP7_75t_R _25395_ (.A1(_07073_),
    .A2(_07112_),
    .B(_07179_),
    .Y(_07180_));
 TAPCELL_ASAP7_75t_R TAP_787 ();
 NOR2x1_ASAP7_75t_R _25397_ (.A(_01709_),
    .B(_06924_),
    .Y(_07182_));
 AO21x1_ASAP7_75t_R _25398_ (.A1(_06924_),
    .A2(_07180_),
    .B(_07182_),
    .Y(_02656_));
 TAPCELL_ASAP7_75t_R TAP_786 ();
 AND2x6_ASAP7_75t_R _25400_ (.A(net418),
    .B(_07135_),
    .Y(_07184_));
 TAPCELL_ASAP7_75t_R TAP_785 ();
 AO221x1_ASAP7_75t_R _25402_ (.A1(net35),
    .A2(_07122_),
    .B1(_07184_),
    .B2(net58),
    .C(_07117_),
    .Y(_07186_));
 INVx1_ASAP7_75t_R _25403_ (.A(_01862_),
    .Y(_07187_));
 INVx1_ASAP7_75t_R _25404_ (.A(_01870_),
    .Y(_07188_));
 AO221x1_ASAP7_75t_R _25405_ (.A1(_07187_),
    .A2(_07122_),
    .B1(_07184_),
    .B2(_07188_),
    .C(_07115_),
    .Y(_07189_));
 INVx1_ASAP7_75t_R _25406_ (.A(net44),
    .Y(_07190_));
 OAI22x1_ASAP7_75t_R _25407_ (.A1(_07190_),
    .A2(_01730_),
    .B1(_01854_),
    .B2(_07129_),
    .Y(_07191_));
 TAPCELL_ASAP7_75t_R TAP_784 ();
 AND2x4_ASAP7_75t_R _25409_ (.A(net418),
    .B(net419),
    .Y(_07193_));
 AO222x2_ASAP7_75t_R _25410_ (.A1(_07186_),
    .A2(_07189_),
    .B1(_07191_),
    .B2(_07128_),
    .C1(net38),
    .C2(_07193_),
    .Y(_07194_));
 TAPCELL_ASAP7_75t_R TAP_783 ();
 NAND2x2_ASAP7_75t_R _25412_ (.A(_00279_),
    .B(_07077_),
    .Y(_07196_));
 TAPCELL_ASAP7_75t_R TAP_782 ();
 TAPCELL_ASAP7_75t_R TAP_781 ();
 AND3x1_ASAP7_75t_R _25415_ (.A(_00279_),
    .B(_01360_),
    .C(_07077_),
    .Y(_07199_));
 AOI21x1_ASAP7_75t_R _25416_ (.A1(_00291_),
    .A2(_07196_),
    .B(_07199_),
    .Y(_07200_));
 NAND2x1_ASAP7_75t_R _25417_ (.A(_00075_),
    .B(_07089_),
    .Y(_07201_));
 AND2x6_ASAP7_75t_R _25418_ (.A(_13386_),
    .B(_06574_),
    .Y(_07202_));
 TAPCELL_ASAP7_75t_R TAP_780 ();
 TAPCELL_ASAP7_75t_R TAP_779 ();
 NAND2x1_ASAP7_75t_R _25421_ (.A(_00076_),
    .B(_07202_),
    .Y(_07205_));
 AOI21x1_ASAP7_75t_R _25422_ (.A1(_06576_),
    .A2(_07084_),
    .B(_07085_),
    .Y(_07206_));
 TAPCELL_ASAP7_75t_R TAP_778 ();
 AO21x1_ASAP7_75t_R _25424_ (.A1(_07201_),
    .A2(_07205_),
    .B(_07206_),
    .Y(_07208_));
 OA211x2_ASAP7_75t_R _25425_ (.A1(_02361_),
    .A2(_07086_),
    .B(_07208_),
    .C(_07094_),
    .Y(_07209_));
 TAPCELL_ASAP7_75t_R TAP_777 ();
 TAPCELL_ASAP7_75t_R TAP_776 ();
 AO21x1_ASAP7_75t_R _25428_ (.A1(net279),
    .A2(_07097_),
    .B(_13576_),
    .Y(_07212_));
 AND2x2_ASAP7_75t_R _25429_ (.A(_06935_),
    .B(_06939_),
    .Y(_07213_));
 AND2x2_ASAP7_75t_R _25430_ (.A(_05478_),
    .B(_07103_),
    .Y(_07214_));
 AND2x2_ASAP7_75t_R _25431_ (.A(_07026_),
    .B(_07214_),
    .Y(_07215_));
 AO21x2_ASAP7_75t_R _25432_ (.A1(_06972_),
    .A2(_07213_),
    .B(_07215_),
    .Y(_07216_));
 OA21x2_ASAP7_75t_R _25433_ (.A1(_07100_),
    .A2(_07216_),
    .B(_07109_),
    .Y(_07217_));
 OR3x1_ASAP7_75t_R _25434_ (.A(_07209_),
    .B(_07212_),
    .C(_07217_),
    .Y(_07218_));
 AND2x2_ASAP7_75t_R _25435_ (.A(_07066_),
    .B(_06932_),
    .Y(_07219_));
 AND3x1_ASAP7_75t_R _25436_ (.A(net288),
    .B(_06983_),
    .C(_06984_),
    .Y(_07220_));
 AO21x1_ASAP7_75t_R _25437_ (.A1(_13658_),
    .A2(_06949_),
    .B(_07220_),
    .Y(_07221_));
 OR2x2_ASAP7_75t_R _25438_ (.A(_15104_),
    .B(_06946_),
    .Y(_07222_));
 AO21x1_ASAP7_75t_R _25439_ (.A1(_06985_),
    .A2(_07222_),
    .B(net288),
    .Y(_07223_));
 OR3x1_ASAP7_75t_R _25440_ (.A(_13658_),
    .B(_06992_),
    .C(_06993_),
    .Y(_07224_));
 AND3x1_ASAP7_75t_R _25441_ (.A(_06939_),
    .B(_07223_),
    .C(_07224_),
    .Y(_07225_));
 AO21x1_ASAP7_75t_R _25442_ (.A1(net281),
    .A2(_07221_),
    .B(_07225_),
    .Y(_07226_));
 AOI211x1_ASAP7_75t_R _25443_ (.A1(_18167_),
    .A2(_06943_),
    .B(_07007_),
    .C(_13658_),
    .Y(_07227_));
 AO21x1_ASAP7_75t_R _25444_ (.A1(_13658_),
    .A2(_06990_),
    .B(_07227_),
    .Y(_07228_));
 NAND2x1_ASAP7_75t_R _25445_ (.A(_15897_),
    .B(_06946_),
    .Y(_07229_));
 OA211x2_ASAP7_75t_R _25446_ (.A1(_18178_),
    .A2(_06946_),
    .B(_07229_),
    .C(net288),
    .Y(_07230_));
 OA211x2_ASAP7_75t_R _25447_ (.A1(_18198_),
    .A2(_06943_),
    .B(_07005_),
    .C(_13658_),
    .Y(_07231_));
 OR3x1_ASAP7_75t_R _25448_ (.A(net281),
    .B(_07230_),
    .C(_07231_),
    .Y(_07232_));
 OA211x2_ASAP7_75t_R _25449_ (.A1(_06939_),
    .A2(_07228_),
    .B(_07232_),
    .C(_06935_),
    .Y(_07233_));
 AO21x2_ASAP7_75t_R _25450_ (.A1(_06996_),
    .A2(_07226_),
    .B(_07233_),
    .Y(_07234_));
 AND2x2_ASAP7_75t_R _25451_ (.A(_07066_),
    .B(_06982_),
    .Y(_07235_));
 OA211x2_ASAP7_75t_R _25452_ (.A1(_18253_),
    .A2(_06943_),
    .B(_06977_),
    .C(net290),
    .Y(_07236_));
 OA211x2_ASAP7_75t_R _25453_ (.A1(_13573_),
    .A2(_06946_),
    .B(_06970_),
    .C(_13658_),
    .Y(_07237_));
 OR2x2_ASAP7_75t_R _25454_ (.A(_07236_),
    .B(_07237_),
    .Y(_07238_));
 OA211x2_ASAP7_75t_R _25455_ (.A1(net290),
    .A2(_07103_),
    .B(_06968_),
    .C(_06953_),
    .Y(_07239_));
 AO21x2_ASAP7_75t_R _25456_ (.A1(_06939_),
    .A2(_07238_),
    .B(_07239_),
    .Y(_07240_));
 OA211x2_ASAP7_75t_R _25457_ (.A1(_05045_),
    .A2(_06943_),
    .B(_06956_),
    .C(net290),
    .Y(_07241_));
 OA211x2_ASAP7_75t_R _25458_ (.A1(_14761_),
    .A2(_06946_),
    .B(_06975_),
    .C(_13658_),
    .Y(_07242_));
 OR3x1_ASAP7_75t_R _25459_ (.A(_06939_),
    .B(_07241_),
    .C(_07242_),
    .Y(_07243_));
 OA21x2_ASAP7_75t_R _25460_ (.A1(_06958_),
    .A2(_06959_),
    .B(net288),
    .Y(_07244_));
 OA211x2_ASAP7_75t_R _25461_ (.A1(_18235_),
    .A2(_06943_),
    .B(_06952_),
    .C(_13658_),
    .Y(_07245_));
 OR3x1_ASAP7_75t_R _25462_ (.A(_06953_),
    .B(_07244_),
    .C(_07245_),
    .Y(_07246_));
 AO21x1_ASAP7_75t_R _25463_ (.A1(_07243_),
    .A2(_07246_),
    .B(_06996_),
    .Y(_07247_));
 OA21x2_ASAP7_75t_R _25464_ (.A1(_06935_),
    .A2(_07240_),
    .B(_07247_),
    .Y(_07248_));
 OA211x2_ASAP7_75t_R _25465_ (.A1(_04603_),
    .A2(_06946_),
    .B(_07027_),
    .C(_13658_),
    .Y(_07249_));
 AO21x1_ASAP7_75t_R _25466_ (.A1(net288),
    .A2(_07045_),
    .B(_07249_),
    .Y(_07250_));
 OA21x2_ASAP7_75t_R _25467_ (.A1(_07041_),
    .A2(_07042_),
    .B(_13658_),
    .Y(_07251_));
 OA211x2_ASAP7_75t_R _25468_ (.A1(_18235_),
    .A2(_06946_),
    .B(_07049_),
    .C(net288),
    .Y(_07252_));
 OR3x1_ASAP7_75t_R _25469_ (.A(net281),
    .B(_07251_),
    .C(_07252_),
    .Y(_07253_));
 OA21x2_ASAP7_75t_R _25470_ (.A1(_06939_),
    .A2(_07250_),
    .B(_07253_),
    .Y(_07254_));
 AND3x2_ASAP7_75t_R _25471_ (.A(_06928_),
    .B(_06932_),
    .C(_06996_),
    .Y(_07255_));
 AND2x2_ASAP7_75t_R _25472_ (.A(_07254_),
    .B(_07255_),
    .Y(_07256_));
 AO221x2_ASAP7_75t_R _25473_ (.A1(_07219_),
    .A2(_07234_),
    .B1(_07235_),
    .B2(_07248_),
    .C(_07256_),
    .Y(_07257_));
 TAPCELL_ASAP7_75t_R TAP_775 ();
 AOI21x1_ASAP7_75t_R _25475_ (.A1(_18167_),
    .A2(_06946_),
    .B(_07020_),
    .Y(_07259_));
 OA211x2_ASAP7_75t_R _25476_ (.A1(_16259_),
    .A2(_06946_),
    .B(_07034_),
    .C(net288),
    .Y(_07260_));
 AO21x1_ASAP7_75t_R _25477_ (.A1(_13658_),
    .A2(_07259_),
    .B(_07260_),
    .Y(_07261_));
 OA21x2_ASAP7_75t_R _25478_ (.A1(_15104_),
    .A2(_06943_),
    .B(net288),
    .Y(_07262_));
 AO32x1_ASAP7_75t_R _25479_ (.A1(_13658_),
    .A2(_07031_),
    .A3(_07032_),
    .B1(_07262_),
    .B2(_07029_),
    .Y(_07263_));
 OR2x2_ASAP7_75t_R _25480_ (.A(net281),
    .B(_07263_),
    .Y(_07264_));
 TAPCELL_ASAP7_75t_R TAP_774 ();
 OA211x2_ASAP7_75t_R _25482_ (.A1(_06939_),
    .A2(_07261_),
    .B(_07264_),
    .C(_06935_),
    .Y(_07266_));
 AO21x1_ASAP7_75t_R _25483_ (.A1(_06998_),
    .A2(_07002_),
    .B(_15668_),
    .Y(_07267_));
 NAND3x1_ASAP7_75t_R _25484_ (.A(_18186_),
    .B(_06998_),
    .C(_07002_),
    .Y(_07268_));
 AO21x1_ASAP7_75t_R _25485_ (.A1(_07267_),
    .A2(_07268_),
    .B(_06939_),
    .Y(_07269_));
 OA211x2_ASAP7_75t_R _25486_ (.A1(_18198_),
    .A2(_06946_),
    .B(_07023_),
    .C(net288),
    .Y(_07270_));
 NAND2x1_ASAP7_75t_R _25487_ (.A(_15897_),
    .B(_06943_),
    .Y(_07271_));
 OA211x2_ASAP7_75t_R _25488_ (.A1(_18178_),
    .A2(_06943_),
    .B(_07271_),
    .C(_13658_),
    .Y(_07272_));
 OR3x1_ASAP7_75t_R _25489_ (.A(net281),
    .B(_07270_),
    .C(_07272_),
    .Y(_07273_));
 AND4x1_ASAP7_75t_R _25490_ (.A(_06982_),
    .B(_06996_),
    .C(_07269_),
    .D(_07273_),
    .Y(_07274_));
 NAND2x1_ASAP7_75t_R _25491_ (.A(_18246_),
    .B(_06943_),
    .Y(_07275_));
 OA211x2_ASAP7_75t_R _25492_ (.A1(_14761_),
    .A2(_06943_),
    .B(_07275_),
    .C(net288),
    .Y(_07276_));
 OA211x2_ASAP7_75t_R _25493_ (.A1(_05045_),
    .A2(_06946_),
    .B(_07047_),
    .C(_13658_),
    .Y(_07277_));
 NOR2x2_ASAP7_75t_R _25494_ (.A(_07276_),
    .B(_07277_),
    .Y(_07278_));
 OA211x2_ASAP7_75t_R _25495_ (.A1(_13573_),
    .A2(_06943_),
    .B(_07060_),
    .C(net290),
    .Y(_07279_));
 AOI211x1_ASAP7_75t_R _25496_ (.A1(_13658_),
    .A2(_07058_),
    .B(_07279_),
    .C(_06953_),
    .Y(_07280_));
 NAND2x1_ASAP7_75t_R _25497_ (.A(_06932_),
    .B(_06935_),
    .Y(_07281_));
 AOI211x1_ASAP7_75t_R _25498_ (.A1(_06953_),
    .A2(_07278_),
    .B(_07280_),
    .C(_07281_),
    .Y(_07282_));
 AOI211x1_ASAP7_75t_R _25499_ (.A1(_06982_),
    .A2(_07266_),
    .B(_07274_),
    .C(_07282_),
    .Y(_07283_));
 NOR2x1_ASAP7_75t_R _25500_ (.A(_07066_),
    .B(_07283_),
    .Y(_07284_));
 OA21x2_ASAP7_75t_R _25501_ (.A1(_07257_),
    .A2(_07284_),
    .B(_07071_),
    .Y(_07285_));
 OA22x2_ASAP7_75t_R _25502_ (.A1(net294),
    .A2(_07200_),
    .B1(_07218_),
    .B2(_07285_),
    .Y(_07286_));
 TAPCELL_ASAP7_75t_R TAP_773 ();
 TAPCELL_ASAP7_75t_R TAP_772 ();
 TAPCELL_ASAP7_75t_R TAP_771 ();
 TAPCELL_ASAP7_75t_R TAP_770 ();
 TAPCELL_ASAP7_75t_R TAP_769 ();
 TAPCELL_ASAP7_75t_R TAP_768 ();
 OAI22x1_ASAP7_75t_R _25509_ (.A1(_01518_),
    .A2(net283),
    .B1(net282),
    .B2(_01487_),
    .Y(_07293_));
 NAND2x1_ASAP7_75t_R _25510_ (.A(_06884_),
    .B(_07293_),
    .Y(_07294_));
 TAPCELL_ASAP7_75t_R TAP_767 ();
 OAI22x1_ASAP7_75t_R _25512_ (.A1(_02171_),
    .A2(net283),
    .B1(net282),
    .B2(_02065_),
    .Y(_07296_));
 NAND2x1_ASAP7_75t_R _25513_ (.A(_06886_),
    .B(_07296_),
    .Y(_07297_));
 TAPCELL_ASAP7_75t_R TAP_766 ();
 NAND2x2_ASAP7_75t_R _25515_ (.A(_05582_),
    .B(_05630_),
    .Y(_07299_));
 TAPCELL_ASAP7_75t_R TAP_765 ();
 OA222x2_ASAP7_75t_R _25517_ (.A1(_02097_),
    .A2(_07171_),
    .B1(_07299_),
    .B2(_02138_),
    .C1(_07172_),
    .C2(_01576_),
    .Y(_07301_));
 OA22x2_ASAP7_75t_R _25518_ (.A1(_01944_),
    .A2(_05588_),
    .B1(_07142_),
    .B2(_01912_),
    .Y(_07302_));
 TAPCELL_ASAP7_75t_R TAP_764 ();
 TAPCELL_ASAP7_75t_R TAP_763 ();
 NAND2x2_ASAP7_75t_R _25521_ (.A(_06906_),
    .B(_05679_),
    .Y(_07305_));
 TAPCELL_ASAP7_75t_R TAP_762 ();
 OA222x2_ASAP7_75t_R _25523_ (.A1(_01994_),
    .A2(_07145_),
    .B1(_07146_),
    .B2(_02028_),
    .C1(_07305_),
    .C2(_00658_),
    .Y(_07307_));
 TAPCELL_ASAP7_75t_R TAP_761 ();
 NAND2x1_ASAP7_75t_R _25525_ (.A(net73),
    .B(_07155_),
    .Y(_07309_));
 OA211x2_ASAP7_75t_R _25526_ (.A1(_07140_),
    .A2(_07302_),
    .B(_07307_),
    .C(_07309_),
    .Y(_07310_));
 AND4x2_ASAP7_75t_R _25527_ (.A(_07294_),
    .B(_07297_),
    .C(_07301_),
    .D(_07310_),
    .Y(_07311_));
 NAND2x1_ASAP7_75t_R _25528_ (.A(_06920_),
    .B(_07311_),
    .Y(_07312_));
 OA22x2_ASAP7_75t_R _25529_ (.A1(_06920_),
    .A2(_07194_),
    .B1(_07286_),
    .B2(_07312_),
    .Y(_07313_));
 NOR2x1_ASAP7_75t_R _25530_ (.A(_01708_),
    .B(_06924_),
    .Y(_07314_));
 AO21x1_ASAP7_75t_R _25531_ (.A1(_06924_),
    .A2(_07313_),
    .B(_07314_),
    .Y(_02657_));
 OA21x2_ASAP7_75t_R _25532_ (.A1(_13658_),
    .A2(_06990_),
    .B(_06994_),
    .Y(_07315_));
 OA21x2_ASAP7_75t_R _25533_ (.A1(_07006_),
    .A2(_07008_),
    .B(_06939_),
    .Y(_07316_));
 AO21x1_ASAP7_75t_R _25534_ (.A1(net281),
    .A2(_07315_),
    .B(_07316_),
    .Y(_07317_));
 AND2x2_ASAP7_75t_R _25535_ (.A(_06939_),
    .B(_06987_),
    .Y(_07318_));
 OR3x1_ASAP7_75t_R _25536_ (.A(net288),
    .B(_06958_),
    .C(_06959_),
    .Y(_07319_));
 OA211x2_ASAP7_75t_R _25537_ (.A1(_13658_),
    .A2(_06949_),
    .B(_07319_),
    .C(net281),
    .Y(_07320_));
 OR3x1_ASAP7_75t_R _25538_ (.A(_06935_),
    .B(_07318_),
    .C(_07320_),
    .Y(_07321_));
 OA21x2_ASAP7_75t_R _25539_ (.A1(_06996_),
    .A2(_07317_),
    .B(_07321_),
    .Y(_07322_));
 OR3x1_ASAP7_75t_R _25540_ (.A(_06939_),
    .B(_06976_),
    .C(_06978_),
    .Y(_07323_));
 OA211x2_ASAP7_75t_R _25541_ (.A1(_18235_),
    .A2(_06943_),
    .B(_06952_),
    .C(net290),
    .Y(_07324_));
 OA211x2_ASAP7_75t_R _25542_ (.A1(_05045_),
    .A2(_06943_),
    .B(_06956_),
    .C(_13658_),
    .Y(_07325_));
 OR3x1_ASAP7_75t_R _25543_ (.A(_06953_),
    .B(_07324_),
    .C(_07325_),
    .Y(_07326_));
 AND3x2_ASAP7_75t_R _25544_ (.A(_06935_),
    .B(_07323_),
    .C(_07326_),
    .Y(_07327_));
 OR2x2_ASAP7_75t_R _25545_ (.A(_06939_),
    .B(_07101_),
    .Y(_07328_));
 OA211x2_ASAP7_75t_R _25546_ (.A1(_06953_),
    .A2(_06972_),
    .B(_07328_),
    .C(_06996_),
    .Y(_07329_));
 OA21x2_ASAP7_75t_R _25547_ (.A1(_07327_),
    .A2(_07329_),
    .B(_06982_),
    .Y(_07330_));
 AO21x1_ASAP7_75t_R _25548_ (.A1(_06932_),
    .A2(_07322_),
    .B(_07330_),
    .Y(_07331_));
 OR2x2_ASAP7_75t_R _25549_ (.A(_07021_),
    .B(_07024_),
    .Y(_07332_));
 OR3x1_ASAP7_75t_R _25550_ (.A(net281),
    .B(_07033_),
    .C(_07035_),
    .Y(_07333_));
 OA21x2_ASAP7_75t_R _25551_ (.A1(_06939_),
    .A2(_07332_),
    .B(_07333_),
    .Y(_07334_));
 AO21x1_ASAP7_75t_R _25552_ (.A1(_06999_),
    .A2(_07003_),
    .B(_06939_),
    .Y(_07335_));
 OA211x2_ASAP7_75t_R _25553_ (.A1(net281),
    .A2(_07018_),
    .B(_07335_),
    .C(_06996_),
    .Y(_07336_));
 AO21x1_ASAP7_75t_R _25554_ (.A1(_06935_),
    .A2(_07334_),
    .B(_07336_),
    .Y(_07337_));
 AND2x6_ASAP7_75t_R _25555_ (.A(_06928_),
    .B(_06982_),
    .Y(_07338_));
 OR3x1_ASAP7_75t_R _25556_ (.A(net281),
    .B(_07043_),
    .C(_07046_),
    .Y(_07339_));
 OA31x2_ASAP7_75t_R _25557_ (.A1(_06939_),
    .A2(_07028_),
    .A3(_07030_),
    .B1(_07339_),
    .Y(_07340_));
 AND2x2_ASAP7_75t_R _25558_ (.A(_06928_),
    .B(_07055_),
    .Y(_07341_));
 OR3x1_ASAP7_75t_R _25559_ (.A(_06939_),
    .B(_07048_),
    .C(_07050_),
    .Y(_07342_));
 OA211x2_ASAP7_75t_R _25560_ (.A1(net281),
    .A2(_07059_),
    .B(_07341_),
    .C(_07342_),
    .Y(_07343_));
 AO21x1_ASAP7_75t_R _25561_ (.A1(_07255_),
    .A2(_07340_),
    .B(_07343_),
    .Y(_07344_));
 AO221x1_ASAP7_75t_R _25562_ (.A1(_07066_),
    .A2(_07331_),
    .B1(_07337_),
    .B2(_07338_),
    .C(_07344_),
    .Y(_07345_));
 AO21x1_ASAP7_75t_R _25563_ (.A1(_06932_),
    .A2(_06935_),
    .B(_07101_),
    .Y(_07346_));
 OA21x2_ASAP7_75t_R _25564_ (.A1(_07281_),
    .A2(_07240_),
    .B(_07346_),
    .Y(_07347_));
 AND2x4_ASAP7_75t_R _25565_ (.A(_06928_),
    .B(_06943_),
    .Y(_07348_));
 TAPCELL_ASAP7_75t_R TAP_760 ();
 TAPCELL_ASAP7_75t_R TAP_759 ();
 INVx1_ASAP7_75t_R _25568_ (.A(_00077_),
    .Y(_07351_));
 TAPCELL_ASAP7_75t_R TAP_758 ();
 TAPCELL_ASAP7_75t_R TAP_757 ();
 NAND2x1_ASAP7_75t_R _25571_ (.A(_00078_),
    .B(_07202_),
    .Y(_07354_));
 OA211x2_ASAP7_75t_R _25572_ (.A1(_07351_),
    .A2(_07202_),
    .B(_07354_),
    .C(_07086_),
    .Y(_07355_));
 AO21x1_ASAP7_75t_R _25573_ (.A1(_02362_),
    .A2(_07206_),
    .B(_07355_),
    .Y(_07356_));
 TAPCELL_ASAP7_75t_R TAP_756 ();
 TAPCELL_ASAP7_75t_R TAP_755 ();
 AO222x2_ASAP7_75t_R _25576_ (.A1(net171),
    .A2(_07097_),
    .B1(_07347_),
    .B2(_07348_),
    .C1(_07356_),
    .C2(_07094_),
    .Y(_07359_));
 TAPCELL_ASAP7_75t_R TAP_754 ();
 TAPCELL_ASAP7_75t_R TAP_753 ();
 TAPCELL_ASAP7_75t_R TAP_752 ();
 OAI22x1_ASAP7_75t_R _25580_ (.A1(_01517_),
    .A2(net283),
    .B1(net282),
    .B2(_01486_),
    .Y(_07363_));
 NAND2x1_ASAP7_75t_R _25581_ (.A(_06884_),
    .B(_07363_),
    .Y(_07364_));
 TAPCELL_ASAP7_75t_R TAP_751 ();
 OAI22x1_ASAP7_75t_R _25583_ (.A1(_02137_),
    .A2(_06908_),
    .B1(_07142_),
    .B2(_01911_),
    .Y(_07366_));
 NAND2x1_ASAP7_75t_R _25584_ (.A(_05627_),
    .B(_07366_),
    .Y(_07367_));
 AO221x2_ASAP7_75t_R _25585_ (.A1(_01364_),
    .A2(_07078_),
    .B1(_07080_),
    .B2(_00663_),
    .C(_13318_),
    .Y(_07368_));
 INVx1_ASAP7_75t_R _25586_ (.A(_01993_),
    .Y(_07369_));
 INVx1_ASAP7_75t_R _25587_ (.A(_02027_),
    .Y(_07370_));
 AO22x1_ASAP7_75t_R _25588_ (.A1(_07369_),
    .A2(_05679_),
    .B1(_05627_),
    .B2(_07370_),
    .Y(_07371_));
 NAND2x1_ASAP7_75t_R _25589_ (.A(_07144_),
    .B(_07371_),
    .Y(_07372_));
 AND4x1_ASAP7_75t_R _25590_ (.A(_07364_),
    .B(_07367_),
    .C(_07368_),
    .D(_07372_),
    .Y(_07373_));
 OAI22x1_ASAP7_75t_R _25591_ (.A1(_02170_),
    .A2(net283),
    .B1(net282),
    .B2(_02064_),
    .Y(_07374_));
 INVx1_ASAP7_75t_R _25592_ (.A(_02096_),
    .Y(_07375_));
 INVx1_ASAP7_75t_R _25593_ (.A(_01575_),
    .Y(_07376_));
 INVx1_ASAP7_75t_R _25594_ (.A(_01943_),
    .Y(_07377_));
 AO221x1_ASAP7_75t_R _25595_ (.A1(_07376_),
    .A2(_05679_),
    .B1(_05630_),
    .B2(_07377_),
    .C(_05632_),
    .Y(_07378_));
 AO32x1_ASAP7_75t_R _25596_ (.A1(_07375_),
    .A2(_05679_),
    .A3(_07170_),
    .B1(_07378_),
    .B2(_06906_),
    .Y(_07379_));
 INVx1_ASAP7_75t_R _25597_ (.A(_01315_),
    .Y(_07380_));
 AO33x2_ASAP7_75t_R _25598_ (.A1(_07380_),
    .A2(_05538_),
    .A3(_05584_),
    .B1(_05679_),
    .B2(_05582_),
    .B3(_06870_),
    .Y(_07381_));
 OR2x2_ASAP7_75t_R _25599_ (.A(_07379_),
    .B(_07381_),
    .Y(_07382_));
 AOI221x1_ASAP7_75t_R _25600_ (.A1(net84),
    .A2(_07155_),
    .B1(_06886_),
    .B2(_07374_),
    .C(_07382_),
    .Y(_07383_));
 NAND2x1_ASAP7_75t_R _25601_ (.A(_07373_),
    .B(_07383_),
    .Y(_07384_));
 AO221x1_ASAP7_75t_R _25602_ (.A1(_07071_),
    .A2(_07345_),
    .B1(_07359_),
    .B2(net294),
    .C(_07384_),
    .Y(_07385_));
 TAPCELL_ASAP7_75t_R TAP_750 ();
 TAPCELL_ASAP7_75t_R TAP_749 ();
 NAND2x2_ASAP7_75t_R _25605_ (.A(_07120_),
    .B(net420),
    .Y(_07388_));
 TAPCELL_ASAP7_75t_R TAP_748 ();
 NAND2x1_ASAP7_75t_R _25607_ (.A(net418),
    .B(_07135_),
    .Y(_07390_));
 OAI22x1_ASAP7_75t_R _25608_ (.A1(_01861_),
    .A2(_07388_),
    .B1(_07390_),
    .B2(_01869_),
    .Y(_07391_));
 AO221x1_ASAP7_75t_R _25609_ (.A1(net36),
    .A2(_07122_),
    .B1(_07184_),
    .B2(net28),
    .C(_07117_),
    .Y(_07392_));
 OA21x2_ASAP7_75t_R _25610_ (.A1(_07115_),
    .A2(_07391_),
    .B(_07392_),
    .Y(_07393_));
 NOR2x1_ASAP7_75t_R _25611_ (.A(_01853_),
    .B(_07129_),
    .Y(_07394_));
 AO21x1_ASAP7_75t_R _25612_ (.A1(net45),
    .A2(_05738_),
    .B(_07394_),
    .Y(_07395_));
 AO22x1_ASAP7_75t_R _25613_ (.A1(net49),
    .A2(_07193_),
    .B1(_07395_),
    .B2(_07128_),
    .Y(_07396_));
 OR3x1_ASAP7_75t_R _25614_ (.A(_06920_),
    .B(_07393_),
    .C(_07396_),
    .Y(_07397_));
 OA21x2_ASAP7_75t_R _25615_ (.A1(_07113_),
    .A2(_07385_),
    .B(_07397_),
    .Y(_07398_));
 NOR2x1_ASAP7_75t_R _25616_ (.A(_01707_),
    .B(_06924_),
    .Y(_07399_));
 AO21x1_ASAP7_75t_R _25617_ (.A1(_06924_),
    .A2(_07398_),
    .B(_07399_),
    .Y(_02658_));
 OA21x2_ASAP7_75t_R _25618_ (.A1(_07244_),
    .A2(_07245_),
    .B(_06953_),
    .Y(_07400_));
 AO21x2_ASAP7_75t_R _25619_ (.A1(_06939_),
    .A2(_07221_),
    .B(_07400_),
    .Y(_07401_));
 AO21x1_ASAP7_75t_R _25620_ (.A1(_07223_),
    .A2(_07224_),
    .B(_06939_),
    .Y(_07402_));
 OA211x2_ASAP7_75t_R _25621_ (.A1(net281),
    .A2(_07228_),
    .B(_07402_),
    .C(_06935_),
    .Y(_07403_));
 AOI21x1_ASAP7_75t_R _25622_ (.A1(_06996_),
    .A2(_07401_),
    .B(_07403_),
    .Y(_07404_));
 OR2x2_ASAP7_75t_R _25623_ (.A(_07241_),
    .B(_07242_),
    .Y(_07405_));
 AND2x2_ASAP7_75t_R _25624_ (.A(_06935_),
    .B(_06953_),
    .Y(_07406_));
 OA211x2_ASAP7_75t_R _25625_ (.A1(_07103_),
    .A2(_07104_),
    .B(_06996_),
    .C(_06968_),
    .Y(_07407_));
 AO221x2_ASAP7_75t_R _25626_ (.A1(_07213_),
    .A2(_07405_),
    .B1(_07238_),
    .B2(_07406_),
    .C(_07407_),
    .Y(_07408_));
 NOR2x1_ASAP7_75t_R _25627_ (.A(_06932_),
    .B(_07408_),
    .Y(_07409_));
 AO21x2_ASAP7_75t_R _25628_ (.A1(_06932_),
    .A2(_07404_),
    .B(_07409_),
    .Y(_07410_));
 OR3x1_ASAP7_75t_R _25629_ (.A(_06939_),
    .B(_07270_),
    .C(_07272_),
    .Y(_07411_));
 OA21x2_ASAP7_75t_R _25630_ (.A1(net281),
    .A2(_07261_),
    .B(_07411_),
    .Y(_07412_));
 AO21x1_ASAP7_75t_R _25631_ (.A1(_07267_),
    .A2(_07268_),
    .B(net281),
    .Y(_07413_));
 OR3x1_ASAP7_75t_R _25632_ (.A(_06939_),
    .B(_07230_),
    .C(_07231_),
    .Y(_07414_));
 AND3x1_ASAP7_75t_R _25633_ (.A(_06996_),
    .B(_07413_),
    .C(_07414_),
    .Y(_07415_));
 AO21x1_ASAP7_75t_R _25634_ (.A1(_06935_),
    .A2(_07412_),
    .B(_07415_),
    .Y(_07416_));
 NAND2x1_ASAP7_75t_R _25635_ (.A(_06939_),
    .B(_07278_),
    .Y(_07417_));
 OR3x1_ASAP7_75t_R _25636_ (.A(_06939_),
    .B(_07251_),
    .C(_07252_),
    .Y(_07418_));
 AND2x2_ASAP7_75t_R _25637_ (.A(net281),
    .B(_07263_),
    .Y(_07419_));
 AO21x1_ASAP7_75t_R _25638_ (.A1(_06939_),
    .A2(_07250_),
    .B(_07419_),
    .Y(_07420_));
 AO32x1_ASAP7_75t_R _25639_ (.A1(_07341_),
    .A2(_07417_),
    .A3(_07418_),
    .B1(_07420_),
    .B2(_07255_),
    .Y(_07421_));
 AOI21x1_ASAP7_75t_R _25640_ (.A1(_07338_),
    .A2(_07416_),
    .B(_07421_),
    .Y(_07422_));
 OAI21x1_ASAP7_75t_R _25641_ (.A1(_06928_),
    .A2(_07410_),
    .B(_07422_),
    .Y(_07423_));
 INVx1_ASAP7_75t_R _25642_ (.A(_00079_),
    .Y(_07424_));
 NAND2x1_ASAP7_75t_R _25643_ (.A(_00080_),
    .B(_07202_),
    .Y(_07425_));
 TAPCELL_ASAP7_75t_R TAP_747 ();
 OA211x2_ASAP7_75t_R _25645_ (.A1(_07424_),
    .A2(_07202_),
    .B(_07425_),
    .C(_07086_),
    .Y(_07427_));
 AO21x1_ASAP7_75t_R _25646_ (.A1(_02363_),
    .A2(_07206_),
    .B(_07427_),
    .Y(_07428_));
 AO22x1_ASAP7_75t_R _25647_ (.A1(net275),
    .A2(_07097_),
    .B1(_07428_),
    .B2(_07094_),
    .Y(_07429_));
 NAND2x2_ASAP7_75t_R _25648_ (.A(_06928_),
    .B(_06943_),
    .Y(_07430_));
 NOR2x1_ASAP7_75t_R _25649_ (.A(_07055_),
    .B(_07101_),
    .Y(_07431_));
 AO21x2_ASAP7_75t_R _25650_ (.A1(_06980_),
    .A2(_07055_),
    .B(_07431_),
    .Y(_07432_));
 NOR2x1_ASAP7_75t_R _25651_ (.A(_07430_),
    .B(_07432_),
    .Y(_07433_));
 OA21x2_ASAP7_75t_R _25652_ (.A1(_07429_),
    .A2(_07433_),
    .B(net294),
    .Y(_07434_));
 NAND2x1_ASAP7_75t_R _25653_ (.A(_00665_),
    .B(_07080_),
    .Y(_07435_));
 TAPCELL_ASAP7_75t_R TAP_746 ();
 NAND2x1_ASAP7_75t_R _25655_ (.A(_07076_),
    .B(_07077_),
    .Y(_07437_));
 OA21x2_ASAP7_75t_R _25656_ (.A1(_02231_),
    .A2(_07437_),
    .B(_13576_),
    .Y(_07438_));
 TAPCELL_ASAP7_75t_R TAP_745 ();
 TAPCELL_ASAP7_75t_R TAP_744 ();
 TAPCELL_ASAP7_75t_R TAP_743 ();
 OAI22x1_ASAP7_75t_R _25660_ (.A1(_02169_),
    .A2(net283),
    .B1(net282),
    .B2(_02063_),
    .Y(_07442_));
 AND2x2_ASAP7_75t_R _25661_ (.A(_06886_),
    .B(_07442_),
    .Y(_07443_));
 INVx1_ASAP7_75t_R _25662_ (.A(_02136_),
    .Y(_07444_));
 TAPCELL_ASAP7_75t_R TAP_742 ();
 AO22x1_ASAP7_75t_R _25664_ (.A1(_07444_),
    .A2(_05582_),
    .B1(_06889_),
    .B2(net146),
    .Y(_07446_));
 AND2x2_ASAP7_75t_R _25665_ (.A(_05611_),
    .B(_05678_),
    .Y(_07447_));
 NAND3x2_ASAP7_75t_R _25666_ (.B(_05572_),
    .C(_07447_),
    .Y(_07448_),
    .A(_14497_));
 OAI22x1_ASAP7_75t_R _25667_ (.A1(_01992_),
    .A2(_07448_),
    .B1(_07140_),
    .B2(_02026_),
    .Y(_07449_));
 OA211x2_ASAP7_75t_R _25668_ (.A1(_05558_),
    .A2(_05586_),
    .B(_05576_),
    .C(_06190_),
    .Y(_07450_));
 OA21x2_ASAP7_75t_R _25669_ (.A1(_05539_),
    .A2(_07450_),
    .B(_05582_),
    .Y(_07451_));
 AO221x1_ASAP7_75t_R _25670_ (.A1(net87),
    .A2(_07155_),
    .B1(_07144_),
    .B2(_07449_),
    .C(_07451_),
    .Y(_07452_));
 AO21x1_ASAP7_75t_R _25671_ (.A1(_05630_),
    .A2(_07446_),
    .B(_07452_),
    .Y(_07453_));
 OAI22x1_ASAP7_75t_R _25672_ (.A1(_01516_),
    .A2(net283),
    .B1(net282),
    .B2(_01485_),
    .Y(_07454_));
 OAI22x1_ASAP7_75t_R _25673_ (.A1(_00081_),
    .A2(_07448_),
    .B1(_07140_),
    .B2(_01942_),
    .Y(_07455_));
 OAI22x1_ASAP7_75t_R _25674_ (.A1(_02095_),
    .A2(_07448_),
    .B1(_07140_),
    .B2(_01910_),
    .Y(_07456_));
 AO32x1_ASAP7_75t_R _25675_ (.A1(_06211_),
    .A2(_05632_),
    .A3(_06889_),
    .B1(_07170_),
    .B2(_07456_),
    .Y(_07457_));
 AO221x1_ASAP7_75t_R _25676_ (.A1(_06884_),
    .A2(_07454_),
    .B1(_07455_),
    .B2(_06906_),
    .C(_07457_),
    .Y(_07458_));
 OR3x4_ASAP7_75t_R _25677_ (.A(_07443_),
    .B(_07453_),
    .C(_07458_),
    .Y(_07459_));
 AO21x2_ASAP7_75t_R _25678_ (.A1(_07435_),
    .A2(_07438_),
    .B(_07459_),
    .Y(_07460_));
 AO211x2_ASAP7_75t_R _25679_ (.A1(_07071_),
    .A2(_07423_),
    .B(_07434_),
    .C(_07460_),
    .Y(_07461_));
 OAI22x1_ASAP7_75t_R _25680_ (.A1(_01860_),
    .A2(_07388_),
    .B1(_07390_),
    .B2(_01868_),
    .Y(_07462_));
 AO221x1_ASAP7_75t_R _25681_ (.A1(net37),
    .A2(_07122_),
    .B1(_07184_),
    .B2(net29),
    .C(_07117_),
    .Y(_07463_));
 OA21x2_ASAP7_75t_R _25682_ (.A1(_07115_),
    .A2(_07462_),
    .B(_07463_),
    .Y(_07464_));
 NOR2x1_ASAP7_75t_R _25683_ (.A(_01852_),
    .B(_07129_),
    .Y(_07465_));
 AO21x1_ASAP7_75t_R _25684_ (.A1(net46),
    .A2(_05738_),
    .B(_07465_),
    .Y(_07466_));
 AO22x1_ASAP7_75t_R _25685_ (.A1(net52),
    .A2(_07193_),
    .B1(_07466_),
    .B2(_07128_),
    .Y(_07467_));
 OR3x1_ASAP7_75t_R _25686_ (.A(_06920_),
    .B(_07464_),
    .C(_07467_),
    .Y(_07468_));
 OA21x2_ASAP7_75t_R _25687_ (.A1(_07113_),
    .A2(_07461_),
    .B(_07468_),
    .Y(_07469_));
 NOR2x1_ASAP7_75t_R _25688_ (.A(_01706_),
    .B(_06924_),
    .Y(_07470_));
 AO21x1_ASAP7_75t_R _25689_ (.A1(_06924_),
    .A2(_07469_),
    .B(_07470_),
    .Y(_02659_));
 TAPCELL_ASAP7_75t_R TAP_741 ();
 AO221x1_ASAP7_75t_R _25691_ (.A1(net39),
    .A2(_07122_),
    .B1(_07184_),
    .B2(net30),
    .C(_07117_),
    .Y(_07472_));
 INVx1_ASAP7_75t_R _25692_ (.A(_01859_),
    .Y(_07473_));
 INVx1_ASAP7_75t_R _25693_ (.A(_01867_),
    .Y(_07474_));
 AO221x1_ASAP7_75t_R _25694_ (.A1(_07473_),
    .A2(_07122_),
    .B1(_07184_),
    .B2(_07474_),
    .C(_07115_),
    .Y(_07475_));
 NOR2x1_ASAP7_75t_R _25695_ (.A(_01851_),
    .B(_07129_),
    .Y(_07476_));
 AO21x1_ASAP7_75t_R _25696_ (.A1(net47),
    .A2(_05738_),
    .B(_07476_),
    .Y(_07477_));
 AO222x2_ASAP7_75t_R _25697_ (.A1(net53),
    .A2(_07193_),
    .B1(_07472_),
    .B2(_07475_),
    .C1(_07477_),
    .C2(_07128_),
    .Y(_07478_));
 OR3x1_ASAP7_75t_R _25698_ (.A(_06996_),
    .B(_06988_),
    .C(_06995_),
    .Y(_07479_));
 AO211x2_ASAP7_75t_R _25699_ (.A1(net290),
    .A2(_06955_),
    .B(_06962_),
    .C(_06935_),
    .Y(_07480_));
 AO21x1_ASAP7_75t_R _25700_ (.A1(_07479_),
    .A2(_07480_),
    .B(_06982_),
    .Y(_07481_));
 OA211x2_ASAP7_75t_R _25701_ (.A1(_06939_),
    .A2(_06972_),
    .B(_06979_),
    .C(_06935_),
    .Y(_07482_));
 AO21x1_ASAP7_75t_R _25702_ (.A1(_06996_),
    .A2(_07101_),
    .B(_06932_),
    .Y(_07483_));
 OA21x2_ASAP7_75t_R _25703_ (.A1(_07482_),
    .A2(_07483_),
    .B(_07066_),
    .Y(_07484_));
 OR3x1_ASAP7_75t_R _25704_ (.A(net281),
    .B(_07021_),
    .C(_07024_),
    .Y(_07485_));
 OA211x2_ASAP7_75t_R _25705_ (.A1(_06939_),
    .A2(_07018_),
    .B(_07485_),
    .C(_06935_),
    .Y(_07486_));
 AND3x1_ASAP7_75t_R _25706_ (.A(_06996_),
    .B(_07004_),
    .C(_07009_),
    .Y(_07487_));
 OA21x2_ASAP7_75t_R _25707_ (.A1(_07486_),
    .A2(_07487_),
    .B(_07338_),
    .Y(_07488_));
 OR3x1_ASAP7_75t_R _25708_ (.A(net281),
    .B(_07028_),
    .C(_07030_),
    .Y(_07489_));
 OR3x1_ASAP7_75t_R _25709_ (.A(_06939_),
    .B(_07033_),
    .C(_07035_),
    .Y(_07490_));
 AO32x1_ASAP7_75t_R _25710_ (.A1(_07489_),
    .A2(_07490_),
    .A3(_07255_),
    .B1(_07341_),
    .B2(_07052_),
    .Y(_07491_));
 AO211x2_ASAP7_75t_R _25711_ (.A1(_07481_),
    .A2(_07484_),
    .B(_07488_),
    .C(_07491_),
    .Y(_07492_));
 OAI21x1_ASAP7_75t_R _25712_ (.A1(_07100_),
    .A2(_07408_),
    .B(_07109_),
    .Y(_07493_));
 INVx1_ASAP7_75t_R _25713_ (.A(_00082_),
    .Y(_07494_));
 TAPCELL_ASAP7_75t_R TAP_740 ();
 NAND2x1_ASAP7_75t_R _25715_ (.A(_00083_),
    .B(_07202_),
    .Y(_07496_));
 OA211x2_ASAP7_75t_R _25716_ (.A1(_07494_),
    .A2(_07202_),
    .B(_07496_),
    .C(_07086_),
    .Y(_07497_));
 AO21x1_ASAP7_75t_R _25717_ (.A1(_02364_),
    .A2(_07206_),
    .B(_07497_),
    .Y(_07498_));
 AOI22x1_ASAP7_75t_R _25718_ (.A1(net175),
    .A2(_07097_),
    .B1(_07498_),
    .B2(_07094_),
    .Y(_07499_));
 AO221x2_ASAP7_75t_R _25719_ (.A1(_01376_),
    .A2(_07078_),
    .B1(_07080_),
    .B2(_00668_),
    .C(_13318_),
    .Y(_07500_));
 OA21x2_ASAP7_75t_R _25720_ (.A1(_13576_),
    .A2(_07499_),
    .B(_07500_),
    .Y(_07501_));
 OAI22x1_ASAP7_75t_R _25721_ (.A1(_01515_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01484_),
    .Y(_07502_));
 NAND2x1_ASAP7_75t_R _25722_ (.A(_06884_),
    .B(_07502_),
    .Y(_07503_));
 AND4x2_ASAP7_75t_R _25723_ (.A(_13302_),
    .B(net289),
    .C(_13955_),
    .D(_05542_),
    .Y(_07504_));
 NAND2x2_ASAP7_75t_R _25724_ (.A(_06892_),
    .B(_07504_),
    .Y(_07505_));
 TAPCELL_ASAP7_75t_R TAP_739 ();
 NAND3x2_ASAP7_75t_R _25726_ (.B(_05625_),
    .C(_05626_),
    .Y(_07507_),
    .A(_05537_));
 OR2x6_ASAP7_75t_R _25727_ (.A(_06908_),
    .B(_07507_),
    .Y(_07508_));
 TAPCELL_ASAP7_75t_R TAP_738 ();
 OA22x2_ASAP7_75t_R _25729_ (.A1(_02094_),
    .A2(_07505_),
    .B1(_07508_),
    .B2(_02135_),
    .Y(_07510_));
 NAND3x2_ASAP7_75t_R _25730_ (.B(_05658_),
    .C(_06892_),
    .Y(_07511_),
    .A(_05541_));
 TAPCELL_ASAP7_75t_R TAP_737 ();
 OR4x2_ASAP7_75t_R _25732_ (.A(_13302_),
    .B(net289),
    .C(_13954_),
    .D(_05560_),
    .Y(_07513_));
 TAPCELL_ASAP7_75t_R TAP_736 ();
 INVx2_ASAP7_75t_R _25734_ (.A(_07513_),
    .Y(_07515_));
 NAND2x2_ASAP7_75t_R _25735_ (.A(_06892_),
    .B(_07515_),
    .Y(_07516_));
 TAPCELL_ASAP7_75t_R TAP_735 ();
 OA22x2_ASAP7_75t_R _25737_ (.A1(_01991_),
    .A2(_07511_),
    .B1(_07516_),
    .B2(_00084_),
    .Y(_07518_));
 OAI22x1_ASAP7_75t_R _25738_ (.A1(_02168_),
    .A2(net284),
    .B1(_07162_),
    .B2(_02062_),
    .Y(_07519_));
 OR4x2_ASAP7_75t_R _25739_ (.A(_13301_),
    .B(_13658_),
    .C(_13954_),
    .D(_05560_),
    .Y(_07520_));
 OAI22x1_ASAP7_75t_R _25740_ (.A1(_01941_),
    .A2(_07513_),
    .B1(_07520_),
    .B2(_01909_),
    .Y(_07521_));
 INVx1_ASAP7_75t_R _25741_ (.A(_07507_),
    .Y(_07522_));
 OR4x2_ASAP7_75t_R _25742_ (.A(_13301_),
    .B(net289),
    .C(_13954_),
    .D(_05560_),
    .Y(_07523_));
 OR2x6_ASAP7_75t_R _25743_ (.A(_07507_),
    .B(_07523_),
    .Y(_07524_));
 TAPCELL_ASAP7_75t_R TAP_734 ();
 OAI21x1_ASAP7_75t_R _25745_ (.A1(_02025_),
    .A2(_07524_),
    .B(_07168_),
    .Y(_07526_));
 AOI221x1_ASAP7_75t_R _25746_ (.A1(_06886_),
    .A2(_07519_),
    .B1(_07521_),
    .B2(_07522_),
    .C(_07526_),
    .Y(_07527_));
 TAPCELL_ASAP7_75t_R TAP_733 ();
 NAND2x2_ASAP7_75t_R _25748_ (.A(net88),
    .B(_06891_),
    .Y(_07529_));
 AND5x2_ASAP7_75t_R _25749_ (.A(_07503_),
    .B(_07510_),
    .C(_07518_),
    .D(_07527_),
    .E(_07529_),
    .Y(_07530_));
 AND3x1_ASAP7_75t_R _25750_ (.A(_07493_),
    .B(_07501_),
    .C(_07530_),
    .Y(_07531_));
 NAND2x1_ASAP7_75t_R _25751_ (.A(_06920_),
    .B(_07531_),
    .Y(_07532_));
 AO21x1_ASAP7_75t_R _25752_ (.A1(_07071_),
    .A2(_07492_),
    .B(_07532_),
    .Y(_07533_));
 OA21x2_ASAP7_75t_R _25753_ (.A1(_06920_),
    .A2(_07478_),
    .B(_07533_),
    .Y(_07534_));
 NOR2x1_ASAP7_75t_R _25754_ (.A(_01705_),
    .B(_06924_),
    .Y(_07535_));
 AO21x1_ASAP7_75t_R _25755_ (.A1(_06924_),
    .A2(_07534_),
    .B(_07535_),
    .Y(_02660_));
 AO221x1_ASAP7_75t_R _25756_ (.A1(net40),
    .A2(_07122_),
    .B1(_07184_),
    .B2(net31),
    .C(_07117_),
    .Y(_07536_));
 INVx1_ASAP7_75t_R _25757_ (.A(_01858_),
    .Y(_07537_));
 INVx1_ASAP7_75t_R _25758_ (.A(_01866_),
    .Y(_07538_));
 AO221x1_ASAP7_75t_R _25759_ (.A1(_07537_),
    .A2(_07122_),
    .B1(_07184_),
    .B2(_07538_),
    .C(_07115_),
    .Y(_07539_));
 NOR2x1_ASAP7_75t_R _25760_ (.A(_01850_),
    .B(_07129_),
    .Y(_07540_));
 AO21x1_ASAP7_75t_R _25761_ (.A1(net48),
    .A2(_05738_),
    .B(_07540_),
    .Y(_07541_));
 AO222x2_ASAP7_75t_R _25762_ (.A1(net54),
    .A2(_07193_),
    .B1(_07536_),
    .B2(_07539_),
    .C1(_07541_),
    .C2(_07128_),
    .Y(_07542_));
 NOR2x1_ASAP7_75t_R _25763_ (.A(_06920_),
    .B(_07542_),
    .Y(_07543_));
 INVx2_ASAP7_75t_R _25764_ (.A(_07071_),
    .Y(_07544_));
 TAPCELL_ASAP7_75t_R TAP_732 ();
 AND3x1_ASAP7_75t_R _25766_ (.A(_06996_),
    .B(_07243_),
    .C(_07246_),
    .Y(_07546_));
 AO21x1_ASAP7_75t_R _25767_ (.A1(_06935_),
    .A2(_07226_),
    .B(_07546_),
    .Y(_07547_));
 OR2x2_ASAP7_75t_R _25768_ (.A(_06935_),
    .B(_07101_),
    .Y(_07548_));
 OA211x2_ASAP7_75t_R _25769_ (.A1(_06996_),
    .A2(_07240_),
    .B(_07548_),
    .C(_06982_),
    .Y(_07549_));
 AO21x2_ASAP7_75t_R _25770_ (.A1(_06932_),
    .A2(_07547_),
    .B(_07549_),
    .Y(_07550_));
 OA21x2_ASAP7_75t_R _25771_ (.A1(_06939_),
    .A2(_07228_),
    .B(_07232_),
    .Y(_07551_));
 AND3x1_ASAP7_75t_R _25772_ (.A(_06935_),
    .B(_07269_),
    .C(_07273_),
    .Y(_07552_));
 AO21x2_ASAP7_75t_R _25773_ (.A1(_06996_),
    .A2(_07551_),
    .B(_07552_),
    .Y(_07553_));
 OR2x2_ASAP7_75t_R _25774_ (.A(_06939_),
    .B(_07261_),
    .Y(_07554_));
 AO32x1_ASAP7_75t_R _25775_ (.A1(_07255_),
    .A2(_07264_),
    .A3(_07554_),
    .B1(_07341_),
    .B2(_07254_),
    .Y(_07555_));
 AOI221x1_ASAP7_75t_R _25776_ (.A1(_07066_),
    .A2(_07550_),
    .B1(_07553_),
    .B2(_07338_),
    .C(_07555_),
    .Y(_07556_));
 OAI21x1_ASAP7_75t_R _25777_ (.A1(_06953_),
    .A2(_06972_),
    .B(_06996_),
    .Y(_07557_));
 NAND2x1_ASAP7_75t_R _25778_ (.A(_06932_),
    .B(_07557_),
    .Y(_07558_));
 AO21x1_ASAP7_75t_R _25779_ (.A1(_06932_),
    .A2(_07016_),
    .B(_07101_),
    .Y(_07559_));
 OAI21x1_ASAP7_75t_R _25780_ (.A1(_07327_),
    .A2(_07558_),
    .B(_07559_),
    .Y(_07560_));
 XOR2x1_ASAP7_75t_R _25781_ (.A(_01387_),
    .Y(_07561_),
    .B(_01385_));
 AO32x2_ASAP7_75t_R _25782_ (.A1(_07076_),
    .A2(_07077_),
    .A3(_07561_),
    .B1(_07080_),
    .B2(_00670_),
    .Y(_07562_));
 INVx1_ASAP7_75t_R _25783_ (.A(_00085_),
    .Y(_07563_));
 NAND2x1_ASAP7_75t_R _25784_ (.A(_00086_),
    .B(_07202_),
    .Y(_07564_));
 OA211x2_ASAP7_75t_R _25785_ (.A1(_07563_),
    .A2(_07202_),
    .B(_07564_),
    .C(_07086_),
    .Y(_07565_));
 AO21x1_ASAP7_75t_R _25786_ (.A1(_02365_),
    .A2(_07206_),
    .B(_07565_),
    .Y(_07566_));
 AO221x1_ASAP7_75t_R _25787_ (.A1(net176),
    .A2(_07097_),
    .B1(_07566_),
    .B2(_07094_),
    .C(_13576_),
    .Y(_07567_));
 INVx1_ASAP7_75t_R _25788_ (.A(_07567_),
    .Y(_07568_));
 AO21x1_ASAP7_75t_R _25789_ (.A1(_13576_),
    .A2(_07562_),
    .B(_07568_),
    .Y(_07569_));
 OAI22x1_ASAP7_75t_R _25790_ (.A1(_01514_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01483_),
    .Y(_07570_));
 OAI22x1_ASAP7_75t_R _25791_ (.A1(_02167_),
    .A2(net284),
    .B1(_07162_),
    .B2(_02061_),
    .Y(_07571_));
 AOI22x1_ASAP7_75t_R _25792_ (.A1(_06884_),
    .A2(_07570_),
    .B1(_07571_),
    .B2(_06886_),
    .Y(_07572_));
 NAND2x1_ASAP7_75t_R _25793_ (.A(net89),
    .B(_07155_),
    .Y(_07573_));
 OA222x2_ASAP7_75t_R _25794_ (.A1(_02024_),
    .A2(_07146_),
    .B1(_07171_),
    .B2(_02093_),
    .C1(_05684_),
    .C2(_06908_),
    .Y(_07574_));
 OA21x2_ASAP7_75t_R _25795_ (.A1(_02134_),
    .A2(_07299_),
    .B(_07574_),
    .Y(_07575_));
 TAPCELL_ASAP7_75t_R TAP_731 ();
 OA222x2_ASAP7_75t_R _25797_ (.A1(_01990_),
    .A2(_07145_),
    .B1(_07149_),
    .B2(_01940_),
    .C1(_00087_),
    .C2(_07305_),
    .Y(_07577_));
 AND4x2_ASAP7_75t_R _25798_ (.A(_07572_),
    .B(_07573_),
    .C(_07575_),
    .D(_07577_),
    .Y(_07578_));
 OA211x2_ASAP7_75t_R _25799_ (.A1(_07430_),
    .A2(_07560_),
    .B(_07569_),
    .C(_07578_),
    .Y(_07579_));
 OA211x2_ASAP7_75t_R _25800_ (.A1(_07544_),
    .A2(_07556_),
    .B(_07579_),
    .C(_06920_),
    .Y(_07580_));
 NOR2x2_ASAP7_75t_R _25801_ (.A(_07543_),
    .B(_07580_),
    .Y(_07581_));
 NOR2x1_ASAP7_75t_R _25802_ (.A(_01704_),
    .B(_06924_),
    .Y(_07582_));
 AO21x1_ASAP7_75t_R _25803_ (.A1(_06924_),
    .A2(_07581_),
    .B(_07582_),
    .Y(_02661_));
 AO21x1_ASAP7_75t_R _25804_ (.A1(_07323_),
    .A2(_07326_),
    .B(_06935_),
    .Y(_07583_));
 OR3x1_ASAP7_75t_R _25805_ (.A(_06996_),
    .B(_07318_),
    .C(_07320_),
    .Y(_07584_));
 AND3x1_ASAP7_75t_R _25806_ (.A(_06932_),
    .B(_07583_),
    .C(_07584_),
    .Y(_07585_));
 AO21x1_ASAP7_75t_R _25807_ (.A1(_06982_),
    .A2(_07216_),
    .B(_07585_),
    .Y(_07586_));
 OA211x2_ASAP7_75t_R _25808_ (.A1(net281),
    .A2(_07018_),
    .B(_07335_),
    .C(_06935_),
    .Y(_07587_));
 AO21x1_ASAP7_75t_R _25809_ (.A1(_06996_),
    .A2(_07317_),
    .B(_07587_),
    .Y(_07588_));
 AO32x1_ASAP7_75t_R _25810_ (.A1(_06928_),
    .A2(_07055_),
    .A3(_07340_),
    .B1(_07334_),
    .B2(_07255_),
    .Y(_07589_));
 AO221x1_ASAP7_75t_R _25811_ (.A1(_07066_),
    .A2(_07586_),
    .B1(_07588_),
    .B2(_07338_),
    .C(_07589_),
    .Y(_07590_));
 OAI21x1_ASAP7_75t_R _25812_ (.A1(_06935_),
    .A2(_07240_),
    .B(_07247_),
    .Y(_07591_));
 NAND2x1_ASAP7_75t_R _25813_ (.A(_07107_),
    .B(_07591_),
    .Y(_07592_));
 INVx1_ASAP7_75t_R _25814_ (.A(_00088_),
    .Y(_07593_));
 NAND2x1_ASAP7_75t_R _25815_ (.A(_00089_),
    .B(_07202_),
    .Y(_07594_));
 OA211x2_ASAP7_75t_R _25816_ (.A1(_07593_),
    .A2(_07202_),
    .B(_07594_),
    .C(_07086_),
    .Y(_07595_));
 AO21x1_ASAP7_75t_R _25817_ (.A1(_02366_),
    .A2(_07206_),
    .B(_07595_),
    .Y(_07596_));
 AOI22x1_ASAP7_75t_R _25818_ (.A1(net177),
    .A2(_07097_),
    .B1(_07596_),
    .B2(_07094_),
    .Y(_07597_));
 INVx1_ASAP7_75t_R _25819_ (.A(_02233_),
    .Y(_07598_));
 AO221x2_ASAP7_75t_R _25820_ (.A1(_07598_),
    .A2(_07078_),
    .B1(_07080_),
    .B2(_00672_),
    .C(_13318_),
    .Y(_07599_));
 OA21x2_ASAP7_75t_R _25821_ (.A1(_13576_),
    .A2(_07597_),
    .B(_07599_),
    .Y(_07600_));
 OAI22x1_ASAP7_75t_R _25822_ (.A1(_01513_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01482_),
    .Y(_07601_));
 OAI22x1_ASAP7_75t_R _25823_ (.A1(_02166_),
    .A2(net284),
    .B1(_07162_),
    .B2(_02060_),
    .Y(_07602_));
 AOI22x1_ASAP7_75t_R _25824_ (.A1(_06884_),
    .A2(_07601_),
    .B1(_07602_),
    .B2(_06886_),
    .Y(_07603_));
 OA21x2_ASAP7_75t_R _25825_ (.A1(_02023_),
    .A2(_07146_),
    .B(_07168_),
    .Y(_07604_));
 OA22x2_ASAP7_75t_R _25826_ (.A1(_02092_),
    .A2(_07171_),
    .B1(_07299_),
    .B2(_02133_),
    .Y(_07605_));
 OA211x2_ASAP7_75t_R _25827_ (.A1(_01712_),
    .A2(_07172_),
    .B(_07604_),
    .C(_07605_),
    .Y(_07606_));
 NAND2x1_ASAP7_75t_R _25828_ (.A(net90),
    .B(_07155_),
    .Y(_07607_));
 OA222x2_ASAP7_75t_R _25829_ (.A1(_01989_),
    .A2(_07145_),
    .B1(_07149_),
    .B2(_01939_),
    .C1(_00090_),
    .C2(_07305_),
    .Y(_07608_));
 AND4x2_ASAP7_75t_R _25830_ (.A(_07603_),
    .B(_07606_),
    .C(_07607_),
    .D(_07608_),
    .Y(_07609_));
 NAND2x2_ASAP7_75t_R _25831_ (.A(_07600_),
    .B(_07609_),
    .Y(_07610_));
 AOI221x1_ASAP7_75t_R _25832_ (.A1(_07071_),
    .A2(_07590_),
    .B1(_07592_),
    .B2(_07109_),
    .C(_07610_),
    .Y(_07611_));
 AO221x1_ASAP7_75t_R _25833_ (.A1(net41),
    .A2(_07122_),
    .B1(_07184_),
    .B2(net32),
    .C(_07117_),
    .Y(_07612_));
 INVx1_ASAP7_75t_R _25834_ (.A(_01857_),
    .Y(_07613_));
 INVx1_ASAP7_75t_R _25835_ (.A(_01865_),
    .Y(_07614_));
 AO221x1_ASAP7_75t_R _25836_ (.A1(_07613_),
    .A2(_07122_),
    .B1(_07184_),
    .B2(_07614_),
    .C(_07115_),
    .Y(_07615_));
 NOR2x1_ASAP7_75t_R _25837_ (.A(_01849_),
    .B(_07129_),
    .Y(_07616_));
 AO21x1_ASAP7_75t_R _25838_ (.A1(net50),
    .A2(_05738_),
    .B(_07616_),
    .Y(_07617_));
 AO222x2_ASAP7_75t_R _25839_ (.A1(net55),
    .A2(_07193_),
    .B1(_07612_),
    .B2(_07615_),
    .C1(_07617_),
    .C2(_07128_),
    .Y(_07618_));
 NOR2x1_ASAP7_75t_R _25840_ (.A(_06920_),
    .B(_07618_),
    .Y(_07619_));
 AOI21x1_ASAP7_75t_R _25841_ (.A1(_06920_),
    .A2(_07611_),
    .B(_07619_),
    .Y(_07620_));
 NOR2x1_ASAP7_75t_R _25842_ (.A(_01703_),
    .B(_06924_),
    .Y(_07621_));
 AO21x1_ASAP7_75t_R _25843_ (.A1(_06924_),
    .A2(net253),
    .B(_07621_),
    .Y(_02662_));
 AO221x1_ASAP7_75t_R _25844_ (.A1(net42),
    .A2(_07122_),
    .B1(_07184_),
    .B2(net33),
    .C(_07117_),
    .Y(_07622_));
 INVx1_ASAP7_75t_R _25845_ (.A(_01856_),
    .Y(_07623_));
 INVx1_ASAP7_75t_R _25846_ (.A(_01864_),
    .Y(_07624_));
 AO221x1_ASAP7_75t_R _25847_ (.A1(_07623_),
    .A2(_07122_),
    .B1(_07184_),
    .B2(_07624_),
    .C(_07115_),
    .Y(_07625_));
 INVx1_ASAP7_75t_R _25848_ (.A(net51),
    .Y(_07626_));
 OAI22x1_ASAP7_75t_R _25849_ (.A1(_07626_),
    .A2(_01730_),
    .B1(_01733_),
    .B2(_07129_),
    .Y(_07627_));
 AO222x2_ASAP7_75t_R _25850_ (.A1(net56),
    .A2(_07193_),
    .B1(_07622_),
    .B2(_07625_),
    .C1(_07627_),
    .C2(_07128_),
    .Y(_07628_));
 OR3x1_ASAP7_75t_R _25851_ (.A(_06939_),
    .B(_07236_),
    .C(_07237_),
    .Y(_07629_));
 OA211x2_ASAP7_75t_R _25852_ (.A1(_06953_),
    .A2(_07405_),
    .B(_07629_),
    .C(_06996_),
    .Y(_07630_));
 AOI21x1_ASAP7_75t_R _25853_ (.A1(_06935_),
    .A2(_07401_),
    .B(_07630_),
    .Y(_07631_));
 NOR2x1_ASAP7_75t_R _25854_ (.A(_06932_),
    .B(_07106_),
    .Y(_07632_));
 AOI21x1_ASAP7_75t_R _25855_ (.A1(_06932_),
    .A2(_07631_),
    .B(_07632_),
    .Y(_07633_));
 OA21x2_ASAP7_75t_R _25856_ (.A1(net281),
    .A2(_07228_),
    .B(_07402_),
    .Y(_07634_));
 AND3x1_ASAP7_75t_R _25857_ (.A(_06935_),
    .B(_07413_),
    .C(_07414_),
    .Y(_07635_));
 AO21x1_ASAP7_75t_R _25858_ (.A1(_06996_),
    .A2(_07634_),
    .B(_07635_),
    .Y(_07636_));
 AO32x1_ASAP7_75t_R _25859_ (.A1(_06928_),
    .A2(_07055_),
    .A3(_07420_),
    .B1(_07412_),
    .B2(_07255_),
    .Y(_07637_));
 AO221x1_ASAP7_75t_R _25860_ (.A1(_07066_),
    .A2(_07633_),
    .B1(_07636_),
    .B2(_07338_),
    .C(_07637_),
    .Y(_07638_));
 TAPCELL_ASAP7_75t_R TAP_730 ();
 OR3x1_ASAP7_75t_R _25862_ (.A(_06982_),
    .B(_06964_),
    .C(_06981_),
    .Y(_07640_));
 AND3x1_ASAP7_75t_R _25863_ (.A(_06928_),
    .B(_06932_),
    .C(_06943_),
    .Y(_07641_));
 INVx1_ASAP7_75t_R _25864_ (.A(_00091_),
    .Y(_07642_));
 TAPCELL_ASAP7_75t_R TAP_729 ();
 NAND2x1_ASAP7_75t_R _25866_ (.A(_00092_),
    .B(_07202_),
    .Y(_07644_));
 OA211x2_ASAP7_75t_R _25867_ (.A1(_07642_),
    .A2(_07202_),
    .B(_07644_),
    .C(_07086_),
    .Y(_07645_));
 AO21x1_ASAP7_75t_R _25868_ (.A1(_02367_),
    .A2(_07206_),
    .B(_07645_),
    .Y(_07646_));
 AOI22x1_ASAP7_75t_R _25869_ (.A1(net178),
    .A2(_07097_),
    .B1(_07646_),
    .B2(_07094_),
    .Y(_07647_));
 TAPCELL_ASAP7_75t_R TAP_728 ();
 TAPCELL_ASAP7_75t_R TAP_727 ();
 XOR2x1_ASAP7_75t_R _25872_ (.A(_01410_),
    .Y(_07650_),
    .B(_02232_));
 NOR2x1_ASAP7_75t_R _25873_ (.A(_07079_),
    .B(_07650_),
    .Y(_07651_));
 AO21x1_ASAP7_75t_R _25874_ (.A1(_00674_),
    .A2(_07079_),
    .B(_07651_),
    .Y(_07652_));
 AO21x1_ASAP7_75t_R _25875_ (.A1(_07076_),
    .A2(_07652_),
    .B(_13318_),
    .Y(_07653_));
 AO21x1_ASAP7_75t_R _25876_ (.A1(_00674_),
    .A2(_05743_),
    .B(_07653_),
    .Y(_07654_));
 OAI22x1_ASAP7_75t_R _25877_ (.A1(_02165_),
    .A2(net284),
    .B1(_07162_),
    .B2(_02059_),
    .Y(_07655_));
 NAND2x1_ASAP7_75t_R _25878_ (.A(_06886_),
    .B(_07655_),
    .Y(_07656_));
 OAI22x1_ASAP7_75t_R _25879_ (.A1(_01512_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01481_),
    .Y(_07657_));
 NAND2x1_ASAP7_75t_R _25880_ (.A(_06884_),
    .B(_07657_),
    .Y(_07658_));
 OR4x2_ASAP7_75t_R _25881_ (.A(_13302_),
    .B(_13658_),
    .C(_13955_),
    .D(_05560_),
    .Y(_07659_));
 TAPCELL_ASAP7_75t_R TAP_726 ();
 OR3x4_ASAP7_75t_R _25883_ (.A(_06911_),
    .B(_06910_),
    .C(_07659_),
    .Y(_07661_));
 INVx1_ASAP7_75t_R _25884_ (.A(net147),
    .Y(_07662_));
 NAND2x2_ASAP7_75t_R _25885_ (.A(_05630_),
    .B(_06889_),
    .Y(_07663_));
 OA222x2_ASAP7_75t_R _25886_ (.A1(_02132_),
    .A2(_07299_),
    .B1(_07661_),
    .B2(_01947_),
    .C1(_07662_),
    .C2(_07663_),
    .Y(_07664_));
 AND3x2_ASAP7_75t_R _25887_ (.A(_07656_),
    .B(_07658_),
    .C(_07664_),
    .Y(_07665_));
 OA21x2_ASAP7_75t_R _25888_ (.A1(_02022_),
    .A2(_07146_),
    .B(_07168_),
    .Y(_07666_));
 OR3x4_ASAP7_75t_R _25889_ (.A(_06911_),
    .B(_06908_),
    .C(_06910_),
    .Y(_07667_));
 OA22x2_ASAP7_75t_R _25890_ (.A1(_01711_),
    .A2(_07172_),
    .B1(_07667_),
    .B2(_01454_),
    .Y(_07668_));
 OA211x2_ASAP7_75t_R _25891_ (.A1(_02091_),
    .A2(_07171_),
    .B(_07666_),
    .C(_07668_),
    .Y(_07669_));
 NAND2x1_ASAP7_75t_R _25892_ (.A(net91),
    .B(_07155_),
    .Y(_07670_));
 OA222x2_ASAP7_75t_R _25893_ (.A1(_01988_),
    .A2(_07145_),
    .B1(_07149_),
    .B2(_01938_),
    .C1(_01574_),
    .C2(_07305_),
    .Y(_07671_));
 AND4x2_ASAP7_75t_R _25894_ (.A(_07665_),
    .B(_07669_),
    .C(_07670_),
    .D(_07671_),
    .Y(_07672_));
 OA211x2_ASAP7_75t_R _25895_ (.A1(_13576_),
    .A2(_07647_),
    .B(_07654_),
    .C(_07672_),
    .Y(_07673_));
 NAND2x1_ASAP7_75t_R _25896_ (.A(_06920_),
    .B(_07673_),
    .Y(_07674_));
 AO221x1_ASAP7_75t_R _25897_ (.A1(_07071_),
    .A2(_07638_),
    .B1(_07640_),
    .B2(_07641_),
    .C(_07674_),
    .Y(_07675_));
 OA21x2_ASAP7_75t_R _25898_ (.A1(_06920_),
    .A2(_07628_),
    .B(_07675_),
    .Y(_07676_));
 NOR2x1_ASAP7_75t_R _25899_ (.A(_01702_),
    .B(_06924_),
    .Y(_07677_));
 AO21x1_ASAP7_75t_R _25900_ (.A1(_06924_),
    .A2(_07676_),
    .B(_07677_),
    .Y(_02663_));
 OR2x4_ASAP7_75t_R _25901_ (.A(_06932_),
    .B(_07101_),
    .Y(_07678_));
 OA31x2_ASAP7_75t_R _25902_ (.A1(_06982_),
    .A2(_06964_),
    .A3(_06981_),
    .B1(_07678_),
    .Y(_07679_));
 OAI21x1_ASAP7_75t_R _25903_ (.A1(_06997_),
    .A2(_07010_),
    .B(_06982_),
    .Y(_07680_));
 NAND2x1_ASAP7_75t_R _25904_ (.A(_06932_),
    .B(_07038_),
    .Y(_07681_));
 AOI21x1_ASAP7_75t_R _25905_ (.A1(_07680_),
    .A2(_07681_),
    .B(_07066_),
    .Y(_07682_));
 AOI21x1_ASAP7_75t_R _25906_ (.A1(_07066_),
    .A2(_07679_),
    .B(_07682_),
    .Y(_07683_));
 OR2x2_ASAP7_75t_R _25907_ (.A(_07544_),
    .B(_07683_),
    .Y(_07684_));
 OR3x1_ASAP7_75t_R _25908_ (.A(_06982_),
    .B(_07430_),
    .C(_07631_),
    .Y(_07685_));
 INVx1_ASAP7_75t_R _25909_ (.A(_02235_),
    .Y(_07686_));
 AOI22x1_ASAP7_75t_R _25910_ (.A1(_07686_),
    .A2(_07078_),
    .B1(_07080_),
    .B2(_00677_),
    .Y(_07687_));
 INVx1_ASAP7_75t_R _25911_ (.A(_00093_),
    .Y(_07688_));
 NAND2x1_ASAP7_75t_R _25912_ (.A(_00094_),
    .B(_07202_),
    .Y(_07689_));
 OA211x2_ASAP7_75t_R _25913_ (.A1(_07688_),
    .A2(_07202_),
    .B(_07689_),
    .C(_07086_),
    .Y(_07690_));
 AO21x1_ASAP7_75t_R _25914_ (.A1(_02368_),
    .A2(net285),
    .B(_07690_),
    .Y(_07691_));
 AO221x1_ASAP7_75t_R _25915_ (.A1(net179),
    .A2(_07097_),
    .B1(_07691_),
    .B2(_07094_),
    .C(_13576_),
    .Y(_07692_));
 AND3x1_ASAP7_75t_R _25916_ (.A(_06982_),
    .B(_07106_),
    .C(_07348_),
    .Y(_07693_));
 OAI22x1_ASAP7_75t_R _25917_ (.A1(net294),
    .A2(_07687_),
    .B1(_07692_),
    .B2(_07693_),
    .Y(_07694_));
 OAI22x1_ASAP7_75t_R _25918_ (.A1(_01511_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01480_),
    .Y(_07695_));
 NAND2x1_ASAP7_75t_R _25919_ (.A(_06884_),
    .B(_07695_),
    .Y(_07696_));
 OAI22x1_ASAP7_75t_R _25920_ (.A1(_02164_),
    .A2(net284),
    .B1(_07162_),
    .B2(_02058_),
    .Y(_07697_));
 NAND2x1_ASAP7_75t_R _25921_ (.A(_06886_),
    .B(_07697_),
    .Y(_07698_));
 AND2x6_ASAP7_75t_R _25922_ (.A(_05538_),
    .B(_06907_),
    .Y(_07699_));
 AOI21x1_ASAP7_75t_R _25923_ (.A1(net92),
    .A2(_06891_),
    .B(_07699_),
    .Y(_07700_));
 OR2x6_ASAP7_75t_R _25924_ (.A(_07507_),
    .B(_07513_),
    .Y(_07701_));
 TAPCELL_ASAP7_75t_R TAP_725 ();
 OA222x2_ASAP7_75t_R _25926_ (.A1(_02090_),
    .A2(_07505_),
    .B1(_07508_),
    .B2(_02131_),
    .C1(_07701_),
    .C2(_01937_),
    .Y(_07703_));
 OA211x2_ASAP7_75t_R _25927_ (.A1(_01987_),
    .A2(_07511_),
    .B(_07700_),
    .C(_07703_),
    .Y(_07704_));
 OR3x4_ASAP7_75t_R _25928_ (.A(_06911_),
    .B(_06910_),
    .C(_06909_),
    .Y(_07705_));
 TAPCELL_ASAP7_75t_R TAP_724 ();
 OA22x2_ASAP7_75t_R _25930_ (.A1(_00095_),
    .A2(_07705_),
    .B1(_07524_),
    .B2(_02021_),
    .Y(_07707_));
 NAND2x2_ASAP7_75t_R _25931_ (.A(_05582_),
    .B(_06892_),
    .Y(_07708_));
 OA22x2_ASAP7_75t_R _25932_ (.A1(_01726_),
    .A2(_07708_),
    .B1(_07516_),
    .B2(_01573_),
    .Y(_07709_));
 AND5x2_ASAP7_75t_R _25933_ (.A(_07696_),
    .B(_07698_),
    .C(_07704_),
    .D(_07707_),
    .E(_07709_),
    .Y(_07710_));
 AND4x2_ASAP7_75t_R _25934_ (.A(_06920_),
    .B(_07685_),
    .C(_07694_),
    .D(_07710_),
    .Y(_07711_));
 TAPCELL_ASAP7_75t_R TAP_723 ();
 TAPCELL_ASAP7_75t_R TAP_722 ();
 TAPCELL_ASAP7_75t_R TAP_721 ();
 OR2x2_ASAP7_75t_R _25938_ (.A(net57),
    .B(_07135_),
    .Y(_07715_));
 OA21x2_ASAP7_75t_R _25939_ (.A1(net420),
    .A2(_07116_),
    .B(_07715_),
    .Y(_07716_));
 TAPCELL_ASAP7_75t_R TAP_720 ();
 INVx1_ASAP7_75t_R _25941_ (.A(_01855_),
    .Y(_07718_));
 OR2x2_ASAP7_75t_R _25942_ (.A(net27),
    .B(net420),
    .Y(_07719_));
 TAPCELL_ASAP7_75t_R TAP_719 ();
 OA211x2_ASAP7_75t_R _25944_ (.A1(_07135_),
    .A2(_07718_),
    .B(_07719_),
    .C(_07120_),
    .Y(_07721_));
 AO21x1_ASAP7_75t_R _25945_ (.A1(_01642_),
    .A2(_07716_),
    .B(_07721_),
    .Y(_07722_));
 OA21x2_ASAP7_75t_R _25946_ (.A1(net43),
    .A2(_07135_),
    .B(_07719_),
    .Y(_07723_));
 TAPCELL_ASAP7_75t_R TAP_718 ();
 OAI21x1_ASAP7_75t_R _25948_ (.A1(net34),
    .A2(net420),
    .B(_07715_),
    .Y(_07725_));
 NAND2x1_ASAP7_75t_R _25949_ (.A(_01642_),
    .B(_07725_),
    .Y(_07726_));
 INVx3_ASAP7_75t_R _25950_ (.A(_01731_),
    .Y(_07727_));
 OA211x2_ASAP7_75t_R _25951_ (.A1(_01642_),
    .A2(_07723_),
    .B(_07726_),
    .C(_07727_),
    .Y(_07728_));
 AND2x2_ASAP7_75t_R _25952_ (.A(net56),
    .B(net420),
    .Y(_07729_));
 AO21x1_ASAP7_75t_R _25953_ (.A1(net33),
    .A2(_07135_),
    .B(_07729_),
    .Y(_07730_));
 NAND2x1_ASAP7_75t_R _25954_ (.A(net418),
    .B(_07730_),
    .Y(_07731_));
 NAND2x1_ASAP7_75t_R _25955_ (.A(net42),
    .B(net420),
    .Y(_07732_));
 NAND2x1_ASAP7_75t_R _25956_ (.A(net51),
    .B(_07135_),
    .Y(_07733_));
 AO21x1_ASAP7_75t_R _25957_ (.A1(_07732_),
    .A2(_07733_),
    .B(net418),
    .Y(_07734_));
 AO21x1_ASAP7_75t_R _25958_ (.A1(_07731_),
    .A2(_07734_),
    .B(_01730_),
    .Y(_07735_));
 OAI21x1_ASAP7_75t_R _25959_ (.A1(_01644_),
    .A2(_07735_),
    .B(_07113_),
    .Y(_07736_));
 AOI211x1_ASAP7_75t_R _25960_ (.A1(_07117_),
    .A2(_07722_),
    .B(_07728_),
    .C(_07736_),
    .Y(_07737_));
 AOI21x1_ASAP7_75t_R _25961_ (.A1(_07684_),
    .A2(_07711_),
    .B(_07737_),
    .Y(_07738_));
 TAPCELL_ASAP7_75t_R TAP_717 ();
 NOR2x1_ASAP7_75t_R _25963_ (.A(_01701_),
    .B(_06924_),
    .Y(_07740_));
 AO21x1_ASAP7_75t_R _25964_ (.A1(_06924_),
    .A2(_07738_),
    .B(_07740_),
    .Y(_02664_));
 INVx1_ASAP7_75t_R _25965_ (.A(net58),
    .Y(_07741_));
 NAND2x1_ASAP7_75t_R _25966_ (.A(_07741_),
    .B(_01643_),
    .Y(_07742_));
 OA21x2_ASAP7_75t_R _25967_ (.A1(net35),
    .A2(_01643_),
    .B(_07742_),
    .Y(_07743_));
 TAPCELL_ASAP7_75t_R TAP_716 ();
 NOR2x1_ASAP7_75t_R _25969_ (.A(net38),
    .B(net420),
    .Y(_07745_));
 AO21x1_ASAP7_75t_R _25970_ (.A1(_07190_),
    .A2(net420),
    .B(_07745_),
    .Y(_07746_));
 NOR2x1_ASAP7_75t_R _25971_ (.A(_01642_),
    .B(_07746_),
    .Y(_07747_));
 AO21x1_ASAP7_75t_R _25972_ (.A1(_01642_),
    .A2(_07743_),
    .B(_07747_),
    .Y(_07748_));
 AOI211x1_ASAP7_75t_R _25973_ (.A1(net420),
    .A2(_01854_),
    .B(_07745_),
    .C(_01642_),
    .Y(_07749_));
 OA211x2_ASAP7_75t_R _25974_ (.A1(_01643_),
    .A2(_07187_),
    .B(_07742_),
    .C(_01642_),
    .Y(_07750_));
 OA21x2_ASAP7_75t_R _25975_ (.A1(_07749_),
    .A2(_07750_),
    .B(_07117_),
    .Y(_07751_));
 AOI211x1_ASAP7_75t_R _25976_ (.A1(_07727_),
    .A2(_07748_),
    .B(_07751_),
    .C(_07736_),
    .Y(_07752_));
 AND3x1_ASAP7_75t_R _25977_ (.A(_06996_),
    .B(_07269_),
    .C(_07273_),
    .Y(_07753_));
 OA21x2_ASAP7_75t_R _25978_ (.A1(_07266_),
    .A2(_07753_),
    .B(_07107_),
    .Y(_07754_));
 AOI21x1_ASAP7_75t_R _25979_ (.A1(_07234_),
    .A2(_07338_),
    .B(_07754_),
    .Y(_07755_));
 NAND2x1_ASAP7_75t_R _25980_ (.A(_07066_),
    .B(_07678_),
    .Y(_07756_));
 AO21x1_ASAP7_75t_R _25981_ (.A1(_06932_),
    .A2(_07591_),
    .B(_07756_),
    .Y(_07757_));
 AO21x1_ASAP7_75t_R _25982_ (.A1(_07755_),
    .A2(_07757_),
    .B(_07544_),
    .Y(_07758_));
 XNOR2x2_ASAP7_75t_R _25983_ (.A(_01426_),
    .B(_02234_),
    .Y(_07759_));
 AND3x1_ASAP7_75t_R _25984_ (.A(_00279_),
    .B(_07077_),
    .C(_07759_),
    .Y(_07760_));
 AO21x1_ASAP7_75t_R _25985_ (.A1(_00680_),
    .A2(_07196_),
    .B(_07760_),
    .Y(_07761_));
 INVx1_ASAP7_75t_R _25986_ (.A(_00096_),
    .Y(_07762_));
 NAND2x1_ASAP7_75t_R _25987_ (.A(_00097_),
    .B(_07202_),
    .Y(_07763_));
 OA211x2_ASAP7_75t_R _25988_ (.A1(_07762_),
    .A2(_07202_),
    .B(_07763_),
    .C(_07086_),
    .Y(_07764_));
 AO21x1_ASAP7_75t_R _25989_ (.A1(_02369_),
    .A2(net285),
    .B(_07764_),
    .Y(_07765_));
 AO221x1_ASAP7_75t_R _25990_ (.A1(net180),
    .A2(_07097_),
    .B1(_07765_),
    .B2(_07094_),
    .C(_13576_),
    .Y(_07766_));
 INVx1_ASAP7_75t_R _25991_ (.A(_07766_),
    .Y(_07767_));
 AO21x1_ASAP7_75t_R _25992_ (.A1(_13576_),
    .A2(_07761_),
    .B(_07767_),
    .Y(_07768_));
 OAI22x1_ASAP7_75t_R _25993_ (.A1(_01510_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01479_),
    .Y(_07769_));
 OAI22x1_ASAP7_75t_R _25994_ (.A1(_02163_),
    .A2(net284),
    .B1(_07162_),
    .B2(_02057_),
    .Y(_07770_));
 AOI22x1_ASAP7_75t_R _25995_ (.A1(_06884_),
    .A2(_07769_),
    .B1(_07770_),
    .B2(_06886_),
    .Y(_07771_));
 OA22x2_ASAP7_75t_R _25996_ (.A1(_02020_),
    .A2(_07146_),
    .B1(_07305_),
    .B2(_01572_),
    .Y(_07772_));
 OA22x2_ASAP7_75t_R _25997_ (.A1(_01986_),
    .A2(_07145_),
    .B1(_07149_),
    .B2(_01936_),
    .Y(_07773_));
 NAND2x1_ASAP7_75t_R _25998_ (.A(net93),
    .B(_07155_),
    .Y(_07774_));
 OA222x2_ASAP7_75t_R _25999_ (.A1(_00098_),
    .A2(_07151_),
    .B1(_07299_),
    .B2(_02130_),
    .C1(_05684_),
    .C2(_06908_),
    .Y(_07775_));
 OA21x2_ASAP7_75t_R _26000_ (.A1(_02089_),
    .A2(_07171_),
    .B(_07775_),
    .Y(_07776_));
 AND5x2_ASAP7_75t_R _26001_ (.A(_07771_),
    .B(_07772_),
    .C(_07773_),
    .D(_07774_),
    .E(_07776_),
    .Y(_07777_));
 NAND2x1_ASAP7_75t_R _26002_ (.A(_07348_),
    .B(_07586_),
    .Y(_07778_));
 AND5x2_ASAP7_75t_R _26003_ (.A(_06920_),
    .B(_07758_),
    .C(_07768_),
    .D(_07777_),
    .E(_07778_),
    .Y(_07779_));
 NOR2x2_ASAP7_75t_R _26004_ (.A(_07752_),
    .B(_07779_),
    .Y(_07780_));
 NOR2x1_ASAP7_75t_R _26005_ (.A(_01700_),
    .B(_06924_),
    .Y(_07781_));
 AO21x1_ASAP7_75t_R _26006_ (.A1(_06924_),
    .A2(_07780_),
    .B(_07781_),
    .Y(_02665_));
 TAPCELL_ASAP7_75t_R TAP_715 ();
 OA211x2_ASAP7_75t_R _26008_ (.A1(_07327_),
    .A2(_07558_),
    .B(_07559_),
    .C(_07066_),
    .Y(_07783_));
 AO221x1_ASAP7_75t_R _26009_ (.A1(_07107_),
    .A2(_07337_),
    .B1(_07338_),
    .B2(_07322_),
    .C(_07783_),
    .Y(_07784_));
 INVx1_ASAP7_75t_R _26010_ (.A(_00099_),
    .Y(_07785_));
 NAND2x1_ASAP7_75t_R _26011_ (.A(_00100_),
    .B(_07202_),
    .Y(_07786_));
 OA211x2_ASAP7_75t_R _26012_ (.A1(_07785_),
    .A2(_07202_),
    .B(_07786_),
    .C(_07086_),
    .Y(_07787_));
 AO21x1_ASAP7_75t_R _26013_ (.A1(_02370_),
    .A2(net285),
    .B(_07787_),
    .Y(_07788_));
 AOI221x1_ASAP7_75t_R _26014_ (.A1(net151),
    .A2(_07097_),
    .B1(_07788_),
    .B2(_07094_),
    .C(_13576_),
    .Y(_07789_));
 INVx1_ASAP7_75t_R _26015_ (.A(_02237_),
    .Y(_07790_));
 AO21x1_ASAP7_75t_R _26016_ (.A1(_07790_),
    .A2(_07078_),
    .B(_00682_),
    .Y(_07791_));
 OA211x2_ASAP7_75t_R _26017_ (.A1(_07790_),
    .A2(_07080_),
    .B(_07791_),
    .C(_13576_),
    .Y(_07792_));
 OAI22x1_ASAP7_75t_R _26018_ (.A1(_01509_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01478_),
    .Y(_07793_));
 OAI22x1_ASAP7_75t_R _26019_ (.A1(_02162_),
    .A2(net284),
    .B1(_07162_),
    .B2(_02056_),
    .Y(_07794_));
 AOI22x1_ASAP7_75t_R _26020_ (.A1(_06884_),
    .A2(_07793_),
    .B1(_07794_),
    .B2(_06886_),
    .Y(_07795_));
 OA22x2_ASAP7_75t_R _26021_ (.A1(_02019_),
    .A2(_07146_),
    .B1(_07305_),
    .B2(_01571_),
    .Y(_07796_));
 OA22x2_ASAP7_75t_R _26022_ (.A1(_01985_),
    .A2(_07145_),
    .B1(_07149_),
    .B2(_01935_),
    .Y(_07797_));
 NAND2x1_ASAP7_75t_R _26023_ (.A(net63),
    .B(_07155_),
    .Y(_07798_));
 OA222x2_ASAP7_75t_R _26024_ (.A1(_00101_),
    .A2(_07151_),
    .B1(_07299_),
    .B2(_02129_),
    .C1(_05684_),
    .C2(_06908_),
    .Y(_07799_));
 OA21x2_ASAP7_75t_R _26025_ (.A1(_02088_),
    .A2(_07171_),
    .B(_07799_),
    .Y(_07800_));
 AND5x2_ASAP7_75t_R _26026_ (.A(_07795_),
    .B(_07796_),
    .C(_07797_),
    .D(_07798_),
    .E(_07800_),
    .Y(_07801_));
 OA21x2_ASAP7_75t_R _26027_ (.A1(_07789_),
    .A2(_07792_),
    .B(_07801_),
    .Y(_07802_));
 NAND2x1_ASAP7_75t_R _26028_ (.A(_06920_),
    .B(_07802_),
    .Y(_07803_));
 AO221x1_ASAP7_75t_R _26029_ (.A1(_07348_),
    .A2(_07550_),
    .B1(_07784_),
    .B2(_07071_),
    .C(_07803_),
    .Y(_07804_));
 OR2x2_ASAP7_75t_R _26030_ (.A(net49),
    .B(net419),
    .Y(_07805_));
 OA21x2_ASAP7_75t_R _26031_ (.A1(net45),
    .A2(_07135_),
    .B(_07805_),
    .Y(_07806_));
 OR2x2_ASAP7_75t_R _26032_ (.A(net28),
    .B(_07135_),
    .Y(_07807_));
 OAI21x1_ASAP7_75t_R _26033_ (.A1(net36),
    .A2(net419),
    .B(_07807_),
    .Y(_07808_));
 NAND2x1_ASAP7_75t_R _26034_ (.A(net418),
    .B(_07808_),
    .Y(_07809_));
 OA211x2_ASAP7_75t_R _26035_ (.A1(net418),
    .A2(_07806_),
    .B(_07809_),
    .C(_07727_),
    .Y(_07810_));
 INVx1_ASAP7_75t_R _26036_ (.A(_01853_),
    .Y(_07811_));
 OA211x2_ASAP7_75t_R _26037_ (.A1(_07135_),
    .A2(_07811_),
    .B(_07805_),
    .C(_07120_),
    .Y(_07812_));
 INVx1_ASAP7_75t_R _26038_ (.A(_01861_),
    .Y(_07813_));
 OA211x2_ASAP7_75t_R _26039_ (.A1(net419),
    .A2(_07813_),
    .B(_07807_),
    .C(net418),
    .Y(_07814_));
 OA21x2_ASAP7_75t_R _26040_ (.A1(_07812_),
    .A2(_07814_),
    .B(_07117_),
    .Y(_07815_));
 OR3x1_ASAP7_75t_R _26041_ (.A(_07736_),
    .B(_07810_),
    .C(_07815_),
    .Y(_07816_));
 AND2x6_ASAP7_75t_R _26042_ (.A(_07804_),
    .B(_07816_),
    .Y(_07817_));
 NOR2x1_ASAP7_75t_R _26043_ (.A(_01699_),
    .B(_06924_),
    .Y(_07818_));
 AO21x1_ASAP7_75t_R _26044_ (.A1(_06924_),
    .A2(_07817_),
    .B(_07818_),
    .Y(_02666_));
 OA21x2_ASAP7_75t_R _26045_ (.A1(_07482_),
    .A2(_07483_),
    .B(_07481_),
    .Y(_07819_));
 NAND2x1_ASAP7_75t_R _26046_ (.A(_06928_),
    .B(_06982_),
    .Y(_07820_));
 INVx1_ASAP7_75t_R _26047_ (.A(_07404_),
    .Y(_07821_));
 OA21x2_ASAP7_75t_R _26048_ (.A1(_06982_),
    .A2(_07408_),
    .B(_07678_),
    .Y(_07822_));
 OA222x2_ASAP7_75t_R _26049_ (.A1(_07820_),
    .A2(_07821_),
    .B1(_07416_),
    .B2(_07100_),
    .C1(_06928_),
    .C2(_07822_),
    .Y(_07823_));
 XOR2x1_ASAP7_75t_R _26050_ (.A(_01436_),
    .Y(_07824_),
    .B(_02236_));
 NOR2x1_ASAP7_75t_R _26051_ (.A(_07079_),
    .B(_07824_),
    .Y(_07825_));
 AO21x1_ASAP7_75t_R _26052_ (.A1(_00684_),
    .A2(_07079_),
    .B(_07825_),
    .Y(_07826_));
 AND2x2_ASAP7_75t_R _26053_ (.A(_07076_),
    .B(_07826_),
    .Y(_07827_));
 AO21x2_ASAP7_75t_R _26054_ (.A1(_00684_),
    .A2(_05743_),
    .B(_07827_),
    .Y(_07828_));
 INVx1_ASAP7_75t_R _26055_ (.A(_00102_),
    .Y(_07829_));
 NAND2x1_ASAP7_75t_R _26056_ (.A(_00103_),
    .B(_07202_),
    .Y(_07830_));
 OA211x2_ASAP7_75t_R _26057_ (.A1(_07829_),
    .A2(_07202_),
    .B(_07830_),
    .C(_07086_),
    .Y(_07831_));
 AO21x1_ASAP7_75t_R _26058_ (.A1(_02371_),
    .A2(_07206_),
    .B(_07831_),
    .Y(_07832_));
 AO221x1_ASAP7_75t_R _26059_ (.A1(net152),
    .A2(_07097_),
    .B1(_07832_),
    .B2(_07094_),
    .C(_13576_),
    .Y(_07833_));
 INVx1_ASAP7_75t_R _26060_ (.A(_07833_),
    .Y(_07834_));
 AO21x1_ASAP7_75t_R _26061_ (.A1(_13576_),
    .A2(_07828_),
    .B(_07834_),
    .Y(_07835_));
 OAI22x1_ASAP7_75t_R _26062_ (.A1(_02161_),
    .A2(net284),
    .B1(_07162_),
    .B2(_02055_),
    .Y(_07836_));
 NAND2x1_ASAP7_75t_R _26063_ (.A(_06886_),
    .B(_07836_),
    .Y(_07837_));
 OAI22x1_ASAP7_75t_R _26064_ (.A1(_01508_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01477_),
    .Y(_07838_));
 NAND2x1_ASAP7_75t_R _26065_ (.A(_06884_),
    .B(_07838_),
    .Y(_07839_));
 OA22x2_ASAP7_75t_R _26066_ (.A1(_01934_),
    .A2(_07701_),
    .B1(_07508_),
    .B2(_02128_),
    .Y(_07840_));
 NOR2x2_ASAP7_75t_R _26067_ (.A(_07507_),
    .B(_07659_),
    .Y(_07841_));
 NAND2x1_ASAP7_75t_R _26068_ (.A(net129),
    .B(_07841_),
    .Y(_07842_));
 OA211x2_ASAP7_75t_R _26069_ (.A1(_02018_),
    .A2(_07524_),
    .B(_07840_),
    .C(_07842_),
    .Y(_07843_));
 OA222x2_ASAP7_75t_R _26070_ (.A1(_00657_),
    .A2(_07705_),
    .B1(_07661_),
    .B2(_01948_),
    .C1(_02087_),
    .C2(_07505_),
    .Y(_07844_));
 OA211x2_ASAP7_75t_R _26071_ (.A1(_01570_),
    .A2(_07516_),
    .B(_07843_),
    .C(_07844_),
    .Y(_07845_));
 OA22x2_ASAP7_75t_R _26072_ (.A1(_02033_),
    .A2(_07708_),
    .B1(_07667_),
    .B2(_01456_),
    .Y(_07846_));
 OA211x2_ASAP7_75t_R _26073_ (.A1(_01984_),
    .A2(_07511_),
    .B(_07846_),
    .C(_07168_),
    .Y(_07847_));
 NAND2x1_ASAP7_75t_R _26074_ (.A(net64),
    .B(_06891_),
    .Y(_07848_));
 AND5x2_ASAP7_75t_R _26075_ (.A(_07837_),
    .B(_07839_),
    .C(_07845_),
    .D(_07847_),
    .E(_07848_),
    .Y(_07849_));
 NAND3x2_ASAP7_75t_R _26076_ (.B(_07835_),
    .C(_07849_),
    .Y(_07850_),
    .A(_06920_));
 AO221x1_ASAP7_75t_R _26077_ (.A1(_07348_),
    .A2(_07819_),
    .B1(_07823_),
    .B2(_07071_),
    .C(_07850_),
    .Y(_07851_));
 OR2x2_ASAP7_75t_R _26078_ (.A(net52),
    .B(net420),
    .Y(_07852_));
 OA21x2_ASAP7_75t_R _26079_ (.A1(net46),
    .A2(_07135_),
    .B(_07852_),
    .Y(_07853_));
 INVx1_ASAP7_75t_R _26080_ (.A(net29),
    .Y(_07854_));
 NAND2x1_ASAP7_75t_R _26081_ (.A(_07854_),
    .B(net420),
    .Y(_07855_));
 OAI21x1_ASAP7_75t_R _26082_ (.A1(net37),
    .A2(net420),
    .B(_07855_),
    .Y(_07856_));
 NAND2x1_ASAP7_75t_R _26083_ (.A(_01642_),
    .B(_07856_),
    .Y(_07857_));
 OA211x2_ASAP7_75t_R _26084_ (.A1(_01642_),
    .A2(_07853_),
    .B(_07857_),
    .C(_07727_),
    .Y(_07858_));
 INVx1_ASAP7_75t_R _26085_ (.A(_01852_),
    .Y(_07859_));
 OA211x2_ASAP7_75t_R _26086_ (.A1(_07135_),
    .A2(_07859_),
    .B(_07852_),
    .C(_07120_),
    .Y(_07860_));
 INVx1_ASAP7_75t_R _26087_ (.A(_01860_),
    .Y(_07861_));
 OA211x2_ASAP7_75t_R _26088_ (.A1(net420),
    .A2(_07861_),
    .B(_07855_),
    .C(_01642_),
    .Y(_07862_));
 OA21x2_ASAP7_75t_R _26089_ (.A1(_07860_),
    .A2(_07862_),
    .B(_07117_),
    .Y(_07863_));
 OR3x1_ASAP7_75t_R _26090_ (.A(_07736_),
    .B(_07858_),
    .C(_07863_),
    .Y(_07864_));
 AND2x6_ASAP7_75t_R _26091_ (.A(_07851_),
    .B(_07864_),
    .Y(_07865_));
 NOR2x1_ASAP7_75t_R _26092_ (.A(_01698_),
    .B(_06924_),
    .Y(_07866_));
 AO21x1_ASAP7_75t_R _26093_ (.A1(_06924_),
    .A2(_07865_),
    .B(_07866_),
    .Y(_02667_));
 AND2x2_ASAP7_75t_R _26094_ (.A(_07479_),
    .B(_07480_),
    .Y(_07867_));
 NAND2x1_ASAP7_75t_R _26095_ (.A(_07066_),
    .B(_07432_),
    .Y(_07868_));
 OR3x1_ASAP7_75t_R _26096_ (.A(_07100_),
    .B(_07486_),
    .C(_07487_),
    .Y(_07869_));
 OA211x2_ASAP7_75t_R _26097_ (.A1(_07820_),
    .A2(_07867_),
    .B(_07868_),
    .C(_07869_),
    .Y(_07870_));
 AND2x2_ASAP7_75t_R _26098_ (.A(_07071_),
    .B(_07870_),
    .Y(_07871_));
 INVx1_ASAP7_75t_R _26099_ (.A(_02239_),
    .Y(_07872_));
 AO32x2_ASAP7_75t_R _26100_ (.A1(_07872_),
    .A2(_07076_),
    .A3(_07077_),
    .B1(_07080_),
    .B2(_00686_),
    .Y(_07873_));
 INVx1_ASAP7_75t_R _26101_ (.A(_00104_),
    .Y(_07874_));
 NAND2x1_ASAP7_75t_R _26102_ (.A(_00105_),
    .B(_07202_),
    .Y(_07875_));
 OA211x2_ASAP7_75t_R _26103_ (.A1(_07874_),
    .A2(_07202_),
    .B(_07875_),
    .C(_07086_),
    .Y(_07876_));
 AO21x1_ASAP7_75t_R _26104_ (.A1(_02372_),
    .A2(_07206_),
    .B(_07876_),
    .Y(_07877_));
 AO221x1_ASAP7_75t_R _26105_ (.A1(net153),
    .A2(_07097_),
    .B1(_07877_),
    .B2(_07094_),
    .C(_13576_),
    .Y(_07878_));
 INVx1_ASAP7_75t_R _26106_ (.A(_07878_),
    .Y(_07879_));
 AO21x1_ASAP7_75t_R _26107_ (.A1(_13576_),
    .A2(_07873_),
    .B(_07879_),
    .Y(_07880_));
 TAPCELL_ASAP7_75t_R TAP_714 ();
 TAPCELL_ASAP7_75t_R TAP_713 ();
 OAI22x1_ASAP7_75t_R _26110_ (.A1(_02160_),
    .A2(net284),
    .B1(_07162_),
    .B2(_02054_),
    .Y(_07883_));
 NAND2x1_ASAP7_75t_R _26111_ (.A(_06886_),
    .B(_07883_),
    .Y(_07884_));
 OAI22x1_ASAP7_75t_R _26112_ (.A1(_01507_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01476_),
    .Y(_07885_));
 NAND2x1_ASAP7_75t_R _26113_ (.A(_06884_),
    .B(_07885_),
    .Y(_07886_));
 OA222x2_ASAP7_75t_R _26114_ (.A1(_00656_),
    .A2(_07705_),
    .B1(_07701_),
    .B2(_01933_),
    .C1(_07516_),
    .C2(_01569_),
    .Y(_07887_));
 OR3x1_ASAP7_75t_R _26115_ (.A(_02127_),
    .B(_06908_),
    .C(_07507_),
    .Y(_07888_));
 OA22x2_ASAP7_75t_R _26116_ (.A1(_02017_),
    .A2(_07524_),
    .B1(_07667_),
    .B2(_01455_),
    .Y(_07889_));
 OA211x2_ASAP7_75t_R _26117_ (.A1(_02032_),
    .A2(_07708_),
    .B(_07888_),
    .C(_07889_),
    .Y(_07890_));
 OAI22x1_ASAP7_75t_R _26118_ (.A1(_02086_),
    .A2(_07520_),
    .B1(_07523_),
    .B2(_01983_),
    .Y(_07891_));
 AO221x1_ASAP7_75t_R _26119_ (.A1(net65),
    .A2(_06891_),
    .B1(_07891_),
    .B2(_06892_),
    .C(_07699_),
    .Y(_07892_));
 INVx1_ASAP7_75t_R _26120_ (.A(_07892_),
    .Y(_07893_));
 AND5x2_ASAP7_75t_R _26121_ (.A(_07884_),
    .B(_07886_),
    .C(_07887_),
    .D(_07890_),
    .E(_07893_),
    .Y(_07894_));
 AND3x2_ASAP7_75t_R _26122_ (.A(_06920_),
    .B(_07880_),
    .C(_07894_),
    .Y(_07895_));
 OAI21x1_ASAP7_75t_R _26123_ (.A1(_07430_),
    .A2(_07410_),
    .B(_07895_),
    .Y(_07896_));
 OR2x2_ASAP7_75t_R _26124_ (.A(net53),
    .B(net419),
    .Y(_07897_));
 OA21x2_ASAP7_75t_R _26125_ (.A1(net47),
    .A2(_07135_),
    .B(_07897_),
    .Y(_07898_));
 OR2x2_ASAP7_75t_R _26126_ (.A(net30),
    .B(_07135_),
    .Y(_07899_));
 OAI21x1_ASAP7_75t_R _26127_ (.A1(net39),
    .A2(net419),
    .B(_07899_),
    .Y(_07900_));
 NAND2x1_ASAP7_75t_R _26128_ (.A(net418),
    .B(_07900_),
    .Y(_07901_));
 OA211x2_ASAP7_75t_R _26129_ (.A1(net418),
    .A2(_07898_),
    .B(_07901_),
    .C(_07727_),
    .Y(_07902_));
 INVx1_ASAP7_75t_R _26130_ (.A(_01851_),
    .Y(_07903_));
 OA211x2_ASAP7_75t_R _26131_ (.A1(_07135_),
    .A2(_07903_),
    .B(_07897_),
    .C(_07120_),
    .Y(_07904_));
 OA211x2_ASAP7_75t_R _26132_ (.A1(net419),
    .A2(_07473_),
    .B(_07899_),
    .C(net418),
    .Y(_07905_));
 OA21x2_ASAP7_75t_R _26133_ (.A1(_07904_),
    .A2(_07905_),
    .B(_07117_),
    .Y(_07906_));
 OR3x1_ASAP7_75t_R _26134_ (.A(_07736_),
    .B(_07902_),
    .C(_07906_),
    .Y(_07907_));
 OA21x2_ASAP7_75t_R _26135_ (.A1(_07871_),
    .A2(_07896_),
    .B(_07907_),
    .Y(_07908_));
 NOR2x1_ASAP7_75t_R _26136_ (.A(_01697_),
    .B(_06924_),
    .Y(_07909_));
 AO21x1_ASAP7_75t_R _26137_ (.A1(_06924_),
    .A2(_07908_),
    .B(_07909_),
    .Y(_02668_));
 INVx1_ASAP7_75t_R _26138_ (.A(_00106_),
    .Y(_07910_));
 NAND2x1_ASAP7_75t_R _26139_ (.A(_00107_),
    .B(_07202_),
    .Y(_07911_));
 OA211x2_ASAP7_75t_R _26140_ (.A1(_07910_),
    .A2(_07202_),
    .B(_07911_),
    .C(_07086_),
    .Y(_07912_));
 AO21x1_ASAP7_75t_R _26141_ (.A1(_02373_),
    .A2(net285),
    .B(_07912_),
    .Y(_07913_));
 AOI22x1_ASAP7_75t_R _26142_ (.A1(net154),
    .A2(_07097_),
    .B1(_07913_),
    .B2(_07094_),
    .Y(_07914_));
 TAPCELL_ASAP7_75t_R TAP_712 ();
 XOR2x2_ASAP7_75t_R _26144_ (.A(_00015_),
    .B(_02238_),
    .Y(_07916_));
 NAND2x1_ASAP7_75t_R _26145_ (.A(_00718_),
    .B(_07079_),
    .Y(_07917_));
 OA21x2_ASAP7_75t_R _26146_ (.A1(_07079_),
    .A2(_07916_),
    .B(_07917_),
    .Y(_07918_));
 OA21x2_ASAP7_75t_R _26147_ (.A1(_05745_),
    .A2(_07918_),
    .B(_13576_),
    .Y(_07919_));
 INVx1_ASAP7_75t_R _26148_ (.A(_07919_),
    .Y(_07920_));
 AO21x1_ASAP7_75t_R _26149_ (.A1(_00718_),
    .A2(_05743_),
    .B(_07920_),
    .Y(_07921_));
 OAI22x1_ASAP7_75t_R _26150_ (.A1(_01506_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01475_),
    .Y(_07922_));
 NAND2x1_ASAP7_75t_R _26151_ (.A(_06884_),
    .B(_07922_),
    .Y(_07923_));
 OAI22x1_ASAP7_75t_R _26152_ (.A1(_02159_),
    .A2(net284),
    .B1(_07162_),
    .B2(_02053_),
    .Y(_07924_));
 NAND2x1_ASAP7_75t_R _26153_ (.A(_06886_),
    .B(_07924_),
    .Y(_07925_));
 NAND2x1_ASAP7_75t_R _26154_ (.A(net66),
    .B(_06891_),
    .Y(_07926_));
 OA21x2_ASAP7_75t_R _26155_ (.A1(_02016_),
    .A2(_07524_),
    .B(_07168_),
    .Y(_07927_));
 OA22x2_ASAP7_75t_R _26156_ (.A1(_01982_),
    .A2(_07511_),
    .B1(_07701_),
    .B2(_01932_),
    .Y(_07928_));
 OA22x2_ASAP7_75t_R _26157_ (.A1(_02031_),
    .A2(_07708_),
    .B1(_07508_),
    .B2(_02126_),
    .Y(_07929_));
 AND4x1_ASAP7_75t_R _26158_ (.A(_07926_),
    .B(_07927_),
    .C(_07928_),
    .D(_07929_),
    .Y(_07930_));
 OA222x2_ASAP7_75t_R _26159_ (.A1(_00108_),
    .A2(_07705_),
    .B1(_07516_),
    .B2(_01568_),
    .C1(_02085_),
    .C2(_07505_),
    .Y(_07931_));
 AND4x2_ASAP7_75t_R _26160_ (.A(_07923_),
    .B(_07925_),
    .C(_07930_),
    .D(_07931_),
    .Y(_07932_));
 OA211x2_ASAP7_75t_R _26161_ (.A1(_13576_),
    .A2(_07914_),
    .B(_07921_),
    .C(_07932_),
    .Y(_07933_));
 NAND2x1_ASAP7_75t_R _26162_ (.A(_06920_),
    .B(_07933_),
    .Y(_07934_));
 TAPCELL_ASAP7_75t_R TAP_711 ();
 OA222x2_ASAP7_75t_R _26164_ (.A1(_06928_),
    .A2(_07347_),
    .B1(_07547_),
    .B2(_07820_),
    .C1(_07553_),
    .C2(_07100_),
    .Y(_07936_));
 AO32x1_ASAP7_75t_R _26165_ (.A1(_06928_),
    .A2(_06943_),
    .A3(_07331_),
    .B1(_07936_),
    .B2(_07071_),
    .Y(_07937_));
 OR2x2_ASAP7_75t_R _26166_ (.A(net54),
    .B(net420),
    .Y(_07938_));
 OA21x2_ASAP7_75t_R _26167_ (.A1(net48),
    .A2(_07135_),
    .B(_07938_),
    .Y(_07939_));
 INVx1_ASAP7_75t_R _26168_ (.A(net31),
    .Y(_07940_));
 NAND2x1_ASAP7_75t_R _26169_ (.A(_07940_),
    .B(net420),
    .Y(_07941_));
 OAI21x1_ASAP7_75t_R _26170_ (.A1(net40),
    .A2(net420),
    .B(_07941_),
    .Y(_07942_));
 NAND2x1_ASAP7_75t_R _26171_ (.A(_01642_),
    .B(_07942_),
    .Y(_07943_));
 OA211x2_ASAP7_75t_R _26172_ (.A1(_01642_),
    .A2(_07939_),
    .B(_07943_),
    .C(_07727_),
    .Y(_07944_));
 INVx1_ASAP7_75t_R _26173_ (.A(_01850_),
    .Y(_07945_));
 OA211x2_ASAP7_75t_R _26174_ (.A1(_07135_),
    .A2(_07945_),
    .B(_07938_),
    .C(_07120_),
    .Y(_07946_));
 OA211x2_ASAP7_75t_R _26175_ (.A1(net420),
    .A2(_07537_),
    .B(_07941_),
    .C(_01642_),
    .Y(_07947_));
 OA21x2_ASAP7_75t_R _26176_ (.A1(_07946_),
    .A2(_07947_),
    .B(_07117_),
    .Y(_07948_));
 OR3x1_ASAP7_75t_R _26177_ (.A(_07736_),
    .B(_07944_),
    .C(_07948_),
    .Y(_07949_));
 OA21x2_ASAP7_75t_R _26178_ (.A1(_07934_),
    .A2(_07937_),
    .B(_07949_),
    .Y(_07950_));
 NOR2x1_ASAP7_75t_R _26179_ (.A(_01696_),
    .B(_06924_),
    .Y(_07951_));
 AO21x1_ASAP7_75t_R _26180_ (.A1(_06924_),
    .A2(_07950_),
    .B(_07951_),
    .Y(_02669_));
 NAND2x1_ASAP7_75t_R _26181_ (.A(_06982_),
    .B(_07591_),
    .Y(_07952_));
 OA211x2_ASAP7_75t_R _26182_ (.A1(_06982_),
    .A2(_07234_),
    .B(_07952_),
    .C(_07348_),
    .Y(_07953_));
 AND3x1_ASAP7_75t_R _26183_ (.A(_00279_),
    .B(_02241_),
    .C(_07077_),
    .Y(_07954_));
 AO21x1_ASAP7_75t_R _26184_ (.A1(_06787_),
    .A2(_07196_),
    .B(_07954_),
    .Y(_07955_));
 INVx1_ASAP7_75t_R _26185_ (.A(_00109_),
    .Y(_07956_));
 NAND2x1_ASAP7_75t_R _26186_ (.A(_00110_),
    .B(_07202_),
    .Y(_07957_));
 OA211x2_ASAP7_75t_R _26187_ (.A1(_07956_),
    .A2(_07202_),
    .B(_07957_),
    .C(_07086_),
    .Y(_07958_));
 AO21x1_ASAP7_75t_R _26188_ (.A1(_02374_),
    .A2(net285),
    .B(_07958_),
    .Y(_07959_));
 AO221x1_ASAP7_75t_R _26189_ (.A1(net155),
    .A2(_07097_),
    .B1(_07959_),
    .B2(_07094_),
    .C(_13576_),
    .Y(_07960_));
 OA21x2_ASAP7_75t_R _26190_ (.A1(net294),
    .A2(_07955_),
    .B(_07960_),
    .Y(_07961_));
 OAI22x1_ASAP7_75t_R _26191_ (.A1(_01505_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01474_),
    .Y(_07962_));
 OAI22x1_ASAP7_75t_R _26192_ (.A1(_02158_),
    .A2(net284),
    .B1(_07162_),
    .B2(_02052_),
    .Y(_07963_));
 AOI22x1_ASAP7_75t_R _26193_ (.A1(_06884_),
    .A2(_07962_),
    .B1(_07963_),
    .B2(_06886_),
    .Y(_07964_));
 OA222x2_ASAP7_75t_R _26194_ (.A1(_00111_),
    .A2(_07151_),
    .B1(_07299_),
    .B2(_02125_),
    .C1(_05684_),
    .C2(_06908_),
    .Y(_07965_));
 OA22x2_ASAP7_75t_R _26195_ (.A1(_01981_),
    .A2(_07145_),
    .B1(_07305_),
    .B2(_01567_),
    .Y(_07966_));
 OA22x2_ASAP7_75t_R _26196_ (.A1(_02015_),
    .A2(_07146_),
    .B1(_07149_),
    .B2(_01931_),
    .Y(_07967_));
 NAND2x1_ASAP7_75t_R _26197_ (.A(net67),
    .B(_07155_),
    .Y(_07968_));
 OA21x2_ASAP7_75t_R _26198_ (.A1(_02084_),
    .A2(_07171_),
    .B(_07968_),
    .Y(_07969_));
 AND5x2_ASAP7_75t_R _26199_ (.A(_07964_),
    .B(_07965_),
    .C(_07966_),
    .D(_07967_),
    .E(_07969_),
    .Y(_07970_));
 INVx1_ASAP7_75t_R _26200_ (.A(_07970_),
    .Y(_07971_));
 AND3x1_ASAP7_75t_R _26201_ (.A(_07071_),
    .B(_07066_),
    .C(_07678_),
    .Y(_07972_));
 OA21x2_ASAP7_75t_R _26202_ (.A1(_06982_),
    .A2(_07216_),
    .B(_07972_),
    .Y(_07973_));
 AND2x2_ASAP7_75t_R _26203_ (.A(_07071_),
    .B(_06928_),
    .Y(_07974_));
 AO21x1_ASAP7_75t_R _26204_ (.A1(_07583_),
    .A2(_07584_),
    .B(_06932_),
    .Y(_07975_));
 OA211x2_ASAP7_75t_R _26205_ (.A1(_06982_),
    .A2(_07588_),
    .B(_07974_),
    .C(_07975_),
    .Y(_07976_));
 OR5x1_ASAP7_75t_R _26206_ (.A(_07113_),
    .B(_07961_),
    .C(_07971_),
    .D(_07973_),
    .E(_07976_),
    .Y(_07977_));
 OR2x2_ASAP7_75t_R _26207_ (.A(net55),
    .B(net419),
    .Y(_07978_));
 OA21x2_ASAP7_75t_R _26208_ (.A1(net50),
    .A2(_07135_),
    .B(_07978_),
    .Y(_07979_));
 INVx1_ASAP7_75t_R _26209_ (.A(net32),
    .Y(_07980_));
 NAND2x1_ASAP7_75t_R _26210_ (.A(_07980_),
    .B(net419),
    .Y(_07981_));
 OAI21x1_ASAP7_75t_R _26211_ (.A1(net41),
    .A2(net419),
    .B(_07981_),
    .Y(_07982_));
 NAND2x1_ASAP7_75t_R _26212_ (.A(net418),
    .B(_07982_),
    .Y(_07983_));
 OA211x2_ASAP7_75t_R _26213_ (.A1(net418),
    .A2(_07979_),
    .B(_07983_),
    .C(_07727_),
    .Y(_07984_));
 INVx1_ASAP7_75t_R _26214_ (.A(_01849_),
    .Y(_07985_));
 OA211x2_ASAP7_75t_R _26215_ (.A1(_07135_),
    .A2(_07985_),
    .B(_07978_),
    .C(_07120_),
    .Y(_07986_));
 OA211x2_ASAP7_75t_R _26216_ (.A1(net419),
    .A2(_07613_),
    .B(_07981_),
    .C(net418),
    .Y(_07987_));
 OA21x2_ASAP7_75t_R _26217_ (.A1(_07986_),
    .A2(_07987_),
    .B(_07117_),
    .Y(_07988_));
 OR3x1_ASAP7_75t_R _26218_ (.A(_07736_),
    .B(_07984_),
    .C(_07988_),
    .Y(_07989_));
 OA21x2_ASAP7_75t_R _26219_ (.A1(_07953_),
    .A2(_07977_),
    .B(_07989_),
    .Y(_07990_));
 NOR2x1_ASAP7_75t_R _26220_ (.A(_01695_),
    .B(_06924_),
    .Y(_07991_));
 AO21x1_ASAP7_75t_R _26221_ (.A1(_06924_),
    .A2(_07990_),
    .B(_07991_),
    .Y(_02670_));
 AO211x2_ASAP7_75t_R _26222_ (.A1(_06935_),
    .A2(_07401_),
    .B(_07630_),
    .C(_06932_),
    .Y(_07992_));
 OA21x2_ASAP7_75t_R _26223_ (.A1(_06982_),
    .A2(_07636_),
    .B(_07992_),
    .Y(_07993_));
 OA21x2_ASAP7_75t_R _26224_ (.A1(_06982_),
    .A2(_07106_),
    .B(_07678_),
    .Y(_07994_));
 AND3x1_ASAP7_75t_R _26225_ (.A(_07071_),
    .B(_07066_),
    .C(_07994_),
    .Y(_07995_));
 INVx1_ASAP7_75t_R _26226_ (.A(_00112_),
    .Y(_07996_));
 NAND2x1_ASAP7_75t_R _26227_ (.A(_00113_),
    .B(_07202_),
    .Y(_07997_));
 OA211x2_ASAP7_75t_R _26228_ (.A1(_07996_),
    .A2(_07202_),
    .B(_07997_),
    .C(_07086_),
    .Y(_07998_));
 AO21x1_ASAP7_75t_R _26229_ (.A1(_02375_),
    .A2(net285),
    .B(_07998_),
    .Y(_07999_));
 AO22x1_ASAP7_75t_R _26230_ (.A1(net156),
    .A2(_07097_),
    .B1(_07999_),
    .B2(_07094_),
    .Y(_08000_));
 NAND2x1_ASAP7_75t_R _26231_ (.A(_00783_),
    .B(_07079_),
    .Y(_08001_));
 XOR2x2_ASAP7_75t_R _26232_ (.A(_00024_),
    .B(_02240_),
    .Y(_08002_));
 OR2x2_ASAP7_75t_R _26233_ (.A(_07079_),
    .B(_08002_),
    .Y(_08003_));
 AO21x1_ASAP7_75t_R _26234_ (.A1(_08001_),
    .A2(_08003_),
    .B(_05745_),
    .Y(_08004_));
 OA211x2_ASAP7_75t_R _26235_ (.A1(_00279_),
    .A2(_06789_),
    .B(_13313_),
    .C(_13317_),
    .Y(_08005_));
 AO22x1_ASAP7_75t_R _26236_ (.A1(net294),
    .A2(_08000_),
    .B1(_08004_),
    .B2(_08005_),
    .Y(_08006_));
 OAI22x1_ASAP7_75t_R _26237_ (.A1(_01504_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01473_),
    .Y(_08007_));
 NAND2x1_ASAP7_75t_R _26238_ (.A(_06884_),
    .B(_08007_),
    .Y(_08008_));
 OAI22x1_ASAP7_75t_R _26239_ (.A1(_02157_),
    .A2(net284),
    .B1(_07162_),
    .B2(_02051_),
    .Y(_08009_));
 NAND2x1_ASAP7_75t_R _26240_ (.A(_06886_),
    .B(_08009_),
    .Y(_08010_));
 NAND2x1_ASAP7_75t_R _26241_ (.A(net68),
    .B(_06891_),
    .Y(_08011_));
 OA211x2_ASAP7_75t_R _26242_ (.A1(_02014_),
    .A2(_07524_),
    .B(_08011_),
    .C(_07168_),
    .Y(_08012_));
 OR2x2_ASAP7_75t_R _26243_ (.A(_01980_),
    .B(_07511_),
    .Y(_08013_));
 OA22x2_ASAP7_75t_R _26244_ (.A1(_02030_),
    .A2(_07708_),
    .B1(_07508_),
    .B2(_02124_),
    .Y(_08014_));
 OA211x2_ASAP7_75t_R _26245_ (.A1(_01930_),
    .A2(_07701_),
    .B(_08013_),
    .C(_08014_),
    .Y(_08015_));
 OA222x2_ASAP7_75t_R _26246_ (.A1(_00114_),
    .A2(_07705_),
    .B1(_07516_),
    .B2(_01566_),
    .C1(_02083_),
    .C2(_07505_),
    .Y(_08016_));
 AND5x2_ASAP7_75t_R _26247_ (.A(_08008_),
    .B(_08010_),
    .C(_08012_),
    .D(_08015_),
    .E(_08016_),
    .Y(_08017_));
 INVx1_ASAP7_75t_R _26248_ (.A(_08017_),
    .Y(_08018_));
 OR4x1_ASAP7_75t_R _26249_ (.A(_07113_),
    .B(_07995_),
    .C(_08006_),
    .D(_08018_),
    .Y(_08019_));
 AO221x1_ASAP7_75t_R _26250_ (.A1(_07012_),
    .A2(_07348_),
    .B1(_07974_),
    .B2(_07993_),
    .C(_08019_),
    .Y(_08020_));
 OR2x2_ASAP7_75t_R _26251_ (.A(net33),
    .B(_07135_),
    .Y(_08021_));
 OA211x2_ASAP7_75t_R _26252_ (.A1(net42),
    .A2(net419),
    .B(_08021_),
    .C(net418),
    .Y(_08022_));
 INVx1_ASAP7_75t_R _26253_ (.A(_08022_),
    .Y(_08023_));
 NOR2x1_ASAP7_75t_R _26254_ (.A(net56),
    .B(net419),
    .Y(_08024_));
 AO21x1_ASAP7_75t_R _26255_ (.A1(_07626_),
    .A2(net419),
    .B(_08024_),
    .Y(_08025_));
 OR2x2_ASAP7_75t_R _26256_ (.A(net418),
    .B(_08025_),
    .Y(_08026_));
 AO21x1_ASAP7_75t_R _26257_ (.A1(_08023_),
    .A2(_08026_),
    .B(_01731_),
    .Y(_08027_));
 INVx1_ASAP7_75t_R _26258_ (.A(_08027_),
    .Y(_08028_));
 TAPCELL_ASAP7_75t_R TAP_710 ();
 AOI211x1_ASAP7_75t_R _26260_ (.A1(net419),
    .A2(_01733_),
    .B(_08024_),
    .C(net418),
    .Y(_08030_));
 OA211x2_ASAP7_75t_R _26261_ (.A1(net419),
    .A2(_07623_),
    .B(_08021_),
    .C(net418),
    .Y(_08031_));
 OA21x2_ASAP7_75t_R _26262_ (.A1(_08030_),
    .A2(_08031_),
    .B(_07117_),
    .Y(_08032_));
 OR3x1_ASAP7_75t_R _26263_ (.A(_07736_),
    .B(_08028_),
    .C(_08032_),
    .Y(_08033_));
 AND2x6_ASAP7_75t_R _26264_ (.A(_08020_),
    .B(_08033_),
    .Y(_08034_));
 NOR2x1_ASAP7_75t_R _26265_ (.A(_01694_),
    .B(_06924_),
    .Y(_08035_));
 AO21x1_ASAP7_75t_R _26266_ (.A1(_06924_),
    .A2(_08034_),
    .B(_08035_),
    .Y(_02671_));
 AO21x2_ASAP7_75t_R _26267_ (.A1(_07735_),
    .A2(_08027_),
    .B(_01644_),
    .Y(_08036_));
 NAND2x2_ASAP7_75t_R _26268_ (.A(_07113_),
    .B(_08036_),
    .Y(_08037_));
 AO21x1_ASAP7_75t_R _26269_ (.A1(net57),
    .A2(_07135_),
    .B(_07133_),
    .Y(_08038_));
 NAND2x1_ASAP7_75t_R _26270_ (.A(net34),
    .B(net420),
    .Y(_08039_));
 OA211x2_ASAP7_75t_R _26271_ (.A1(net420),
    .A2(_01855_),
    .B(_08039_),
    .C(_01642_),
    .Y(_08040_));
 INVx1_ASAP7_75t_R _26272_ (.A(_08040_),
    .Y(_08041_));
 OA211x2_ASAP7_75t_R _26273_ (.A1(_01642_),
    .A2(_08038_),
    .B(_08041_),
    .C(_07117_),
    .Y(_08042_));
 AND2x2_ASAP7_75t_R _26274_ (.A(_07066_),
    .B(_07994_),
    .Y(_08043_));
 AO21x1_ASAP7_75t_R _26275_ (.A1(_06928_),
    .A2(_07993_),
    .B(_08043_),
    .Y(_08044_));
 INVx1_ASAP7_75t_R _26276_ (.A(_00115_),
    .Y(_08045_));
 NAND2x1_ASAP7_75t_R _26277_ (.A(_00116_),
    .B(_07202_),
    .Y(_08046_));
 OA211x2_ASAP7_75t_R _26278_ (.A1(_08045_),
    .A2(_07202_),
    .B(_08046_),
    .C(_07086_),
    .Y(_08047_));
 AO21x1_ASAP7_75t_R _26279_ (.A1(_02376_),
    .A2(net285),
    .B(_08047_),
    .Y(_08048_));
 AO22x1_ASAP7_75t_R _26280_ (.A1(net157),
    .A2(_07097_),
    .B1(_08048_),
    .B2(_07094_),
    .Y(_08049_));
 AND2x2_ASAP7_75t_R _26281_ (.A(_01356_),
    .B(_07079_),
    .Y(_08050_));
 AO21x1_ASAP7_75t_R _26282_ (.A1(_00030_),
    .A2(_07077_),
    .B(_08050_),
    .Y(_08051_));
 AOI21x1_ASAP7_75t_R _26283_ (.A1(_07076_),
    .A2(_08051_),
    .B(_13318_),
    .Y(_08052_));
 NAND2x1_ASAP7_75t_R _26284_ (.A(_00816_),
    .B(_05743_),
    .Y(_08053_));
 AO22x1_ASAP7_75t_R _26285_ (.A1(net294),
    .A2(_08049_),
    .B1(_08052_),
    .B2(_08053_),
    .Y(_08054_));
 NOR2x1_ASAP7_75t_R _26286_ (.A(_02082_),
    .B(_07171_),
    .Y(_08055_));
 OAI21x1_ASAP7_75t_R _26287_ (.A1(_00117_),
    .A2(_07151_),
    .B(_07168_),
    .Y(_08056_));
 OAI22x1_ASAP7_75t_R _26288_ (.A1(_01979_),
    .A2(_07145_),
    .B1(_07305_),
    .B2(_01565_),
    .Y(_08057_));
 OAI22x1_ASAP7_75t_R _26289_ (.A1(_02013_),
    .A2(_07146_),
    .B1(_07149_),
    .B2(_01929_),
    .Y(_08058_));
 OR4x2_ASAP7_75t_R _26290_ (.A(_08055_),
    .B(_08056_),
    .C(_08057_),
    .D(_08058_),
    .Y(_08059_));
 AO21x1_ASAP7_75t_R _26291_ (.A1(net69),
    .A2(_07155_),
    .B(_08059_),
    .Y(_08060_));
 OAI22x1_ASAP7_75t_R _26292_ (.A1(_01503_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01472_),
    .Y(_08061_));
 AND2x2_ASAP7_75t_R _26293_ (.A(_06884_),
    .B(_08061_),
    .Y(_08062_));
 OAI22x1_ASAP7_75t_R _26294_ (.A1(_02156_),
    .A2(net284),
    .B1(_07162_),
    .B2(_02050_),
    .Y(_08063_));
 AND2x2_ASAP7_75t_R _26295_ (.A(_06886_),
    .B(_08063_),
    .Y(_08064_));
 AND3x1_ASAP7_75t_R _26296_ (.A(net130),
    .B(_05630_),
    .C(_06889_),
    .Y(_08065_));
 TAPCELL_ASAP7_75t_R TAP_709 ();
 OAI22x1_ASAP7_75t_R _26298_ (.A1(_02123_),
    .A2(_07299_),
    .B1(_07661_),
    .B2(_01963_),
    .Y(_08067_));
 OR5x2_ASAP7_75t_R _26299_ (.A(_08060_),
    .B(_08062_),
    .C(_08064_),
    .D(_08065_),
    .E(_08067_),
    .Y(_08068_));
 AND2x2_ASAP7_75t_R _26300_ (.A(_07066_),
    .B(_07101_),
    .Y(_08069_));
 OR2x2_ASAP7_75t_R _26301_ (.A(_07113_),
    .B(_08069_),
    .Y(_08070_));
 OR3x1_ASAP7_75t_R _26302_ (.A(_08054_),
    .B(_08068_),
    .C(_08070_),
    .Y(_08071_));
 AO221x1_ASAP7_75t_R _26303_ (.A1(_07012_),
    .A2(_07974_),
    .B1(_08044_),
    .B2(_06943_),
    .C(_08071_),
    .Y(_08072_));
 OA21x2_ASAP7_75t_R _26304_ (.A1(_08037_),
    .A2(_08042_),
    .B(_08072_),
    .Y(_08073_));
 NOR2x1_ASAP7_75t_R _26305_ (.A(_01693_),
    .B(_06924_),
    .Y(_08074_));
 AO21x1_ASAP7_75t_R _26306_ (.A1(_06924_),
    .A2(_08073_),
    .B(_08074_),
    .Y(_02672_));
 AND2x2_ASAP7_75t_R _26307_ (.A(_06982_),
    .B(_07101_),
    .Y(_08075_));
 AO21x1_ASAP7_75t_R _26308_ (.A1(_06932_),
    .A2(_07216_),
    .B(_08075_),
    .Y(_08076_));
 AO32x1_ASAP7_75t_R _26309_ (.A1(_07338_),
    .A2(_07583_),
    .A3(_07584_),
    .B1(_08076_),
    .B2(_07066_),
    .Y(_08077_));
 AND2x2_ASAP7_75t_R _26310_ (.A(_06943_),
    .B(_08077_),
    .Y(_08078_));
 OA211x2_ASAP7_75t_R _26311_ (.A1(_06982_),
    .A2(_07234_),
    .B(_07952_),
    .C(_07974_),
    .Y(_08079_));
 AND2x2_ASAP7_75t_R _26312_ (.A(_07588_),
    .B(_07641_),
    .Y(_08080_));
 INVx1_ASAP7_75t_R _26313_ (.A(_00118_),
    .Y(_08081_));
 NAND2x1_ASAP7_75t_R _26314_ (.A(_00119_),
    .B(_07202_),
    .Y(_08082_));
 OA211x2_ASAP7_75t_R _26315_ (.A1(_08081_),
    .A2(_07202_),
    .B(_08082_),
    .C(_07086_),
    .Y(_08083_));
 AO21x1_ASAP7_75t_R _26316_ (.A1(_02377_),
    .A2(net285),
    .B(_08083_),
    .Y(_08084_));
 AO22x1_ASAP7_75t_R _26317_ (.A1(net158),
    .A2(_07097_),
    .B1(_08084_),
    .B2(_07094_),
    .Y(_08085_));
 OR2x2_ASAP7_75t_R _26318_ (.A(_08069_),
    .B(_08085_),
    .Y(_08086_));
 XNOR2x1_ASAP7_75t_R _26319_ (.B(_00031_),
    .Y(_08087_),
    .A(_00033_));
 NOR2x1_ASAP7_75t_R _26320_ (.A(_01360_),
    .B(_07077_),
    .Y(_08088_));
 AO221x1_ASAP7_75t_R _26321_ (.A1(_13317_),
    .A2(_05743_),
    .B1(_07077_),
    .B2(_08087_),
    .C(_08088_),
    .Y(_08089_));
 NAND2x1_ASAP7_75t_R _26322_ (.A(_00849_),
    .B(_05743_),
    .Y(_08090_));
 AND3x1_ASAP7_75t_R _26323_ (.A(_13576_),
    .B(_08089_),
    .C(_08090_),
    .Y(_08091_));
 AO21x1_ASAP7_75t_R _26324_ (.A1(net294),
    .A2(_08086_),
    .B(_08091_),
    .Y(_08092_));
 OAI22x1_ASAP7_75t_R _26325_ (.A1(_02155_),
    .A2(net284),
    .B1(_07162_),
    .B2(_02049_),
    .Y(_08093_));
 NAND2x1_ASAP7_75t_R _26326_ (.A(_06886_),
    .B(_08093_),
    .Y(_08094_));
 OAI22x1_ASAP7_75t_R _26327_ (.A1(_01502_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01471_),
    .Y(_08095_));
 NAND2x1_ASAP7_75t_R _26328_ (.A(_06884_),
    .B(_08095_),
    .Y(_08096_));
 OA22x2_ASAP7_75t_R _26329_ (.A1(_02081_),
    .A2(_07505_),
    .B1(_07667_),
    .B2(_01996_),
    .Y(_08097_));
 OR2x2_ASAP7_75t_R _26330_ (.A(_07507_),
    .B(_07659_),
    .Y(_08098_));
 INVx1_ASAP7_75t_R _26331_ (.A(net136),
    .Y(_08099_));
 OA222x2_ASAP7_75t_R _26332_ (.A1(_00120_),
    .A2(_07705_),
    .B1(_07701_),
    .B2(_01928_),
    .C1(_08098_),
    .C2(_08099_),
    .Y(_08100_));
 OA22x2_ASAP7_75t_R _26333_ (.A1(_01978_),
    .A2(_07511_),
    .B1(_07524_),
    .B2(_02012_),
    .Y(_08101_));
 AND3x2_ASAP7_75t_R _26334_ (.A(_08097_),
    .B(_08100_),
    .C(_08101_),
    .Y(_08102_));
 OA22x2_ASAP7_75t_R _26335_ (.A1(_02122_),
    .A2(_07508_),
    .B1(_07661_),
    .B2(_01962_),
    .Y(_08103_));
 OA211x2_ASAP7_75t_R _26336_ (.A1(_01564_),
    .A2(_07516_),
    .B(_08103_),
    .C(_07168_),
    .Y(_08104_));
 NAND2x1_ASAP7_75t_R _26337_ (.A(net70),
    .B(_06891_),
    .Y(_08105_));
 AND5x2_ASAP7_75t_R _26338_ (.A(_08094_),
    .B(_08096_),
    .C(_08102_),
    .D(_08104_),
    .E(_08105_),
    .Y(_08106_));
 INVx1_ASAP7_75t_R _26339_ (.A(_08106_),
    .Y(_08107_));
 OR5x1_ASAP7_75t_R _26340_ (.A(_07113_),
    .B(_08079_),
    .C(_08080_),
    .D(_08092_),
    .E(_08107_),
    .Y(_08108_));
 AND2x6_ASAP7_75t_R _26341_ (.A(_07113_),
    .B(_08036_),
    .Y(_08109_));
 NAND2x1_ASAP7_75t_R _26342_ (.A(net38),
    .B(_01643_),
    .Y(_08110_));
 OA211x2_ASAP7_75t_R _26343_ (.A1(_07741_),
    .A2(_01643_),
    .B(_08110_),
    .C(_07120_),
    .Y(_08111_));
 NAND2x1_ASAP7_75t_R _26344_ (.A(net35),
    .B(_01643_),
    .Y(_08112_));
 OA211x2_ASAP7_75t_R _26345_ (.A1(_01643_),
    .A2(_01854_),
    .B(_08112_),
    .C(_01642_),
    .Y(_08113_));
 OR3x1_ASAP7_75t_R _26346_ (.A(_07115_),
    .B(_08111_),
    .C(_08113_),
    .Y(_08114_));
 NAND2x1_ASAP7_75t_R _26347_ (.A(_08109_),
    .B(_08114_),
    .Y(_08115_));
 OA21x2_ASAP7_75t_R _26348_ (.A1(_08078_),
    .A2(_08108_),
    .B(_08115_),
    .Y(_08116_));
 NOR2x1_ASAP7_75t_R _26349_ (.A(_01692_),
    .B(_06924_),
    .Y(_08117_));
 AO21x1_ASAP7_75t_R _26350_ (.A1(_06924_),
    .A2(_08116_),
    .B(_08117_),
    .Y(_02673_));
 TAPCELL_ASAP7_75t_R TAP_708 ();
 NOR2x1_ASAP7_75t_R _26352_ (.A(_02243_),
    .B(_07079_),
    .Y(_08119_));
 AO21x1_ASAP7_75t_R _26353_ (.A1(_01364_),
    .A2(_07079_),
    .B(_08119_),
    .Y(_08120_));
 AO21x1_ASAP7_75t_R _26354_ (.A1(_07076_),
    .A2(_08120_),
    .B(_13318_),
    .Y(_08121_));
 AO21x1_ASAP7_75t_R _26355_ (.A1(_00881_),
    .A2(_05743_),
    .B(_08121_),
    .Y(_08122_));
 OA222x2_ASAP7_75t_R _26356_ (.A1(_00123_),
    .A2(_07705_),
    .B1(_07701_),
    .B2(_01927_),
    .C1(_02080_),
    .C2(_07505_),
    .Y(_08123_));
 OA21x2_ASAP7_75t_R _26357_ (.A1(_01563_),
    .A2(_07516_),
    .B(_08123_),
    .Y(_08124_));
 NAND2x1_ASAP7_75t_R _26358_ (.A(net71),
    .B(_06891_),
    .Y(_08125_));
 OA211x2_ASAP7_75t_R _26359_ (.A1(_02121_),
    .A2(_07508_),
    .B(_08125_),
    .C(_07168_),
    .Y(_08126_));
 OA22x2_ASAP7_75t_R _26360_ (.A1(_01977_),
    .A2(_07511_),
    .B1(_07661_),
    .B2(_01961_),
    .Y(_08127_));
 NAND2x1_ASAP7_75t_R _26361_ (.A(net137),
    .B(_07841_),
    .Y(_08128_));
 OA211x2_ASAP7_75t_R _26362_ (.A1(_02011_),
    .A2(_07524_),
    .B(_08127_),
    .C(_08128_),
    .Y(_08129_));
 OAI22x1_ASAP7_75t_R _26363_ (.A1(_01501_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01470_),
    .Y(_08130_));
 OAI22x1_ASAP7_75t_R _26364_ (.A1(_02154_),
    .A2(net283),
    .B1(net282),
    .B2(_02048_),
    .Y(_08131_));
 AOI22x1_ASAP7_75t_R _26365_ (.A1(_06884_),
    .A2(_08130_),
    .B1(_08131_),
    .B2(_06886_),
    .Y(_08132_));
 AND4x2_ASAP7_75t_R _26366_ (.A(_08124_),
    .B(_08126_),
    .C(_08129_),
    .D(_08132_),
    .Y(_08133_));
 NAND2x1_ASAP7_75t_R _26367_ (.A(_06943_),
    .B(_07936_),
    .Y(_08134_));
 AND4x1_ASAP7_75t_R _26368_ (.A(_06920_),
    .B(_08122_),
    .C(_08133_),
    .D(_08134_),
    .Y(_08135_));
 INVx1_ASAP7_75t_R _26369_ (.A(_00121_),
    .Y(_08136_));
 NAND2x1_ASAP7_75t_R _26370_ (.A(_00122_),
    .B(_07202_),
    .Y(_08137_));
 OA211x2_ASAP7_75t_R _26371_ (.A1(_08136_),
    .A2(_07202_),
    .B(_08137_),
    .C(_07086_),
    .Y(_08138_));
 AO21x1_ASAP7_75t_R _26372_ (.A1(_02378_),
    .A2(net285),
    .B(_08138_),
    .Y(_08139_));
 AOI22x1_ASAP7_75t_R _26373_ (.A1(net159),
    .A2(_07097_),
    .B1(_08139_),
    .B2(_07094_),
    .Y(_08140_));
 OA21x2_ASAP7_75t_R _26374_ (.A1(_06928_),
    .A2(_07214_),
    .B(_07071_),
    .Y(_08141_));
 OAI21x1_ASAP7_75t_R _26375_ (.A1(_07066_),
    .A2(_07331_),
    .B(_08141_),
    .Y(_08142_));
 AO21x1_ASAP7_75t_R _26376_ (.A1(_08140_),
    .A2(_08142_),
    .B(_13576_),
    .Y(_08143_));
 AND2x2_ASAP7_75t_R _26377_ (.A(net49),
    .B(net419),
    .Y(_08144_));
 AO21x1_ASAP7_75t_R _26378_ (.A1(net28),
    .A2(_07135_),
    .B(_08144_),
    .Y(_08145_));
 NAND2x1_ASAP7_75t_R _26379_ (.A(_07135_),
    .B(_01853_),
    .Y(_08146_));
 OA211x2_ASAP7_75t_R _26380_ (.A1(net36),
    .A2(_07135_),
    .B(_08146_),
    .C(net418),
    .Y(_08147_));
 AO21x1_ASAP7_75t_R _26381_ (.A1(_07120_),
    .A2(_08145_),
    .B(_08147_),
    .Y(_08148_));
 AOI21x1_ASAP7_75t_R _26382_ (.A1(_07117_),
    .A2(_08148_),
    .B(_08037_),
    .Y(_08149_));
 AOI21x1_ASAP7_75t_R _26383_ (.A1(_08135_),
    .A2(_08143_),
    .B(_08149_),
    .Y(_08150_));
 TAPCELL_ASAP7_75t_R TAP_707 ();
 NOR2x1_ASAP7_75t_R _26385_ (.A(_01691_),
    .B(_06924_),
    .Y(_08152_));
 AO21x1_ASAP7_75t_R _26386_ (.A1(_06924_),
    .A2(_08150_),
    .B(_08152_),
    .Y(_02674_));
 AND2x2_ASAP7_75t_R _26387_ (.A(_06943_),
    .B(_07870_),
    .Y(_08153_));
 NOR3x1_ASAP7_75t_R _26388_ (.A(_07544_),
    .B(_07066_),
    .C(_07410_),
    .Y(_08154_));
 INVx1_ASAP7_75t_R _26389_ (.A(_00124_),
    .Y(_08155_));
 NAND2x1_ASAP7_75t_R _26390_ (.A(_00125_),
    .B(_07202_),
    .Y(_08156_));
 OA211x2_ASAP7_75t_R _26391_ (.A1(_08155_),
    .A2(_07202_),
    .B(_08156_),
    .C(_07086_),
    .Y(_08157_));
 AO21x1_ASAP7_75t_R _26392_ (.A1(_02379_),
    .A2(net285),
    .B(_08157_),
    .Y(_08158_));
 AO22x1_ASAP7_75t_R _26393_ (.A1(net257),
    .A2(_07097_),
    .B1(_08158_),
    .B2(_07094_),
    .Y(_08159_));
 OR2x2_ASAP7_75t_R _26394_ (.A(_02231_),
    .B(_07077_),
    .Y(_08160_));
 XNOR2x1_ASAP7_75t_R _26395_ (.B(_02242_),
    .Y(_08161_),
    .A(_00038_));
 NAND2x1_ASAP7_75t_R _26396_ (.A(_07077_),
    .B(_08161_),
    .Y(_08162_));
 AO21x1_ASAP7_75t_R _26397_ (.A1(_08160_),
    .A2(_08162_),
    .B(_05745_),
    .Y(_08163_));
 NAND2x1_ASAP7_75t_R _26398_ (.A(_00914_),
    .B(_05743_),
    .Y(_08164_));
 AND3x1_ASAP7_75t_R _26399_ (.A(_13576_),
    .B(_08163_),
    .C(_08164_),
    .Y(_08165_));
 AO21x1_ASAP7_75t_R _26400_ (.A1(net294),
    .A2(_08159_),
    .B(_08165_),
    .Y(_08166_));
 OAI22x1_ASAP7_75t_R _26401_ (.A1(_02153_),
    .A2(net283),
    .B1(net282),
    .B2(_02047_),
    .Y(_08167_));
 NAND2x1_ASAP7_75t_R _26402_ (.A(_06886_),
    .B(_08167_),
    .Y(_08168_));
 OAI22x1_ASAP7_75t_R _26403_ (.A1(_01500_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01469_),
    .Y(_08169_));
 NAND2x1_ASAP7_75t_R _26404_ (.A(_06884_),
    .B(_08169_),
    .Y(_08170_));
 NAND2x1_ASAP7_75t_R _26405_ (.A(net72),
    .B(_06891_),
    .Y(_08171_));
 OA211x2_ASAP7_75t_R _26406_ (.A1(_01976_),
    .A2(_07511_),
    .B(_08171_),
    .C(_07168_),
    .Y(_08172_));
 OA222x2_ASAP7_75t_R _26407_ (.A1(_01926_),
    .A2(_07701_),
    .B1(_07524_),
    .B2(_02010_),
    .C1(_02079_),
    .C2(_07505_),
    .Y(_08173_));
 OA211x2_ASAP7_75t_R _26408_ (.A1(_01960_),
    .A2(_07661_),
    .B(_08172_),
    .C(_08173_),
    .Y(_08174_));
 OA22x2_ASAP7_75t_R _26409_ (.A1(_00126_),
    .A2(_07705_),
    .B1(_07516_),
    .B2(_01562_),
    .Y(_08175_));
 NAND2x1_ASAP7_75t_R _26410_ (.A(net138),
    .B(_07841_),
    .Y(_08176_));
 OA211x2_ASAP7_75t_R _26411_ (.A1(_02120_),
    .A2(_07508_),
    .B(_08175_),
    .C(_08176_),
    .Y(_08177_));
 AND4x2_ASAP7_75t_R _26412_ (.A(_08168_),
    .B(_08170_),
    .C(_08174_),
    .D(_08177_),
    .Y(_08178_));
 INVx1_ASAP7_75t_R _26413_ (.A(_08178_),
    .Y(_08179_));
 OR4x1_ASAP7_75t_R _26414_ (.A(_08070_),
    .B(_08154_),
    .C(_08166_),
    .D(_08179_),
    .Y(_08180_));
 NAND2x1_ASAP7_75t_R _26415_ (.A(net52),
    .B(net420),
    .Y(_08181_));
 OA211x2_ASAP7_75t_R _26416_ (.A1(_07854_),
    .A2(net420),
    .B(_08181_),
    .C(_07120_),
    .Y(_08182_));
 NAND2x1_ASAP7_75t_R _26417_ (.A(net37),
    .B(net420),
    .Y(_08183_));
 OA211x2_ASAP7_75t_R _26418_ (.A1(net420),
    .A2(_01852_),
    .B(_08183_),
    .C(_01642_),
    .Y(_08184_));
 OR3x1_ASAP7_75t_R _26419_ (.A(_07115_),
    .B(_08182_),
    .C(_08184_),
    .Y(_08185_));
 NAND2x1_ASAP7_75t_R _26420_ (.A(_08109_),
    .B(_08185_),
    .Y(_08186_));
 OA21x2_ASAP7_75t_R _26421_ (.A1(_08153_),
    .A2(_08180_),
    .B(_08186_),
    .Y(_08187_));
 NOR2x1_ASAP7_75t_R _26422_ (.A(_01690_),
    .B(_06924_),
    .Y(_08188_));
 AO21x1_ASAP7_75t_R _26423_ (.A1(_06924_),
    .A2(_08187_),
    .B(_08188_),
    .Y(_02675_));
 TAPCELL_ASAP7_75t_R TAP_706 ();
 AND2x2_ASAP7_75t_R _26425_ (.A(net53),
    .B(net419),
    .Y(_08190_));
 AO21x1_ASAP7_75t_R _26426_ (.A1(net30),
    .A2(_07135_),
    .B(_08190_),
    .Y(_08191_));
 NAND2x1_ASAP7_75t_R _26427_ (.A(net39),
    .B(net419),
    .Y(_08192_));
 OA211x2_ASAP7_75t_R _26428_ (.A1(net419),
    .A2(_01851_),
    .B(_08192_),
    .C(net418),
    .Y(_08193_));
 INVx1_ASAP7_75t_R _26429_ (.A(_08193_),
    .Y(_08194_));
 OA211x2_ASAP7_75t_R _26430_ (.A1(net418),
    .A2(_08191_),
    .B(_08194_),
    .C(_07117_),
    .Y(_08195_));
 INVx1_ASAP7_75t_R _26431_ (.A(_00127_),
    .Y(_08196_));
 NAND2x1_ASAP7_75t_R _26432_ (.A(_00128_),
    .B(_07202_),
    .Y(_08197_));
 OA211x2_ASAP7_75t_R _26433_ (.A1(_08196_),
    .A2(_07202_),
    .B(_08197_),
    .C(_07086_),
    .Y(_08198_));
 AO21x1_ASAP7_75t_R _26434_ (.A1(_02380_),
    .A2(net285),
    .B(_08198_),
    .Y(_08199_));
 AO22x1_ASAP7_75t_R _26435_ (.A1(net161),
    .A2(_07097_),
    .B1(_08199_),
    .B2(_07094_),
    .Y(_08200_));
 NOR2x1_ASAP7_75t_R _26436_ (.A(_01376_),
    .B(_07077_),
    .Y(_08201_));
 AO21x1_ASAP7_75t_R _26437_ (.A1(_02245_),
    .A2(_07077_),
    .B(_08201_),
    .Y(_08202_));
 OA21x2_ASAP7_75t_R _26438_ (.A1(_05745_),
    .A2(_08202_),
    .B(_13576_),
    .Y(_08203_));
 NAND2x1_ASAP7_75t_R _26439_ (.A(_00946_),
    .B(_05743_),
    .Y(_08204_));
 AO22x1_ASAP7_75t_R _26440_ (.A1(net295),
    .A2(_08200_),
    .B1(_08203_),
    .B2(_08204_),
    .Y(_08205_));
 OAI22x1_ASAP7_75t_R _26441_ (.A1(_01499_),
    .A2(net283),
    .B1(net282),
    .B2(_01468_),
    .Y(_08206_));
 NAND2x1_ASAP7_75t_R _26442_ (.A(_06884_),
    .B(_08206_),
    .Y(_08207_));
 OAI22x1_ASAP7_75t_R _26443_ (.A1(_02152_),
    .A2(net283),
    .B1(net282),
    .B2(_02046_),
    .Y(_08208_));
 NAND2x1_ASAP7_75t_R _26444_ (.A(_06886_),
    .B(_08208_),
    .Y(_08209_));
 OA222x2_ASAP7_75t_R _26445_ (.A1(_02078_),
    .A2(_07171_),
    .B1(_07661_),
    .B2(_01959_),
    .C1(_06239_),
    .C2(_07663_),
    .Y(_08210_));
 AND3x1_ASAP7_75t_R _26446_ (.A(_08207_),
    .B(_08209_),
    .C(_08210_),
    .Y(_08211_));
 AOI21x1_ASAP7_75t_R _26447_ (.A1(net74),
    .A2(_07155_),
    .B(_07699_),
    .Y(_08212_));
 OA222x2_ASAP7_75t_R _26448_ (.A1(_01925_),
    .A2(_07149_),
    .B1(_07299_),
    .B2(_02119_),
    .C1(_07305_),
    .C2(_01561_),
    .Y(_08213_));
 OA222x2_ASAP7_75t_R _26449_ (.A1(_01975_),
    .A2(_07145_),
    .B1(_07146_),
    .B2(_02009_),
    .C1(_07151_),
    .C2(_00129_),
    .Y(_08214_));
 AND4x2_ASAP7_75t_R _26450_ (.A(_08211_),
    .B(_08212_),
    .C(_08213_),
    .D(_08214_),
    .Y(_08215_));
 INVx1_ASAP7_75t_R _26451_ (.A(_08215_),
    .Y(_08216_));
 OR3x2_ASAP7_75t_R _26452_ (.A(_08070_),
    .B(_08205_),
    .C(_08216_),
    .Y(_08217_));
 AO221x1_ASAP7_75t_R _26453_ (.A1(_06943_),
    .A2(_07823_),
    .B1(_08141_),
    .B2(_07819_),
    .C(_08217_),
    .Y(_08218_));
 OA21x2_ASAP7_75t_R _26454_ (.A1(_08037_),
    .A2(_08195_),
    .B(_08218_),
    .Y(_08219_));
 NOR2x1_ASAP7_75t_R _26455_ (.A(_01689_),
    .B(_06924_),
    .Y(_08220_));
 AO21x1_ASAP7_75t_R _26456_ (.A1(_06924_),
    .A2(_08219_),
    .B(_08220_),
    .Y(_02676_));
 OA21x2_ASAP7_75t_R _26457_ (.A1(_07066_),
    .A2(_07550_),
    .B(_08141_),
    .Y(_08221_));
 INVx1_ASAP7_75t_R _26458_ (.A(_00130_),
    .Y(_08222_));
 NAND2x1_ASAP7_75t_R _26459_ (.A(_00131_),
    .B(_07202_),
    .Y(_08223_));
 OA211x2_ASAP7_75t_R _26460_ (.A1(_08222_),
    .A2(_07202_),
    .B(_08223_),
    .C(_07086_),
    .Y(_08224_));
 AO21x1_ASAP7_75t_R _26461_ (.A1(_02381_),
    .A2(net285),
    .B(_08224_),
    .Y(_08225_));
 AOI22x1_ASAP7_75t_R _26462_ (.A1(net255),
    .A2(_07097_),
    .B1(_08225_),
    .B2(_07094_),
    .Y(_08226_));
 XOR2x1_ASAP7_75t_R _26463_ (.A(_00044_),
    .Y(_08227_),
    .B(_02244_));
 NAND2x1_ASAP7_75t_R _26464_ (.A(_07079_),
    .B(_07561_),
    .Y(_08228_));
 OA21x2_ASAP7_75t_R _26465_ (.A1(_07079_),
    .A2(_08227_),
    .B(_08228_),
    .Y(_08229_));
 OA21x2_ASAP7_75t_R _26466_ (.A1(_05745_),
    .A2(_08229_),
    .B(_13576_),
    .Y(_08230_));
 INVx1_ASAP7_75t_R _26467_ (.A(_08230_),
    .Y(_08231_));
 AO21x1_ASAP7_75t_R _26468_ (.A1(_00979_),
    .A2(_05743_),
    .B(_08231_),
    .Y(_08232_));
 OAI22x1_ASAP7_75t_R _26469_ (.A1(_02151_),
    .A2(net283),
    .B1(net282),
    .B2(_02045_),
    .Y(_08233_));
 NAND2x1_ASAP7_75t_R _26470_ (.A(_06886_),
    .B(_08233_),
    .Y(_08234_));
 OAI22x1_ASAP7_75t_R _26471_ (.A1(_01498_),
    .A2(net284),
    .B1(_07162_),
    .B2(_01467_),
    .Y(_08235_));
 NAND2x1_ASAP7_75t_R _26472_ (.A(_06884_),
    .B(_08235_),
    .Y(_08236_));
 INVx1_ASAP7_75t_R _26473_ (.A(net140),
    .Y(_08237_));
 OA222x2_ASAP7_75t_R _26474_ (.A1(_00132_),
    .A2(_07705_),
    .B1(_07516_),
    .B2(_01560_),
    .C1(_08098_),
    .C2(_08237_),
    .Y(_08238_));
 OA222x2_ASAP7_75t_R _26475_ (.A1(_01924_),
    .A2(_07701_),
    .B1(_07661_),
    .B2(_01958_),
    .C1(_02077_),
    .C2(_07505_),
    .Y(_08239_));
 OA211x2_ASAP7_75t_R _26476_ (.A1(_02118_),
    .A2(_07508_),
    .B(_08238_),
    .C(_08239_),
    .Y(_08240_));
 OA22x2_ASAP7_75t_R _26477_ (.A1(_02008_),
    .A2(_07524_),
    .B1(_07667_),
    .B2(_01997_),
    .Y(_08241_));
 OA211x2_ASAP7_75t_R _26478_ (.A1(_01974_),
    .A2(_07511_),
    .B(_08241_),
    .C(_07168_),
    .Y(_08242_));
 NAND2x1_ASAP7_75t_R _26479_ (.A(net75),
    .B(_06891_),
    .Y(_08243_));
 AND5x2_ASAP7_75t_R _26480_ (.A(_08234_),
    .B(_08236_),
    .C(_08240_),
    .D(_08242_),
    .E(_08243_),
    .Y(_08244_));
 OA211x2_ASAP7_75t_R _26481_ (.A1(_13576_),
    .A2(_08226_),
    .B(_08232_),
    .C(_08244_),
    .Y(_08245_));
 NAND2x1_ASAP7_75t_R _26482_ (.A(_06920_),
    .B(_08245_),
    .Y(_08246_));
 AND2x2_ASAP7_75t_R _26483_ (.A(_06943_),
    .B(_07784_),
    .Y(_08247_));
 NAND2x1_ASAP7_75t_R _26484_ (.A(net54),
    .B(net420),
    .Y(_08248_));
 OA211x2_ASAP7_75t_R _26485_ (.A1(_07940_),
    .A2(net420),
    .B(_08248_),
    .C(_07120_),
    .Y(_08249_));
 NAND2x1_ASAP7_75t_R _26486_ (.A(net40),
    .B(net420),
    .Y(_08250_));
 OA211x2_ASAP7_75t_R _26487_ (.A1(net420),
    .A2(_01850_),
    .B(_08250_),
    .C(_01642_),
    .Y(_08251_));
 OR3x1_ASAP7_75t_R _26488_ (.A(_07115_),
    .B(_08249_),
    .C(_08251_),
    .Y(_08252_));
 NAND2x1_ASAP7_75t_R _26489_ (.A(_08109_),
    .B(_08252_),
    .Y(_08253_));
 OA31x2_ASAP7_75t_R _26490_ (.A1(_08221_),
    .A2(_08246_),
    .A3(_08247_),
    .B1(_08253_),
    .Y(_08254_));
 NOR2x1_ASAP7_75t_R _26491_ (.A(_01688_),
    .B(_06924_),
    .Y(_08255_));
 AO21x1_ASAP7_75t_R _26492_ (.A1(_06924_),
    .A2(_08254_),
    .B(_08255_),
    .Y(_02677_));
 NAND2x1_ASAP7_75t_R _26493_ (.A(net41),
    .B(net419),
    .Y(_08256_));
 OA211x2_ASAP7_75t_R _26494_ (.A1(net419),
    .A2(_01849_),
    .B(_08256_),
    .C(net418),
    .Y(_08257_));
 NAND2x1_ASAP7_75t_R _26495_ (.A(net55),
    .B(net419),
    .Y(_08258_));
 OA211x2_ASAP7_75t_R _26496_ (.A1(_07980_),
    .A2(net419),
    .B(_08258_),
    .C(_07120_),
    .Y(_08259_));
 OR3x1_ASAP7_75t_R _26497_ (.A(_07115_),
    .B(_08257_),
    .C(_08259_),
    .Y(_08260_));
 AO21x1_ASAP7_75t_R _26498_ (.A1(_07755_),
    .A2(_07757_),
    .B(_06946_),
    .Y(_08261_));
 OAI22x1_ASAP7_75t_R _26499_ (.A1(_02150_),
    .A2(net283),
    .B1(net282),
    .B2(_02044_),
    .Y(_08262_));
 NAND2x1_ASAP7_75t_R _26500_ (.A(_06886_),
    .B(_08262_),
    .Y(_08263_));
 OAI22x1_ASAP7_75t_R _26501_ (.A1(_01497_),
    .A2(net283),
    .B1(net282),
    .B2(_01466_),
    .Y(_08264_));
 NAND2x1_ASAP7_75t_R _26502_ (.A(_06884_),
    .B(_08264_),
    .Y(_08265_));
 INVx1_ASAP7_75t_R _26503_ (.A(net141),
    .Y(_08266_));
 OA222x2_ASAP7_75t_R _26504_ (.A1(_02076_),
    .A2(_07171_),
    .B1(_07299_),
    .B2(_02117_),
    .C1(_07663_),
    .C2(_08266_),
    .Y(_08267_));
 OA222x2_ASAP7_75t_R _26505_ (.A1(_01923_),
    .A2(_07149_),
    .B1(_07661_),
    .B2(_01957_),
    .C1(_05684_),
    .C2(_06908_),
    .Y(_08268_));
 OA22x2_ASAP7_75t_R _26506_ (.A1(_00135_),
    .A2(_07151_),
    .B1(_07305_),
    .B2(_01559_),
    .Y(_08269_));
 OA22x2_ASAP7_75t_R _26507_ (.A1(_01973_),
    .A2(_07145_),
    .B1(_07146_),
    .B2(_02007_),
    .Y(_08270_));
 NAND2x1_ASAP7_75t_R _26508_ (.A(net76),
    .B(_07155_),
    .Y(_08271_));
 AND4x2_ASAP7_75t_R _26509_ (.A(_08268_),
    .B(_08269_),
    .C(_08270_),
    .D(_08271_),
    .Y(_08272_));
 AND4x2_ASAP7_75t_R _26510_ (.A(_08263_),
    .B(_08265_),
    .C(_08267_),
    .D(_08272_),
    .Y(_08273_));
 INVx1_ASAP7_75t_R _26511_ (.A(_00133_),
    .Y(_08274_));
 NAND2x1_ASAP7_75t_R _26512_ (.A(_00134_),
    .B(_07202_),
    .Y(_08275_));
 OA211x2_ASAP7_75t_R _26513_ (.A1(_08274_),
    .A2(_07202_),
    .B(_08275_),
    .C(_07086_),
    .Y(_08276_));
 AO21x1_ASAP7_75t_R _26514_ (.A1(_02382_),
    .A2(net285),
    .B(_08276_),
    .Y(_08277_));
 AO22x1_ASAP7_75t_R _26515_ (.A1(net163),
    .A2(_07097_),
    .B1(_08277_),
    .B2(_07094_),
    .Y(_08278_));
 AND2x2_ASAP7_75t_R _26516_ (.A(_02233_),
    .B(_07079_),
    .Y(_08279_));
 AO21x2_ASAP7_75t_R _26517_ (.A1(_02247_),
    .A2(_07077_),
    .B(_08279_),
    .Y(_08280_));
 NAND2x1_ASAP7_75t_R _26518_ (.A(_01011_),
    .B(_05743_),
    .Y(_08281_));
 OA211x2_ASAP7_75t_R _26519_ (.A1(_05745_),
    .A2(_08280_),
    .B(_08281_),
    .C(_13576_),
    .Y(_08282_));
 AO21x2_ASAP7_75t_R _26520_ (.A1(net295),
    .A2(_08278_),
    .B(_08282_),
    .Y(_08283_));
 NOR2x2_ASAP7_75t_R _26521_ (.A(_08069_),
    .B(_08283_),
    .Y(_08284_));
 NAND2x1_ASAP7_75t_R _26522_ (.A(_07586_),
    .B(_07974_),
    .Y(_08285_));
 AND5x2_ASAP7_75t_R _26523_ (.A(_06920_),
    .B(_08261_),
    .C(_08273_),
    .D(_08284_),
    .E(_08285_),
    .Y(_08286_));
 AOI21x1_ASAP7_75t_R _26524_ (.A1(_08109_),
    .A2(_08260_),
    .B(_08286_),
    .Y(_08287_));
 NOR2x1_ASAP7_75t_R _26525_ (.A(_01687_),
    .B(_06924_),
    .Y(_08288_));
 AO21x1_ASAP7_75t_R _26526_ (.A1(_06924_),
    .A2(_08287_),
    .B(_08288_),
    .Y(_02678_));
 OA211x2_ASAP7_75t_R _26527_ (.A1(net420),
    .A2(_01733_),
    .B(_07732_),
    .C(net418),
    .Y(_08289_));
 INVx1_ASAP7_75t_R _26528_ (.A(_08289_),
    .Y(_08290_));
 OA211x2_ASAP7_75t_R _26529_ (.A1(_01642_),
    .A2(_07730_),
    .B(_08290_),
    .C(_07117_),
    .Y(_08291_));
 NOR2x1_ASAP7_75t_R _26530_ (.A(_06946_),
    .B(_07683_),
    .Y(_08292_));
 INVx1_ASAP7_75t_R _26531_ (.A(_00136_),
    .Y(_08293_));
 NAND2x1_ASAP7_75t_R _26532_ (.A(_00137_),
    .B(_07202_),
    .Y(_08294_));
 OA211x2_ASAP7_75t_R _26533_ (.A1(_08293_),
    .A2(_07202_),
    .B(_08294_),
    .C(_07086_),
    .Y(_08295_));
 AO21x1_ASAP7_75t_R _26534_ (.A1(_02383_),
    .A2(net285),
    .B(_08295_),
    .Y(_08296_));
 AO22x1_ASAP7_75t_R _26535_ (.A1(net164),
    .A2(_07097_),
    .B1(_08296_),
    .B2(_07094_),
    .Y(_08297_));
 NAND2x1_ASAP7_75t_R _26536_ (.A(_01045_),
    .B(_05743_),
    .Y(_08298_));
 XNOR2x1_ASAP7_75t_R _26537_ (.B(_02246_),
    .Y(_08299_),
    .A(_00052_));
 NAND2x1_ASAP7_75t_R _26538_ (.A(_07077_),
    .B(_08299_),
    .Y(_08300_));
 OA21x2_ASAP7_75t_R _26539_ (.A1(_07077_),
    .A2(_07650_),
    .B(_08300_),
    .Y(_08301_));
 OA21x2_ASAP7_75t_R _26540_ (.A1(_05745_),
    .A2(_08301_),
    .B(_13576_),
    .Y(_08302_));
 AO22x1_ASAP7_75t_R _26541_ (.A1(net295),
    .A2(_08297_),
    .B1(_08298_),
    .B2(_08302_),
    .Y(_08303_));
 OA222x2_ASAP7_75t_R _26542_ (.A1(_00138_),
    .A2(_07151_),
    .B1(_07171_),
    .B2(_02075_),
    .C1(_05684_),
    .C2(_06908_),
    .Y(_08304_));
 OA22x2_ASAP7_75t_R _26543_ (.A1(_01972_),
    .A2(_07145_),
    .B1(_07305_),
    .B2(_01558_),
    .Y(_08305_));
 OA22x2_ASAP7_75t_R _26544_ (.A1(_02006_),
    .A2(_07146_),
    .B1(_07149_),
    .B2(_01922_),
    .Y(_08306_));
 NAND2x1_ASAP7_75t_R _26545_ (.A(net77),
    .B(_07155_),
    .Y(_08307_));
 AND4x2_ASAP7_75t_R _26546_ (.A(_08304_),
    .B(_08305_),
    .C(_08306_),
    .D(_08307_),
    .Y(_08308_));
 OAI22x1_ASAP7_75t_R _26547_ (.A1(_01496_),
    .A2(net283),
    .B1(net282),
    .B2(_01465_),
    .Y(_08309_));
 NAND2x1_ASAP7_75t_R _26548_ (.A(_06884_),
    .B(_08309_),
    .Y(_08310_));
 OAI22x1_ASAP7_75t_R _26549_ (.A1(_02149_),
    .A2(net283),
    .B1(net282),
    .B2(_02043_),
    .Y(_08311_));
 NAND2x1_ASAP7_75t_R _26550_ (.A(_06886_),
    .B(_08311_),
    .Y(_08312_));
 INVx1_ASAP7_75t_R _26551_ (.A(net142),
    .Y(_08313_));
 OA222x2_ASAP7_75t_R _26552_ (.A1(_02116_),
    .A2(_07299_),
    .B1(_07661_),
    .B2(_01956_),
    .C1(_08313_),
    .C2(_07663_),
    .Y(_08314_));
 AND4x2_ASAP7_75t_R _26553_ (.A(_08308_),
    .B(_08310_),
    .C(_08312_),
    .D(_08314_),
    .Y(_08315_));
 INVx1_ASAP7_75t_R _26554_ (.A(_08315_),
    .Y(_08316_));
 OA21x2_ASAP7_75t_R _26555_ (.A1(_07066_),
    .A2(_07633_),
    .B(_08141_),
    .Y(_08317_));
 OR4x2_ASAP7_75t_R _26556_ (.A(_07113_),
    .B(_08303_),
    .C(_08316_),
    .D(_08317_),
    .Y(_08318_));
 OA22x2_ASAP7_75t_R _26557_ (.A1(_08037_),
    .A2(_08291_),
    .B1(_08292_),
    .B2(_08318_),
    .Y(_08319_));
 NOR2x1_ASAP7_75t_R _26558_ (.A(_01686_),
    .B(_06924_),
    .Y(_08320_));
 AO21x1_ASAP7_75t_R _26559_ (.A1(_06924_),
    .A2(_08319_),
    .B(_08320_),
    .Y(_02679_));
 NAND2x1_ASAP7_75t_R _26560_ (.A(_01642_),
    .B(_07723_),
    .Y(_08321_));
 OR2x2_ASAP7_75t_R _26561_ (.A(_01642_),
    .B(_07725_),
    .Y(_08322_));
 AO21x1_ASAP7_75t_R _26562_ (.A1(_08321_),
    .A2(_08322_),
    .B(_07115_),
    .Y(_08323_));
 NAND2x1_ASAP7_75t_R _26563_ (.A(_06943_),
    .B(_07638_),
    .Y(_08324_));
 OA21x2_ASAP7_75t_R _26564_ (.A1(_07107_),
    .A2(_07101_),
    .B(_07071_),
    .Y(_08325_));
 INVx1_ASAP7_75t_R _26565_ (.A(_00139_),
    .Y(_08326_));
 NAND2x1_ASAP7_75t_R _26566_ (.A(_00140_),
    .B(_07202_),
    .Y(_08327_));
 OA211x2_ASAP7_75t_R _26567_ (.A1(_08326_),
    .A2(_07202_),
    .B(_08327_),
    .C(_07086_),
    .Y(_08328_));
 AO21x1_ASAP7_75t_R _26568_ (.A1(_02384_),
    .A2(_07206_),
    .B(_08328_),
    .Y(_08329_));
 AO22x1_ASAP7_75t_R _26569_ (.A1(net165),
    .A2(_07097_),
    .B1(_08329_),
    .B2(_07094_),
    .Y(_08330_));
 AO221x1_ASAP7_75t_R _26570_ (.A1(_07066_),
    .A2(_07101_),
    .B1(_07640_),
    .B2(_08325_),
    .C(_08330_),
    .Y(_08331_));
 XNOR2x1_ASAP7_75t_R _26571_ (.B(_14025_),
    .Y(_08332_),
    .A(_13656_));
 OR3x1_ASAP7_75t_R _26572_ (.A(_13301_),
    .B(_13656_),
    .C(_14025_),
    .Y(_08333_));
 OA21x2_ASAP7_75t_R _26573_ (.A1(_13302_),
    .A2(_08332_),
    .B(_08333_),
    .Y(_08334_));
 NAND2x1_ASAP7_75t_R _26574_ (.A(_06908_),
    .B(_07523_),
    .Y(_08335_));
 AND4x1_ASAP7_75t_R _26575_ (.A(_14084_),
    .B(_14140_),
    .C(_05661_),
    .D(_08335_),
    .Y(_08336_));
 OR4x1_ASAP7_75t_R _26576_ (.A(_13954_),
    .B(_05558_),
    .C(_08334_),
    .D(_08336_),
    .Y(_08337_));
 NAND2x1_ASAP7_75t_R _26577_ (.A(_05625_),
    .B(_08337_),
    .Y(_08338_));
 OR4x1_ASAP7_75t_R _26578_ (.A(_14139_),
    .B(_05558_),
    .C(_05620_),
    .D(_05664_),
    .Y(_08339_));
 OAI22x1_ASAP7_75t_R _26579_ (.A1(_02148_),
    .A2(net283),
    .B1(net282),
    .B2(_02042_),
    .Y(_08340_));
 NAND2x1_ASAP7_75t_R _26580_ (.A(_05661_),
    .B(_08340_),
    .Y(_08341_));
 AOI21x1_ASAP7_75t_R _26581_ (.A1(_08338_),
    .A2(_08339_),
    .B(_08341_),
    .Y(_08342_));
 NAND2x1_ASAP7_75t_R _26582_ (.A(net143),
    .B(_06889_),
    .Y(_08343_));
 OA22x2_ASAP7_75t_R _26583_ (.A1(_02115_),
    .A2(_06908_),
    .B1(_07523_),
    .B2(_02005_),
    .Y(_08344_));
 OA211x2_ASAP7_75t_R _26584_ (.A1(_01921_),
    .A2(_07513_),
    .B(_08343_),
    .C(_08344_),
    .Y(_08345_));
 OA222x2_ASAP7_75t_R _26585_ (.A1(_01971_),
    .A2(_07145_),
    .B1(_07171_),
    .B2(_02074_),
    .C1(_07305_),
    .C2(_01557_),
    .Y(_08346_));
 OAI21x1_ASAP7_75t_R _26586_ (.A1(_07140_),
    .A2(_08345_),
    .B(_08346_),
    .Y(_08347_));
 OAI22x1_ASAP7_75t_R _26587_ (.A1(_01495_),
    .A2(net283),
    .B1(net282),
    .B2(_01464_),
    .Y(_08348_));
 NAND2x1_ASAP7_75t_R _26588_ (.A(_02249_),
    .B(_07077_),
    .Y(_08349_));
 OA211x2_ASAP7_75t_R _26589_ (.A1(_07686_),
    .A2(_07077_),
    .B(_08349_),
    .C(_07076_),
    .Y(_08350_));
 AO21x1_ASAP7_75t_R _26590_ (.A1(_01077_),
    .A2(_05743_),
    .B(net295),
    .Y(_08351_));
 OA222x2_ASAP7_75t_R _26591_ (.A1(_05684_),
    .A2(_06908_),
    .B1(_08350_),
    .B2(_08351_),
    .C1(_07661_),
    .C2(_01955_),
    .Y(_08352_));
 OAI21x1_ASAP7_75t_R _26592_ (.A1(_00141_),
    .A2(_07151_),
    .B(_08352_),
    .Y(_08353_));
 AO221x1_ASAP7_75t_R _26593_ (.A1(net78),
    .A2(_07155_),
    .B1(_08348_),
    .B2(_06884_),
    .C(_08353_),
    .Y(_08354_));
 OR4x2_ASAP7_75t_R _26594_ (.A(_07113_),
    .B(_08342_),
    .C(_08347_),
    .D(_08354_),
    .Y(_08355_));
 AOI21x1_ASAP7_75t_R _26595_ (.A1(net294),
    .A2(_08331_),
    .B(_08355_),
    .Y(_08356_));
 AOI22x1_ASAP7_75t_R _26596_ (.A1(_08109_),
    .A2(_08323_),
    .B1(_08324_),
    .B2(_08356_),
    .Y(_08357_));
 NOR2x1_ASAP7_75t_R _26597_ (.A(_01685_),
    .B(_06924_),
    .Y(_08358_));
 AO21x1_ASAP7_75t_R _26598_ (.A1(_06924_),
    .A2(_08357_),
    .B(_08358_),
    .Y(_02680_));
 NAND2x1_ASAP7_75t_R _26599_ (.A(_01642_),
    .B(_07746_),
    .Y(_08359_));
 OA211x2_ASAP7_75t_R _26600_ (.A1(_01642_),
    .A2(_07743_),
    .B(_08359_),
    .C(_07117_),
    .Y(_08360_));
 AND2x2_ASAP7_75t_R _26601_ (.A(_06943_),
    .B(_07590_),
    .Y(_08361_));
 AND2x2_ASAP7_75t_R _26602_ (.A(_07592_),
    .B(_08325_),
    .Y(_08362_));
 INVx1_ASAP7_75t_R _26603_ (.A(_00142_),
    .Y(_08363_));
 NAND2x1_ASAP7_75t_R _26604_ (.A(_00143_),
    .B(_07202_),
    .Y(_08364_));
 OA211x2_ASAP7_75t_R _26605_ (.A1(_08363_),
    .A2(_07202_),
    .B(_08364_),
    .C(_07086_),
    .Y(_08365_));
 AO21x1_ASAP7_75t_R _26606_ (.A1(_02385_),
    .A2(net285),
    .B(_08365_),
    .Y(_08366_));
 AO22x1_ASAP7_75t_R _26607_ (.A1(net166),
    .A2(_07097_),
    .B1(_08366_),
    .B2(_07094_),
    .Y(_08367_));
 XOR2x1_ASAP7_75t_R _26608_ (.A(_00055_),
    .Y(_08368_),
    .B(_02248_));
 NAND2x1_ASAP7_75t_R _26609_ (.A(_07079_),
    .B(_07759_),
    .Y(_08369_));
 OA21x2_ASAP7_75t_R _26610_ (.A1(_07079_),
    .A2(_08368_),
    .B(_08369_),
    .Y(_08370_));
 OA21x2_ASAP7_75t_R _26611_ (.A1(_05745_),
    .A2(_08370_),
    .B(_13576_),
    .Y(_08371_));
 NAND2x1_ASAP7_75t_R _26612_ (.A(_01110_),
    .B(_05743_),
    .Y(_08372_));
 AO22x1_ASAP7_75t_R _26613_ (.A1(net295),
    .A2(_08367_),
    .B1(_08371_),
    .B2(_08372_),
    .Y(_08373_));
 OAI22x1_ASAP7_75t_R _26614_ (.A1(_01494_),
    .A2(net283),
    .B1(net282),
    .B2(_01463_),
    .Y(_08374_));
 NAND2x1_ASAP7_75t_R _26615_ (.A(_06884_),
    .B(_08374_),
    .Y(_08375_));
 OAI22x1_ASAP7_75t_R _26616_ (.A1(_02147_),
    .A2(net283),
    .B1(net282),
    .B2(_02041_),
    .Y(_08376_));
 NAND2x1_ASAP7_75t_R _26617_ (.A(_06886_),
    .B(_08376_),
    .Y(_08377_));
 OA222x2_ASAP7_75t_R _26618_ (.A1(_01920_),
    .A2(_07149_),
    .B1(_07171_),
    .B2(_02073_),
    .C1(_05684_),
    .C2(_06908_),
    .Y(_08378_));
 INVx1_ASAP7_75t_R _26619_ (.A(_02114_),
    .Y(_08379_));
 AO22x1_ASAP7_75t_R _26620_ (.A1(_08379_),
    .A2(_05582_),
    .B1(_06889_),
    .B2(net144),
    .Y(_08380_));
 OAI22x1_ASAP7_75t_R _26621_ (.A1(_01954_),
    .A2(_07659_),
    .B1(_07150_),
    .B2(_00144_),
    .Y(_08381_));
 AO222x2_ASAP7_75t_R _26622_ (.A1(net79),
    .A2(_07155_),
    .B1(_08380_),
    .B2(_05630_),
    .C1(_08381_),
    .C2(_05632_),
    .Y(_08382_));
 INVx1_ASAP7_75t_R _26623_ (.A(_08382_),
    .Y(_08383_));
 OA222x2_ASAP7_75t_R _26624_ (.A1(_01970_),
    .A2(_07145_),
    .B1(_07146_),
    .B2(_02004_),
    .C1(_07305_),
    .C2(_01556_),
    .Y(_08384_));
 AND5x2_ASAP7_75t_R _26625_ (.A(_08375_),
    .B(_08377_),
    .C(_08378_),
    .D(_08383_),
    .E(_08384_),
    .Y(_08385_));
 INVx1_ASAP7_75t_R _26626_ (.A(_08385_),
    .Y(_08386_));
 OR4x2_ASAP7_75t_R _26627_ (.A(_07113_),
    .B(_08362_),
    .C(_08373_),
    .D(_08386_),
    .Y(_08387_));
 OA22x2_ASAP7_75t_R _26628_ (.A1(_08037_),
    .A2(_08360_),
    .B1(_08361_),
    .B2(_08387_),
    .Y(_08388_));
 NOR2x1_ASAP7_75t_R _26629_ (.A(_01684_),
    .B(_06924_),
    .Y(_08389_));
 AO21x1_ASAP7_75t_R _26630_ (.A1(_06924_),
    .A2(_08388_),
    .B(_08389_),
    .Y(_02681_));
 AO221x1_ASAP7_75t_R _26631_ (.A1(_07066_),
    .A2(_07550_),
    .B1(_07553_),
    .B2(_07338_),
    .C(_07555_),
    .Y(_08390_));
 NAND2x1_ASAP7_75t_R _26632_ (.A(_06928_),
    .B(_07560_),
    .Y(_08391_));
 INVx1_ASAP7_75t_R _26633_ (.A(_00145_),
    .Y(_08392_));
 NAND2x1_ASAP7_75t_R _26634_ (.A(_00146_),
    .B(_07202_),
    .Y(_08393_));
 OA211x2_ASAP7_75t_R _26635_ (.A1(_08392_),
    .A2(_07202_),
    .B(_08393_),
    .C(_07086_),
    .Y(_08394_));
 AO21x1_ASAP7_75t_R _26636_ (.A1(_02386_),
    .A2(net285),
    .B(_08394_),
    .Y(_08395_));
 AOI22x1_ASAP7_75t_R _26637_ (.A1(net167),
    .A2(_07097_),
    .B1(_08395_),
    .B2(_07094_),
    .Y(_08396_));
 AND2x2_ASAP7_75t_R _26638_ (.A(_02237_),
    .B(_07079_),
    .Y(_08397_));
 AO221x2_ASAP7_75t_R _26639_ (.A1(_13317_),
    .A2(_05743_),
    .B1(_07077_),
    .B2(_02251_),
    .C(_08397_),
    .Y(_08398_));
 NAND2x1_ASAP7_75t_R _26640_ (.A(_13576_),
    .B(_08398_),
    .Y(_08399_));
 AO21x1_ASAP7_75t_R _26641_ (.A1(_01142_),
    .A2(_05743_),
    .B(_08399_),
    .Y(_08400_));
 OAI22x1_ASAP7_75t_R _26642_ (.A1(_02146_),
    .A2(net283),
    .B1(net282),
    .B2(_02040_),
    .Y(_08401_));
 NAND2x1_ASAP7_75t_R _26643_ (.A(_06886_),
    .B(_08401_),
    .Y(_08402_));
 OAI22x1_ASAP7_75t_R _26644_ (.A1(_01493_),
    .A2(net283),
    .B1(net282),
    .B2(_01462_),
    .Y(_08403_));
 NAND2x1_ASAP7_75t_R _26645_ (.A(_06884_),
    .B(_08403_),
    .Y(_08404_));
 OR3x1_ASAP7_75t_R _26646_ (.A(_06236_),
    .B(_07507_),
    .C(_07659_),
    .Y(_08405_));
 NAND2x1_ASAP7_75t_R _26647_ (.A(net80),
    .B(_06891_),
    .Y(_08406_));
 OA21x2_ASAP7_75t_R _26648_ (.A1(_02113_),
    .A2(_07508_),
    .B(_07168_),
    .Y(_08407_));
 OA222x2_ASAP7_75t_R _26649_ (.A1(_01919_),
    .A2(_07701_),
    .B1(_07524_),
    .B2(_02003_),
    .C1(_02072_),
    .C2(_07505_),
    .Y(_08408_));
 AND4x1_ASAP7_75t_R _26650_ (.A(_08405_),
    .B(_08406_),
    .C(_08407_),
    .D(_08408_),
    .Y(_08409_));
 OA22x2_ASAP7_75t_R _26651_ (.A1(_00147_),
    .A2(_07705_),
    .B1(_07516_),
    .B2(_01555_),
    .Y(_08410_));
 OA22x2_ASAP7_75t_R _26652_ (.A1(_01969_),
    .A2(_07511_),
    .B1(_07661_),
    .B2(_01953_),
    .Y(_08411_));
 AND5x2_ASAP7_75t_R _26653_ (.A(_08402_),
    .B(_08404_),
    .C(_08409_),
    .D(_08410_),
    .E(_08411_),
    .Y(_08412_));
 OA211x2_ASAP7_75t_R _26654_ (.A1(_13576_),
    .A2(_08396_),
    .B(_08400_),
    .C(_08412_),
    .Y(_08413_));
 NAND2x1_ASAP7_75t_R _26655_ (.A(_06920_),
    .B(_08413_),
    .Y(_08414_));
 AO221x1_ASAP7_75t_R _26656_ (.A1(_06943_),
    .A2(_08390_),
    .B1(_08141_),
    .B2(_08391_),
    .C(_08414_),
    .Y(_08415_));
 NOR2x1_ASAP7_75t_R _26657_ (.A(net418),
    .B(_07808_),
    .Y(_08416_));
 AO21x1_ASAP7_75t_R _26658_ (.A1(net418),
    .A2(_07806_),
    .B(_08416_),
    .Y(_08417_));
 AO21x1_ASAP7_75t_R _26659_ (.A1(_07117_),
    .A2(_08417_),
    .B(_08037_),
    .Y(_08418_));
 AND2x6_ASAP7_75t_R _26660_ (.A(_08415_),
    .B(_08418_),
    .Y(_08419_));
 NOR2x1_ASAP7_75t_R _26661_ (.A(_01683_),
    .B(_06924_),
    .Y(_08420_));
 AO21x1_ASAP7_75t_R _26662_ (.A1(_06924_),
    .A2(_08419_),
    .B(_08420_),
    .Y(_02682_));
 INVx1_ASAP7_75t_R _26663_ (.A(_00148_),
    .Y(_08421_));
 NAND2x1_ASAP7_75t_R _26664_ (.A(_00149_),
    .B(_07202_),
    .Y(_08422_));
 OA211x2_ASAP7_75t_R _26665_ (.A1(_08421_),
    .A2(_07202_),
    .B(_08422_),
    .C(_07086_),
    .Y(_08423_));
 AO21x1_ASAP7_75t_R _26666_ (.A1(_02387_),
    .A2(_07206_),
    .B(_08423_),
    .Y(_08424_));
 AO221x1_ASAP7_75t_R _26667_ (.A1(net168),
    .A2(_07097_),
    .B1(_08424_),
    .B2(_07094_),
    .C(_13576_),
    .Y(_08425_));
 OA21x2_ASAP7_75t_R _26668_ (.A1(_07100_),
    .A2(_07408_),
    .B(_08325_),
    .Y(_08426_));
 XNOR2x1_ASAP7_75t_R _26669_ (.B(_02250_),
    .Y(_08427_),
    .A(_00058_));
 NAND2x1_ASAP7_75t_R _26670_ (.A(_07077_),
    .B(_08427_),
    .Y(_08428_));
 OAI21x1_ASAP7_75t_R _26671_ (.A1(_07077_),
    .A2(_07824_),
    .B(_08428_),
    .Y(_08429_));
 NAND2x1_ASAP7_75t_R _26672_ (.A(_07076_),
    .B(_08429_),
    .Y(_08430_));
 NAND2x1_ASAP7_75t_R _26673_ (.A(_01176_),
    .B(_05743_),
    .Y(_08431_));
 AO21x1_ASAP7_75t_R _26674_ (.A1(_08430_),
    .A2(_08431_),
    .B(net295),
    .Y(_08432_));
 OAI21x1_ASAP7_75t_R _26675_ (.A1(_08425_),
    .A2(_08426_),
    .B(_08432_),
    .Y(_08433_));
 OAI22x1_ASAP7_75t_R _26676_ (.A1(_02145_),
    .A2(net283),
    .B1(net282),
    .B2(_02039_),
    .Y(_08434_));
 NAND2x1_ASAP7_75t_R _26677_ (.A(_06886_),
    .B(_08434_),
    .Y(_08435_));
 OAI22x1_ASAP7_75t_R _26678_ (.A1(_01492_),
    .A2(net283),
    .B1(net282),
    .B2(_01461_),
    .Y(_08436_));
 NAND2x1_ASAP7_75t_R _26679_ (.A(_06884_),
    .B(_08436_),
    .Y(_08437_));
 NAND2x1_ASAP7_75t_R _26680_ (.A(net81),
    .B(_06891_),
    .Y(_08438_));
 OA211x2_ASAP7_75t_R _26681_ (.A1(_01952_),
    .A2(_07661_),
    .B(_08438_),
    .C(_07168_),
    .Y(_08439_));
 INVx1_ASAP7_75t_R _26682_ (.A(net132),
    .Y(_08440_));
 OA222x2_ASAP7_75t_R _26683_ (.A1(_02071_),
    .A2(_07505_),
    .B1(_07511_),
    .B2(_01968_),
    .C1(_08440_),
    .C2(_08098_),
    .Y(_08441_));
 OA211x2_ASAP7_75t_R _26684_ (.A1(_02112_),
    .A2(_07508_),
    .B(_08439_),
    .C(_08441_),
    .Y(_08442_));
 OA22x2_ASAP7_75t_R _26685_ (.A1(_00150_),
    .A2(_07705_),
    .B1(_07701_),
    .B2(_01918_),
    .Y(_08443_));
 OA22x2_ASAP7_75t_R _26686_ (.A1(_02002_),
    .A2(_07524_),
    .B1(_07516_),
    .B2(_01554_),
    .Y(_08444_));
 AND5x2_ASAP7_75t_R _26687_ (.A(_08435_),
    .B(_08437_),
    .C(_08442_),
    .D(_08443_),
    .E(_08444_),
    .Y(_08445_));
 NAND2x1_ASAP7_75t_R _26688_ (.A(_06943_),
    .B(_07492_),
    .Y(_08446_));
 AND4x2_ASAP7_75t_R _26689_ (.A(_06920_),
    .B(_08433_),
    .C(_08445_),
    .D(_08446_),
    .Y(_08447_));
 NAND2x1_ASAP7_75t_R _26690_ (.A(_01642_),
    .B(_07853_),
    .Y(_08448_));
 OA21x2_ASAP7_75t_R _26691_ (.A1(_01642_),
    .A2(_07856_),
    .B(_08448_),
    .Y(_08449_));
 OA21x2_ASAP7_75t_R _26692_ (.A1(_07115_),
    .A2(_08449_),
    .B(_08109_),
    .Y(_08450_));
 NOR2x2_ASAP7_75t_R _26693_ (.A(_08447_),
    .B(_08450_),
    .Y(_08451_));
 NOR2x1_ASAP7_75t_R _26694_ (.A(_01682_),
    .B(_06924_),
    .Y(_08452_));
 AO21x1_ASAP7_75t_R _26695_ (.A1(_06924_),
    .A2(_08451_),
    .B(_08452_),
    .Y(_02683_));
 NOR2x1_ASAP7_75t_R _26696_ (.A(net418),
    .B(_07900_),
    .Y(_08453_));
 AO21x1_ASAP7_75t_R _26697_ (.A1(net418),
    .A2(_07898_),
    .B(_08453_),
    .Y(_08454_));
 AO21x1_ASAP7_75t_R _26698_ (.A1(_07117_),
    .A2(_08454_),
    .B(_08037_),
    .Y(_08455_));
 NAND2x1_ASAP7_75t_R _26699_ (.A(_02253_),
    .B(_07077_),
    .Y(_08456_));
 OA211x2_ASAP7_75t_R _26700_ (.A1(_07872_),
    .A2(_07077_),
    .B(_08456_),
    .C(_07076_),
    .Y(_08457_));
 AO21x1_ASAP7_75t_R _26701_ (.A1(_01208_),
    .A2(_05743_),
    .B(_08457_),
    .Y(_08458_));
 NAND2x1_ASAP7_75t_R _26702_ (.A(_13576_),
    .B(_08458_),
    .Y(_08459_));
 NAND2x1_ASAP7_75t_R _26703_ (.A(_06928_),
    .B(_07432_),
    .Y(_08460_));
 INVx1_ASAP7_75t_R _26704_ (.A(_00151_),
    .Y(_08461_));
 NAND2x1_ASAP7_75t_R _26705_ (.A(_00152_),
    .B(_07202_),
    .Y(_08462_));
 OA211x2_ASAP7_75t_R _26706_ (.A1(_08461_),
    .A2(_07202_),
    .B(_08462_),
    .C(_07086_),
    .Y(_08463_));
 AO21x1_ASAP7_75t_R _26707_ (.A1(_02388_),
    .A2(net285),
    .B(_08463_),
    .Y(_08464_));
 AO22x1_ASAP7_75t_R _26708_ (.A1(net169),
    .A2(_07097_),
    .B1(_08464_),
    .B2(_07094_),
    .Y(_08465_));
 AO221x1_ASAP7_75t_R _26709_ (.A1(_13313_),
    .A2(_13317_),
    .B1(_08141_),
    .B2(_08460_),
    .C(_08465_),
    .Y(_08466_));
 OA222x2_ASAP7_75t_R _26710_ (.A1(_02001_),
    .A2(_07146_),
    .B1(_07299_),
    .B2(_02111_),
    .C1(_05684_),
    .C2(_06908_),
    .Y(_08467_));
 OA22x2_ASAP7_75t_R _26711_ (.A1(_00153_),
    .A2(_07151_),
    .B1(_07149_),
    .B2(_01917_),
    .Y(_08468_));
 OA22x2_ASAP7_75t_R _26712_ (.A1(_01967_),
    .A2(_07145_),
    .B1(_07305_),
    .B2(_01553_),
    .Y(_08469_));
 NAND2x1_ASAP7_75t_R _26713_ (.A(net82),
    .B(_07155_),
    .Y(_08470_));
 AND4x2_ASAP7_75t_R _26714_ (.A(_08467_),
    .B(_08468_),
    .C(_08469_),
    .D(_08470_),
    .Y(_08471_));
 OAI22x1_ASAP7_75t_R _26715_ (.A1(_01491_),
    .A2(net283),
    .B1(net282),
    .B2(_01460_),
    .Y(_08472_));
 NAND2x1_ASAP7_75t_R _26716_ (.A(_06884_),
    .B(_08472_),
    .Y(_08473_));
 OAI22x1_ASAP7_75t_R _26717_ (.A1(_02144_),
    .A2(net283),
    .B1(net282),
    .B2(_02038_),
    .Y(_08474_));
 NAND2x1_ASAP7_75t_R _26718_ (.A(_06886_),
    .B(_08474_),
    .Y(_08475_));
 INVx1_ASAP7_75t_R _26719_ (.A(net133),
    .Y(_08476_));
 OA222x2_ASAP7_75t_R _26720_ (.A1(_02070_),
    .A2(_07171_),
    .B1(_07661_),
    .B2(_01951_),
    .C1(_08476_),
    .C2(_07663_),
    .Y(_08477_));
 AND4x2_ASAP7_75t_R _26721_ (.A(_08471_),
    .B(_08473_),
    .C(_08475_),
    .D(_08477_),
    .Y(_08478_));
 NAND2x1_ASAP7_75t_R _26722_ (.A(_06920_),
    .B(_08478_),
    .Y(_08479_));
 AO221x2_ASAP7_75t_R _26723_ (.A1(_06943_),
    .A2(_07423_),
    .B1(_08459_),
    .B2(_08466_),
    .C(_08479_),
    .Y(_08480_));
 AND2x6_ASAP7_75t_R _26724_ (.A(_08455_),
    .B(_08480_),
    .Y(_08481_));
 NOR2x1_ASAP7_75t_R _26725_ (.A(_01681_),
    .B(_06924_),
    .Y(_08482_));
 AO21x1_ASAP7_75t_R _26726_ (.A1(_06924_),
    .A2(_08481_),
    .B(_08482_),
    .Y(_02684_));
 NOR2x1_ASAP7_75t_R _26727_ (.A(_01642_),
    .B(_07942_),
    .Y(_08483_));
 AO21x1_ASAP7_75t_R _26728_ (.A1(_01642_),
    .A2(_07939_),
    .B(_08483_),
    .Y(_08484_));
 AO21x1_ASAP7_75t_R _26729_ (.A1(_07117_),
    .A2(_08484_),
    .B(_08037_),
    .Y(_08485_));
 INVx1_ASAP7_75t_R _26730_ (.A(_00154_),
    .Y(_08486_));
 NAND2x1_ASAP7_75t_R _26731_ (.A(_00155_),
    .B(_07202_),
    .Y(_08487_));
 OA211x2_ASAP7_75t_R _26732_ (.A1(_08486_),
    .A2(_07202_),
    .B(_08487_),
    .C(_07086_),
    .Y(_08488_));
 AO21x1_ASAP7_75t_R _26733_ (.A1(_02389_),
    .A2(net285),
    .B(_08488_),
    .Y(_08489_));
 OA21x2_ASAP7_75t_R _26734_ (.A1(_07066_),
    .A2(_07347_),
    .B(_08141_),
    .Y(_08490_));
 AO221x1_ASAP7_75t_R _26735_ (.A1(net2114),
    .A2(_07097_),
    .B1(_08489_),
    .B2(_07094_),
    .C(_08490_),
    .Y(_08491_));
 XNOR2x1_ASAP7_75t_R _26736_ (.B(_02252_),
    .Y(_08492_),
    .A(_00061_));
 NAND2x1_ASAP7_75t_R _26737_ (.A(_07077_),
    .B(_08492_),
    .Y(_08493_));
 OAI21x1_ASAP7_75t_R _26738_ (.A1(_07077_),
    .A2(_07916_),
    .B(_08493_),
    .Y(_08494_));
 AO21x1_ASAP7_75t_R _26739_ (.A1(_07076_),
    .A2(_08494_),
    .B(_13318_),
    .Y(_08495_));
 AOI21x1_ASAP7_75t_R _26740_ (.A1(_01242_),
    .A2(_05743_),
    .B(_08495_),
    .Y(_08496_));
 OAI22x1_ASAP7_75t_R _26741_ (.A1(_01490_),
    .A2(net283),
    .B1(net282),
    .B2(_01459_),
    .Y(_08497_));
 OAI22x1_ASAP7_75t_R _26742_ (.A1(_02143_),
    .A2(net283),
    .B1(net282),
    .B2(_02037_),
    .Y(_08498_));
 OAI22x1_ASAP7_75t_R _26743_ (.A1(_02069_),
    .A2(_07171_),
    .B1(_07663_),
    .B2(_06281_),
    .Y(_08499_));
 OAI22x1_ASAP7_75t_R _26744_ (.A1(_01966_),
    .A2(_07145_),
    .B1(_07305_),
    .B2(_01552_),
    .Y(_08500_));
 INVx1_ASAP7_75t_R _26745_ (.A(_02000_),
    .Y(_08501_));
 AO32x1_ASAP7_75t_R _26746_ (.A1(_08501_),
    .A2(_05630_),
    .A3(_07144_),
    .B1(_05539_),
    .B2(_05582_),
    .Y(_08502_));
 OR3x2_ASAP7_75t_R _26747_ (.A(_08499_),
    .B(_08500_),
    .C(_08502_),
    .Y(_08503_));
 AOI221x1_ASAP7_75t_R _26748_ (.A1(_06884_),
    .A2(_08497_),
    .B1(_08498_),
    .B2(_06886_),
    .C(_08503_),
    .Y(_08504_));
 OAI22x1_ASAP7_75t_R _26749_ (.A1(_02110_),
    .A2(_06908_),
    .B1(_07513_),
    .B2(_01916_),
    .Y(_08505_));
 OAI22x1_ASAP7_75t_R _26750_ (.A1(_01950_),
    .A2(_07659_),
    .B1(_07150_),
    .B2(_00156_),
    .Y(_08506_));
 AO222x2_ASAP7_75t_R _26751_ (.A1(net83),
    .A2(_07155_),
    .B1(_08505_),
    .B2(_05630_),
    .C1(_08506_),
    .C2(_05632_),
    .Y(_08507_));
 INVx1_ASAP7_75t_R _26752_ (.A(_08507_),
    .Y(_08508_));
 NAND2x2_ASAP7_75t_R _26753_ (.A(_08504_),
    .B(_08508_),
    .Y(_08509_));
 OR3x1_ASAP7_75t_R _26754_ (.A(_07113_),
    .B(_08496_),
    .C(_08509_),
    .Y(_08510_));
 AO221x1_ASAP7_75t_R _26755_ (.A1(_06943_),
    .A2(_07345_),
    .B1(_08491_),
    .B2(net294),
    .C(_08510_),
    .Y(_08511_));
 AND2x6_ASAP7_75t_R _26756_ (.A(_08485_),
    .B(_08511_),
    .Y(_08512_));
 NOR2x1_ASAP7_75t_R _26757_ (.A(_01680_),
    .B(_06924_),
    .Y(_08513_));
 AO21x1_ASAP7_75t_R _26758_ (.A1(_06924_),
    .A2(_08512_),
    .B(_08513_),
    .Y(_02685_));
 NAND2x1_ASAP7_75t_R _26759_ (.A(net418),
    .B(_07979_),
    .Y(_08514_));
 OA21x2_ASAP7_75t_R _26760_ (.A1(net418),
    .A2(_07982_),
    .B(_08514_),
    .Y(_08515_));
 OA21x2_ASAP7_75t_R _26761_ (.A1(_07115_),
    .A2(_08515_),
    .B(_08109_),
    .Y(_08516_));
 INVx1_ASAP7_75t_R _26762_ (.A(_02241_),
    .Y(_08517_));
 NAND2x1_ASAP7_75t_R _26763_ (.A(_02255_),
    .B(_07077_),
    .Y(_08518_));
 OA211x2_ASAP7_75t_R _26764_ (.A1(_08517_),
    .A2(_07077_),
    .B(_08518_),
    .C(_07076_),
    .Y(_08519_));
 AOI21x1_ASAP7_75t_R _26765_ (.A1(_01274_),
    .A2(_05743_),
    .B(_08519_),
    .Y(_08520_));
 OA21x2_ASAP7_75t_R _26766_ (.A1(_07100_),
    .A2(_07216_),
    .B(_08325_),
    .Y(_08521_));
 INVx1_ASAP7_75t_R _26767_ (.A(_00157_),
    .Y(_08522_));
 NAND2x1_ASAP7_75t_R _26768_ (.A(_00158_),
    .B(_07202_),
    .Y(_08523_));
 OA211x2_ASAP7_75t_R _26769_ (.A1(_08522_),
    .A2(_07202_),
    .B(_08523_),
    .C(_07086_),
    .Y(_08524_));
 AO21x1_ASAP7_75t_R _26770_ (.A1(_02390_),
    .A2(net285),
    .B(_08524_),
    .Y(_08525_));
 AO22x1_ASAP7_75t_R _26771_ (.A1(net172),
    .A2(_07097_),
    .B1(_08525_),
    .B2(_07094_),
    .Y(_08526_));
 OR3x1_ASAP7_75t_R _26772_ (.A(_13576_),
    .B(_08521_),
    .C(_08526_),
    .Y(_08527_));
 OAI21x1_ASAP7_75t_R _26773_ (.A1(net294),
    .A2(_08520_),
    .B(_08527_),
    .Y(_08528_));
 NAND2x1_ASAP7_75t_R _26774_ (.A(_06943_),
    .B(_07257_),
    .Y(_08529_));
 OAI22x1_ASAP7_75t_R _26775_ (.A1(_01489_),
    .A2(net283),
    .B1(net282),
    .B2(_01458_),
    .Y(_08530_));
 NAND2x1_ASAP7_75t_R _26776_ (.A(_06884_),
    .B(_08530_),
    .Y(_08531_));
 OAI22x1_ASAP7_75t_R _26777_ (.A1(_02142_),
    .A2(net283),
    .B1(net282),
    .B2(_02036_),
    .Y(_08532_));
 NAND2x1_ASAP7_75t_R _26778_ (.A(_06886_),
    .B(_08532_),
    .Y(_08533_));
 OA21x2_ASAP7_75t_R _26779_ (.A1(_01551_),
    .A2(_07305_),
    .B(_07172_),
    .Y(_08534_));
 AOI22x1_ASAP7_75t_R _26780_ (.A1(_06206_),
    .A2(_05632_),
    .B1(_05630_),
    .B2(net135),
    .Y(_08535_));
 OA22x2_ASAP7_75t_R _26781_ (.A1(_02068_),
    .A2(_07171_),
    .B1(_08535_),
    .B2(_07659_),
    .Y(_08536_));
 OA211x2_ASAP7_75t_R _26782_ (.A1(_02109_),
    .A2(_07299_),
    .B(_08534_),
    .C(_08536_),
    .Y(_08537_));
 OAI22x1_ASAP7_75t_R _26783_ (.A1(_01999_),
    .A2(_07146_),
    .B1(_07149_),
    .B2(_01915_),
    .Y(_08538_));
 OAI22x1_ASAP7_75t_R _26784_ (.A1(_01965_),
    .A2(_07145_),
    .B1(_07151_),
    .B2(_00159_),
    .Y(_08539_));
 OR3x4_ASAP7_75t_R _26785_ (.A(_07699_),
    .B(_08538_),
    .C(_08539_),
    .Y(_08540_));
 AOI21x1_ASAP7_75t_R _26786_ (.A1(net85),
    .A2(_07155_),
    .B(_08540_),
    .Y(_08541_));
 AND4x2_ASAP7_75t_R _26787_ (.A(_08531_),
    .B(_08533_),
    .C(_08537_),
    .D(_08541_),
    .Y(_08542_));
 OA211x2_ASAP7_75t_R _26788_ (.A1(_07283_),
    .A2(_07430_),
    .B(_08542_),
    .C(_06920_),
    .Y(_08543_));
 AND3x2_ASAP7_75t_R _26789_ (.A(_08528_),
    .B(_08529_),
    .C(_08543_),
    .Y(_08544_));
 NOR2x2_ASAP7_75t_R _26790_ (.A(_08516_),
    .B(_08544_),
    .Y(_08545_));
 NOR2x1_ASAP7_75t_R _26791_ (.A(_01679_),
    .B(_06924_),
    .Y(_08546_));
 AO21x1_ASAP7_75t_R _26792_ (.A1(_06924_),
    .A2(_08545_),
    .B(_08546_),
    .Y(_02686_));
 XNOR2x1_ASAP7_75t_R _26793_ (.B(_02254_),
    .Y(_08547_),
    .A(_00064_));
 NAND2x1_ASAP7_75t_R _26794_ (.A(_07077_),
    .B(_08547_),
    .Y(_08548_));
 OA211x2_ASAP7_75t_R _26795_ (.A1(_07077_),
    .A2(_08002_),
    .B(_08548_),
    .C(_07076_),
    .Y(_08549_));
 AND3x1_ASAP7_75t_R _26796_ (.A(_05503_),
    .B(_13317_),
    .C(_05743_),
    .Y(_08550_));
 OA21x2_ASAP7_75t_R _26797_ (.A1(_07100_),
    .A2(_07106_),
    .B(_08325_),
    .Y(_08551_));
 INVx1_ASAP7_75t_R _26798_ (.A(_01310_),
    .Y(_08552_));
 NAND2x1_ASAP7_75t_R _26799_ (.A(_00160_),
    .B(_07202_),
    .Y(_08553_));
 OA211x2_ASAP7_75t_R _26800_ (.A1(_08552_),
    .A2(_07202_),
    .B(_08553_),
    .C(_07086_),
    .Y(_08554_));
 AO21x1_ASAP7_75t_R _26801_ (.A1(_02282_),
    .A2(_07206_),
    .B(_08554_),
    .Y(_08555_));
 AO221x1_ASAP7_75t_R _26802_ (.A1(net173),
    .A2(_07097_),
    .B1(_08555_),
    .B2(_07094_),
    .C(_13576_),
    .Y(_08556_));
 OA221x2_ASAP7_75t_R _26803_ (.A1(_06928_),
    .A2(_07012_),
    .B1(_07054_),
    .B2(_07068_),
    .C(_06943_),
    .Y(_08557_));
 OA33x2_ASAP7_75t_R _26804_ (.A1(net294),
    .A2(_08549_),
    .A3(_08550_),
    .B1(_08551_),
    .B2(_08556_),
    .B3(_08557_),
    .Y(_08558_));
 OAI22x1_ASAP7_75t_R _26805_ (.A1(_01488_),
    .A2(net283),
    .B1(net282),
    .B2(_01457_),
    .Y(_08559_));
 OAI22x1_ASAP7_75t_R _26806_ (.A1(_02141_),
    .A2(net283),
    .B1(net282),
    .B2(_02035_),
    .Y(_08560_));
 AOI22x1_ASAP7_75t_R _26807_ (.A1(_06884_),
    .A2(_08559_),
    .B1(_08560_),
    .B2(_06886_),
    .Y(_08561_));
 OA22x2_ASAP7_75t_R _26808_ (.A1(_02067_),
    .A2(_07171_),
    .B1(_07299_),
    .B2(_02108_),
    .Y(_08562_));
 OR3x1_ASAP7_75t_R _26809_ (.A(_01908_),
    .B(_07140_),
    .C(_07142_),
    .Y(_08563_));
 OA21x2_ASAP7_75t_R _26810_ (.A1(_01914_),
    .A2(_07149_),
    .B(_08563_),
    .Y(_08564_));
 OA211x2_ASAP7_75t_R _26811_ (.A1(_00161_),
    .A2(_07151_),
    .B(_07168_),
    .C(_08564_),
    .Y(_08565_));
 NAND2x1_ASAP7_75t_R _26812_ (.A(net86),
    .B(_07155_),
    .Y(_08566_));
 OA222x2_ASAP7_75t_R _26813_ (.A1(_01964_),
    .A2(_07145_),
    .B1(_07146_),
    .B2(_01998_),
    .C1(_07305_),
    .C2(_01550_),
    .Y(_08567_));
 AND5x2_ASAP7_75t_R _26814_ (.A(_08561_),
    .B(_08562_),
    .C(_08565_),
    .D(_08566_),
    .E(_08567_),
    .Y(_08568_));
 NAND2x1_ASAP7_75t_R _26815_ (.A(_06920_),
    .B(_08568_),
    .Y(_08569_));
 NOR2x1_ASAP7_75t_R _26816_ (.A(_07120_),
    .B(_08025_),
    .Y(_08570_));
 OA211x2_ASAP7_75t_R _26817_ (.A1(net42),
    .A2(net419),
    .B(_08021_),
    .C(_07120_),
    .Y(_08571_));
 OA21x2_ASAP7_75t_R _26818_ (.A1(_08570_),
    .A2(_08571_),
    .B(_07117_),
    .Y(_08572_));
 OA22x2_ASAP7_75t_R _26819_ (.A1(_08558_),
    .A2(_08569_),
    .B1(_08572_),
    .B2(_08037_),
    .Y(_08573_));
 NOR2x1_ASAP7_75t_R _26820_ (.A(_01678_),
    .B(_06924_),
    .Y(_08574_));
 AO21x1_ASAP7_75t_R _26821_ (.A1(_06924_),
    .A2(_08573_),
    .B(_08574_),
    .Y(_02687_));
 TAPCELL_ASAP7_75t_R TAP_705 ();
 NAND2x2_ASAP7_75t_R _26823_ (.A(_01873_),
    .B(_13527_),
    .Y(_08576_));
 AND2x4_ASAP7_75t_R _26824_ (.A(_05474_),
    .B(_05915_),
    .Y(_08577_));
 NAND2x1_ASAP7_75t_R _26825_ (.A(_00282_),
    .B(_05743_),
    .Y(_08578_));
 NAND2x1_ASAP7_75t_R _26826_ (.A(_05907_),
    .B(_13327_),
    .Y(_08579_));
 AND4x2_ASAP7_75t_R _26827_ (.A(_13313_),
    .B(_05420_),
    .C(_05517_),
    .D(_08579_),
    .Y(_08580_));
 INVx11_ASAP7_75t_R _26828_ (.A(_08580_),
    .Y(_08581_));
 NAND2x2_ASAP7_75t_R _26829_ (.A(_05474_),
    .B(_05915_),
    .Y(_08582_));
 AND4x1_ASAP7_75t_R _26830_ (.A(_00282_),
    .B(_05743_),
    .C(_08582_),
    .D(_08580_),
    .Y(_08583_));
 AO21x1_ASAP7_75t_R _26831_ (.A1(_08577_),
    .A2(_08581_),
    .B(_08583_),
    .Y(_08584_));
 INVx1_ASAP7_75t_R _26832_ (.A(_01519_),
    .Y(_08585_));
 OA211x2_ASAP7_75t_R _26833_ (.A1(_00283_),
    .A2(_13350_),
    .B(_13317_),
    .C(_08585_),
    .Y(_08586_));
 INVx1_ASAP7_75t_R _26834_ (.A(_08586_),
    .Y(_08587_));
 AO221x1_ASAP7_75t_R _26835_ (.A1(_08577_),
    .A2(_08578_),
    .B1(_08584_),
    .B2(_08587_),
    .C(_00285_),
    .Y(_08588_));
 OA21x2_ASAP7_75t_R _26836_ (.A1(_05778_),
    .A2(_08576_),
    .B(_08588_),
    .Y(_08589_));
 OAI21x1_ASAP7_75t_R _26837_ (.A1(_07076_),
    .A2(_08589_),
    .B(_14626_),
    .Y(_08590_));
 CKINVDCx20_ASAP7_75t_R _26838_ (.A(_08590_),
    .Y(_08591_));
 TAPCELL_ASAP7_75t_R TAP_704 ();
 TAPCELL_ASAP7_75t_R TAP_703 ();
 TAPCELL_ASAP7_75t_R TAP_702 ();
 TAPCELL_ASAP7_75t_R TAP_701 ();
 AND2x2_ASAP7_75t_R _26843_ (.A(_00324_),
    .B(_07079_),
    .Y(_08596_));
 AO21x1_ASAP7_75t_R _26844_ (.A1(_01356_),
    .A2(_07077_),
    .B(_08596_),
    .Y(_08597_));
 AND3x4_ASAP7_75t_R _26845_ (.A(_00282_),
    .B(_05517_),
    .C(_05743_),
    .Y(_08598_));
 TAPCELL_ASAP7_75t_R TAP_700 ();
 OR3x4_ASAP7_75t_R _26847_ (.A(_07076_),
    .B(_08576_),
    .C(_08598_),
    .Y(_08600_));
 TAPCELL_ASAP7_75t_R TAP_699 ();
 TAPCELL_ASAP7_75t_R TAP_698 ();
 NOR2x1_ASAP7_75t_R _26850_ (.A(_13758_),
    .B(_08600_),
    .Y(_08603_));
 AO21x1_ASAP7_75t_R _26851_ (.A1(_07076_),
    .A2(_08597_),
    .B(_08603_),
    .Y(_08604_));
 TAPCELL_ASAP7_75t_R TAP_697 ();
 INVx1_ASAP7_75t_R _26853_ (.A(_02202_),
    .Y(_08606_));
 MAJx3_ASAP7_75t_R _26854_ (.A(_01308_),
    .B(_08606_),
    .C(net173),
    .Y(_08607_));
 OR3x4_ASAP7_75t_R _26855_ (.A(_05751_),
    .B(_05750_),
    .C(_08607_),
    .Y(_08608_));
 OA211x2_ASAP7_75t_R _26856_ (.A1(_01321_),
    .A2(_08608_),
    .B(_08598_),
    .C(_01323_),
    .Y(_08609_));
 OR3x4_ASAP7_75t_R _26857_ (.A(_00279_),
    .B(_13323_),
    .C(net295),
    .Y(_08610_));
 TAPCELL_ASAP7_75t_R TAP_696 ();
 TAPCELL_ASAP7_75t_R TAP_695 ();
 TAPCELL_ASAP7_75t_R TAP_694 ();
 MAJx3_ASAP7_75t_R _26861_ (.A(_05503_),
    .B(_02202_),
    .C(_05512_),
    .Y(_08614_));
 TAPCELL_ASAP7_75t_R TAP_693 ();
 AND2x2_ASAP7_75t_R _26863_ (.A(_16503_),
    .B(_08614_),
    .Y(_08616_));
 AO21x1_ASAP7_75t_R _26864_ (.A1(_00324_),
    .A2(_08607_),
    .B(_08616_),
    .Y(_08617_));
 AO21x1_ASAP7_75t_R _26865_ (.A1(_08610_),
    .A2(_08617_),
    .B(_01727_),
    .Y(_08618_));
 TAPCELL_ASAP7_75t_R TAP_692 ();
 TAPCELL_ASAP7_75t_R TAP_691 ();
 INVx3_ASAP7_75t_R _26868_ (.A(net299),
    .Y(_08621_));
 AND2x2_ASAP7_75t_R _26869_ (.A(net299),
    .B(_01674_),
    .Y(_08622_));
 AO21x1_ASAP7_75t_R _26870_ (.A1(_08621_),
    .A2(_01676_),
    .B(_08622_),
    .Y(_08623_));
 TAPCELL_ASAP7_75t_R TAP_690 ();
 INVx1_ASAP7_75t_R _26872_ (.A(_01675_),
    .Y(_08625_));
 NAND2x1_ASAP7_75t_R _26873_ (.A(net299),
    .B(_01673_),
    .Y(_08626_));
 OA211x2_ASAP7_75t_R _26874_ (.A1(net299),
    .A2(_08625_),
    .B(_08626_),
    .C(_17600_),
    .Y(_08627_));
 INVx1_ASAP7_75t_R _26875_ (.A(_08627_),
    .Y(_08628_));
 XNOR2x2_ASAP7_75t_R _26876_ (.A(_01322_),
    .B(_02292_),
    .Y(_08629_));
 OA211x2_ASAP7_75t_R _26877_ (.A1(_17600_),
    .A2(_08623_),
    .B(_08628_),
    .C(_08629_),
    .Y(_08630_));
 AND2x2_ASAP7_75t_R _26878_ (.A(net299),
    .B(_01666_),
    .Y(_08631_));
 AO21x1_ASAP7_75t_R _26879_ (.A1(_08621_),
    .A2(_01668_),
    .B(_08631_),
    .Y(_08632_));
 INVx1_ASAP7_75t_R _26880_ (.A(_01667_),
    .Y(_08633_));
 NAND2x1_ASAP7_75t_R _26881_ (.A(net299),
    .B(_01665_),
    .Y(_08634_));
 OA211x2_ASAP7_75t_R _26882_ (.A1(net299),
    .A2(_08633_),
    .B(_08634_),
    .C(_17600_),
    .Y(_08635_));
 INVx1_ASAP7_75t_R _26883_ (.A(_08635_),
    .Y(_08636_));
 INVx2_ASAP7_75t_R _26884_ (.A(_08629_),
    .Y(_08637_));
 OA211x2_ASAP7_75t_R _26885_ (.A1(_17600_),
    .A2(_08632_),
    .B(_08636_),
    .C(_08637_),
    .Y(_08638_));
 OR3x1_ASAP7_75t_R _26886_ (.A(_02293_),
    .B(_08630_),
    .C(_08638_),
    .Y(_08639_));
 INVx1_ASAP7_75t_R _26887_ (.A(_01672_),
    .Y(_08640_));
 NAND2x1_ASAP7_75t_R _26888_ (.A(net299),
    .B(_01670_),
    .Y(_08641_));
 OA211x2_ASAP7_75t_R _26889_ (.A1(net299),
    .A2(_08640_),
    .B(_08641_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_08642_));
 INVx1_ASAP7_75t_R _26890_ (.A(_01671_),
    .Y(_08643_));
 NAND2x1_ASAP7_75t_R _26891_ (.A(net299),
    .B(_01669_),
    .Y(_08644_));
 OA211x2_ASAP7_75t_R _26892_ (.A1(net299),
    .A2(_08643_),
    .B(_08644_),
    .C(_17600_),
    .Y(_08645_));
 OR3x1_ASAP7_75t_R _26893_ (.A(_08637_),
    .B(_08642_),
    .C(_08645_),
    .Y(_08646_));
 INVx1_ASAP7_75t_R _26894_ (.A(_01664_),
    .Y(_08647_));
 NAND2x1_ASAP7_75t_R _26895_ (.A(_02290_),
    .B(_01662_),
    .Y(_08648_));
 OA211x2_ASAP7_75t_R _26896_ (.A1(_02290_),
    .A2(_08647_),
    .B(_08648_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_08649_));
 INVx1_ASAP7_75t_R _26897_ (.A(_01663_),
    .Y(_08650_));
 NAND2x1_ASAP7_75t_R _26898_ (.A(net299),
    .B(_01661_),
    .Y(_08651_));
 OA211x2_ASAP7_75t_R _26899_ (.A1(net299),
    .A2(_08650_),
    .B(_08651_),
    .C(_17600_),
    .Y(_08652_));
 OR3x1_ASAP7_75t_R _26900_ (.A(_08629_),
    .B(_08649_),
    .C(_08652_),
    .Y(_08653_));
 AND3x1_ASAP7_75t_R _26901_ (.A(_02293_),
    .B(_08646_),
    .C(_08653_),
    .Y(_08654_));
 INVx1_ASAP7_75t_R _26902_ (.A(_08654_),
    .Y(_08655_));
 TAPCELL_ASAP7_75t_R TAP_689 ();
 NOR2x1_ASAP7_75t_R _26904_ (.A(_02291_),
    .B(_05750_),
    .Y(_08657_));
 XNOR2x2_ASAP7_75t_R _26905_ (.A(_01318_),
    .B(_08657_),
    .Y(_08658_));
 AO21x1_ASAP7_75t_R _26906_ (.A1(_08639_),
    .A2(_08655_),
    .B(_08658_),
    .Y(_08659_));
 INVx1_ASAP7_75t_R _26907_ (.A(_02293_),
    .Y(_08660_));
 TAPCELL_ASAP7_75t_R TAP_688 ();
 INVx1_ASAP7_75t_R _26909_ (.A(_01660_),
    .Y(_08662_));
 NAND2x1_ASAP7_75t_R _26910_ (.A(net299),
    .B(_01658_),
    .Y(_08663_));
 OA211x2_ASAP7_75t_R _26911_ (.A1(net299),
    .A2(_08662_),
    .B(_08663_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_08664_));
 INVx1_ASAP7_75t_R _26912_ (.A(_01659_),
    .Y(_08665_));
 NAND2x1_ASAP7_75t_R _26913_ (.A(net299),
    .B(_01657_),
    .Y(_08666_));
 OA211x2_ASAP7_75t_R _26914_ (.A1(net299),
    .A2(_08665_),
    .B(_08666_),
    .C(_17600_),
    .Y(_08667_));
 OR3x1_ASAP7_75t_R _26915_ (.A(_08637_),
    .B(_08664_),
    .C(_08667_),
    .Y(_08668_));
 INVx1_ASAP7_75t_R _26916_ (.A(_01652_),
    .Y(_08669_));
 NAND2x1_ASAP7_75t_R _26917_ (.A(_02290_),
    .B(_01650_),
    .Y(_08670_));
 OA211x2_ASAP7_75t_R _26918_ (.A1(_02290_),
    .A2(_08669_),
    .B(_08670_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_08671_));
 INVx1_ASAP7_75t_R _26919_ (.A(_01651_),
    .Y(_08672_));
 NAND2x1_ASAP7_75t_R _26920_ (.A(_02290_),
    .B(_01649_),
    .Y(_08673_));
 OA211x2_ASAP7_75t_R _26921_ (.A1(_02290_),
    .A2(_08672_),
    .B(_08673_),
    .C(_17600_),
    .Y(_08674_));
 OR3x1_ASAP7_75t_R _26922_ (.A(_08629_),
    .B(_08671_),
    .C(_08674_),
    .Y(_08675_));
 AND3x1_ASAP7_75t_R _26923_ (.A(_08660_),
    .B(_08668_),
    .C(_08675_),
    .Y(_08676_));
 INVx1_ASAP7_75t_R _26924_ (.A(_01645_),
    .Y(_08677_));
 NOR2x1_ASAP7_75t_R _26925_ (.A(_02290_),
    .B(_01647_),
    .Y(_08678_));
 AO21x1_ASAP7_75t_R _26926_ (.A1(_02290_),
    .A2(_08677_),
    .B(_08678_),
    .Y(_08679_));
 INVx1_ASAP7_75t_R _26927_ (.A(_01648_),
    .Y(_08680_));
 NAND2x1_ASAP7_75t_R _26928_ (.A(_02290_),
    .B(_01646_),
    .Y(_08681_));
 OA211x2_ASAP7_75t_R _26929_ (.A1(_02290_),
    .A2(_08680_),
    .B(_08681_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_08682_));
 AO21x1_ASAP7_75t_R _26930_ (.A1(_17600_),
    .A2(_08679_),
    .B(_08682_),
    .Y(_08683_));
 INVx1_ASAP7_75t_R _26931_ (.A(_01654_),
    .Y(_08684_));
 NAND2x1_ASAP7_75t_R _26932_ (.A(_08621_),
    .B(_01656_),
    .Y(_08685_));
 OA211x2_ASAP7_75t_R _26933_ (.A1(_08621_),
    .A2(_08684_),
    .B(_08685_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_08686_));
 INVx1_ASAP7_75t_R _26934_ (.A(_01655_),
    .Y(_08687_));
 NAND2x1_ASAP7_75t_R _26935_ (.A(_02290_),
    .B(_01653_),
    .Y(_08688_));
 OA211x2_ASAP7_75t_R _26936_ (.A1(_02290_),
    .A2(_08687_),
    .B(_08688_),
    .C(_17600_),
    .Y(_08689_));
 OR3x1_ASAP7_75t_R _26937_ (.A(_08637_),
    .B(_08686_),
    .C(_08689_),
    .Y(_08690_));
 OA211x2_ASAP7_75t_R _26938_ (.A1(_08629_),
    .A2(_08683_),
    .B(_08690_),
    .C(_02293_),
    .Y(_08691_));
 OAI21x1_ASAP7_75t_R _26939_ (.A1(_08676_),
    .A2(_08691_),
    .B(_08658_),
    .Y(_08692_));
 TAPCELL_ASAP7_75t_R TAP_687 ();
 AO21x1_ASAP7_75t_R _26941_ (.A1(_08659_),
    .A2(_08692_),
    .B(_01357_),
    .Y(_08694_));
 AND3x4_ASAP7_75t_R _26942_ (.A(_13317_),
    .B(_05743_),
    .C(_08576_),
    .Y(_08695_));
 TAPCELL_ASAP7_75t_R TAP_686 ();
 NAND2x1_ASAP7_75t_R _26944_ (.A(_13530_),
    .B(net280),
    .Y(_08697_));
 OA211x2_ASAP7_75t_R _26945_ (.A1(_01645_),
    .A2(_01873_),
    .B(_08695_),
    .C(_08697_),
    .Y(_08698_));
 OA211x2_ASAP7_75t_R _26946_ (.A1(_08609_),
    .A2(_08618_),
    .B(_08694_),
    .C(_08698_),
    .Y(_08699_));
 OR3x1_ASAP7_75t_R _26947_ (.A(_08590_),
    .B(_08604_),
    .C(_08699_),
    .Y(_08700_));
 OAI21x1_ASAP7_75t_R _26948_ (.A1(_00324_),
    .A2(_08591_),
    .B(_08700_),
    .Y(_02688_));
 AND2x2_ASAP7_75t_R _26949_ (.A(_00291_),
    .B(_07079_),
    .Y(_08701_));
 AO21x1_ASAP7_75t_R _26950_ (.A1(_01360_),
    .A2(_07077_),
    .B(_08701_),
    .Y(_08702_));
 NOR2x1_ASAP7_75t_R _26951_ (.A(_13523_),
    .B(_08600_),
    .Y(_08703_));
 AO21x1_ASAP7_75t_R _26952_ (.A1(_07076_),
    .A2(_08702_),
    .B(_08703_),
    .Y(_08704_));
 TAPCELL_ASAP7_75t_R TAP_685 ();
 TAPCELL_ASAP7_75t_R TAP_684 ();
 TAPCELL_ASAP7_75t_R TAP_683 ();
 OR3x1_ASAP7_75t_R _26956_ (.A(_05750_),
    .B(_05752_),
    .C(_08607_),
    .Y(_08708_));
 AND2x2_ASAP7_75t_R _26957_ (.A(_16499_),
    .B(_08614_),
    .Y(_08709_));
 AO21x1_ASAP7_75t_R _26958_ (.A1(_00291_),
    .A2(_08607_),
    .B(_08709_),
    .Y(_08710_));
 AO32x1_ASAP7_75t_R _26959_ (.A1(_01324_),
    .A2(_08598_),
    .A3(_08708_),
    .B1(_08710_),
    .B2(_08610_),
    .Y(_08711_));
 TAPCELL_ASAP7_75t_R TAP_682 ();
 TAPCELL_ASAP7_75t_R TAP_681 ();
 OA21x2_ASAP7_75t_R _26962_ (.A1(_00285_),
    .A2(_16499_),
    .B(_08695_),
    .Y(_08714_));
 OA21x2_ASAP7_75t_R _26963_ (.A1(_01357_),
    .A2(_08617_),
    .B(_08714_),
    .Y(_08715_));
 OA21x2_ASAP7_75t_R _26964_ (.A1(_01727_),
    .A2(_08711_),
    .B(_08715_),
    .Y(_08716_));
 OR3x1_ASAP7_75t_R _26965_ (.A(_08590_),
    .B(_08704_),
    .C(_08716_),
    .Y(_08717_));
 OAI21x1_ASAP7_75t_R _26966_ (.A1(_00291_),
    .A2(_08591_),
    .B(_08717_),
    .Y(_02689_));
 AND2x2_ASAP7_75t_R _26967_ (.A(_00663_),
    .B(_07079_),
    .Y(_08718_));
 AO21x1_ASAP7_75t_R _26968_ (.A1(_01364_),
    .A2(_07077_),
    .B(_08718_),
    .Y(_08719_));
 NOR2x1_ASAP7_75t_R _26969_ (.A(_14684_),
    .B(_08600_),
    .Y(_08720_));
 AO21x1_ASAP7_75t_R _26970_ (.A1(_07076_),
    .A2(_08719_),
    .B(_08720_),
    .Y(_08721_));
 OA211x2_ASAP7_75t_R _26971_ (.A1(_01326_),
    .A2(_08608_),
    .B(_08598_),
    .C(_01325_),
    .Y(_08722_));
 TAPCELL_ASAP7_75t_R TAP_680 ();
 TAPCELL_ASAP7_75t_R TAP_679 ();
 AND2x2_ASAP7_75t_R _26974_ (.A(_05767_),
    .B(_08614_),
    .Y(_08725_));
 AO21x1_ASAP7_75t_R _26975_ (.A1(_00663_),
    .A2(_08607_),
    .B(_08725_),
    .Y(_08726_));
 AO21x1_ASAP7_75t_R _26976_ (.A1(_08610_),
    .A2(_08726_),
    .B(_01727_),
    .Y(_08727_));
 OA21x2_ASAP7_75t_R _26977_ (.A1(_00285_),
    .A2(_05767_),
    .B(_08695_),
    .Y(_08728_));
 OA21x2_ASAP7_75t_R _26978_ (.A1(_01357_),
    .A2(_08710_),
    .B(_08728_),
    .Y(_08729_));
 OA21x2_ASAP7_75t_R _26979_ (.A1(_08722_),
    .A2(_08727_),
    .B(_08729_),
    .Y(_08730_));
 OR3x1_ASAP7_75t_R _26980_ (.A(_08590_),
    .B(_08721_),
    .C(_08730_),
    .Y(_08731_));
 OAI21x1_ASAP7_75t_R _26981_ (.A1(_00663_),
    .A2(_08591_),
    .B(_08731_),
    .Y(_02690_));
 TAPCELL_ASAP7_75t_R TAP_678 ();
 NAND2x1_ASAP7_75t_R _26983_ (.A(_02231_),
    .B(_07077_),
    .Y(_08733_));
 OA211x2_ASAP7_75t_R _26984_ (.A1(_00665_),
    .A2(_07077_),
    .B(_08733_),
    .C(_07076_),
    .Y(_08734_));
 NOR2x1_ASAP7_75t_R _26985_ (.A(_14752_),
    .B(_08600_),
    .Y(_08735_));
 AND2x2_ASAP7_75t_R _26986_ (.A(_06277_),
    .B(_08614_),
    .Y(_08736_));
 AO21x1_ASAP7_75t_R _26987_ (.A1(_00665_),
    .A2(_08607_),
    .B(_08736_),
    .Y(_08737_));
 AND3x4_ASAP7_75t_R _26988_ (.A(_13325_),
    .B(_00282_),
    .C(_13576_),
    .Y(_08738_));
 OA211x2_ASAP7_75t_R _26989_ (.A1(_01320_),
    .A2(_08608_),
    .B(_08738_),
    .C(_01327_),
    .Y(_08739_));
 AO21x1_ASAP7_75t_R _26990_ (.A1(_08610_),
    .A2(_08737_),
    .B(_08739_),
    .Y(_08740_));
 TAPCELL_ASAP7_75t_R TAP_677 ();
 OA21x2_ASAP7_75t_R _26992_ (.A1(_00285_),
    .A2(_06277_),
    .B(_08695_),
    .Y(_08742_));
 OA21x2_ASAP7_75t_R _26993_ (.A1(_01357_),
    .A2(_08726_),
    .B(_08742_),
    .Y(_08743_));
 OA21x2_ASAP7_75t_R _26994_ (.A1(_01727_),
    .A2(_08740_),
    .B(_08743_),
    .Y(_08744_));
 OR4x1_ASAP7_75t_R _26995_ (.A(_08590_),
    .B(_08734_),
    .C(_08735_),
    .D(_08744_),
    .Y(_08745_));
 OAI21x1_ASAP7_75t_R _26996_ (.A1(_00665_),
    .A2(_08591_),
    .B(_08745_),
    .Y(_02691_));
 INVx3_ASAP7_75t_R _26997_ (.A(_01322_),
    .Y(_08746_));
 INVx1_ASAP7_75t_R _26998_ (.A(_17607_),
    .Y(_08747_));
 NAND2x2_ASAP7_75t_R _26999_ (.A(_08747_),
    .B(_08614_),
    .Y(_08748_));
 TAPCELL_ASAP7_75t_R TAP_676 ();
 OR3x4_ASAP7_75t_R _27001_ (.A(_05751_),
    .B(_08746_),
    .C(_08748_),
    .Y(_08750_));
 OA211x2_ASAP7_75t_R _27002_ (.A1(_01321_),
    .A2(_08750_),
    .B(_08598_),
    .C(_01328_),
    .Y(_08751_));
 TAPCELL_ASAP7_75t_R TAP_675 ();
 TAPCELL_ASAP7_75t_R TAP_674 ();
 TAPCELL_ASAP7_75t_R TAP_673 ();
 AND2x2_ASAP7_75t_R _27006_ (.A(_05766_),
    .B(_08614_),
    .Y(_08755_));
 AO21x1_ASAP7_75t_R _27007_ (.A1(_00668_),
    .A2(_08607_),
    .B(_08755_),
    .Y(_08756_));
 AO21x1_ASAP7_75t_R _27008_ (.A1(_08610_),
    .A2(_08756_),
    .B(_01727_),
    .Y(_08757_));
 TAPCELL_ASAP7_75t_R TAP_672 ();
 OA21x2_ASAP7_75t_R _27010_ (.A1(_00285_),
    .A2(_05766_),
    .B(_08695_),
    .Y(_08759_));
 OA21x2_ASAP7_75t_R _27011_ (.A1(_01357_),
    .A2(_08737_),
    .B(_08759_),
    .Y(_08760_));
 OAI21x1_ASAP7_75t_R _27012_ (.A1(_08751_),
    .A2(_08757_),
    .B(_08760_),
    .Y(_08761_));
 NAND2x1_ASAP7_75t_R _27013_ (.A(_00668_),
    .B(_07079_),
    .Y(_08762_));
 NAND2x1_ASAP7_75t_R _27014_ (.A(_01376_),
    .B(_07077_),
    .Y(_08763_));
 AO21x1_ASAP7_75t_R _27015_ (.A1(_08762_),
    .A2(_08763_),
    .B(_05745_),
    .Y(_08764_));
 OA211x2_ASAP7_75t_R _27016_ (.A1(_14820_),
    .A2(_08600_),
    .B(_08764_),
    .C(_08591_),
    .Y(_08765_));
 AO22x1_ASAP7_75t_R _27017_ (.A1(_06699_),
    .A2(_08590_),
    .B1(_08761_),
    .B2(_08765_),
    .Y(_02692_));
 TAPCELL_ASAP7_75t_R TAP_671 ();
 INVx1_ASAP7_75t_R _27019_ (.A(net176),
    .Y(_08767_));
 OA21x2_ASAP7_75t_R _27020_ (.A1(_00285_),
    .A2(_08767_),
    .B(_08695_),
    .Y(_08768_));
 OAI21x1_ASAP7_75t_R _27021_ (.A1(_01357_),
    .A2(_08756_),
    .B(_08768_),
    .Y(_08769_));
 AND2x2_ASAP7_75t_R _27022_ (.A(_08767_),
    .B(_08614_),
    .Y(_08770_));
 AO21x1_ASAP7_75t_R _27023_ (.A1(_00670_),
    .A2(_08607_),
    .B(_08770_),
    .Y(_08771_));
 OR3x1_ASAP7_75t_R _27024_ (.A(_08746_),
    .B(_05752_),
    .C(_08748_),
    .Y(_08772_));
 AND3x1_ASAP7_75t_R _27025_ (.A(_01329_),
    .B(_08598_),
    .C(_08772_),
    .Y(_08773_));
 AOI211x1_ASAP7_75t_R _27026_ (.A1(_08610_),
    .A2(_08771_),
    .B(_08773_),
    .C(_01727_),
    .Y(_08774_));
 AND2x2_ASAP7_75t_R _27027_ (.A(_07077_),
    .B(_07561_),
    .Y(_08775_));
 AOI21x1_ASAP7_75t_R _27028_ (.A1(_00670_),
    .A2(_07079_),
    .B(_08775_),
    .Y(_08776_));
 OA222x2_ASAP7_75t_R _27029_ (.A1(_14873_),
    .A2(_08600_),
    .B1(_08769_),
    .B2(_08774_),
    .C1(_08776_),
    .C2(_05745_),
    .Y(_08777_));
 NAND2x1_ASAP7_75t_R _27030_ (.A(_00670_),
    .B(_08590_),
    .Y(_08778_));
 OA21x2_ASAP7_75t_R _27031_ (.A1(_08590_),
    .A2(_08777_),
    .B(_08778_),
    .Y(_02693_));
 OR2x2_ASAP7_75t_R _27032_ (.A(_07079_),
    .B(_08590_),
    .Y(_08779_));
 AO32x1_ASAP7_75t_R _27033_ (.A1(_07598_),
    .A2(_14626_),
    .A3(_07078_),
    .B1(_08779_),
    .B2(_00672_),
    .Y(_08780_));
 AND2x2_ASAP7_75t_R _27034_ (.A(_05768_),
    .B(_08614_),
    .Y(_08781_));
 AO21x1_ASAP7_75t_R _27035_ (.A1(_00672_),
    .A2(_08607_),
    .B(_08781_),
    .Y(_08782_));
 TAPCELL_ASAP7_75t_R TAP_670 ();
 OA211x2_ASAP7_75t_R _27037_ (.A1(_01326_),
    .A2(_08750_),
    .B(_08738_),
    .C(_01330_),
    .Y(_08784_));
 AO21x1_ASAP7_75t_R _27038_ (.A1(_08610_),
    .A2(_08782_),
    .B(_08784_),
    .Y(_08785_));
 AND3x4_ASAP7_75t_R _27039_ (.A(_14626_),
    .B(_05745_),
    .C(_08589_),
    .Y(_08786_));
 TAPCELL_ASAP7_75t_R TAP_669 ();
 OR2x6_ASAP7_75t_R _27041_ (.A(_08576_),
    .B(_08598_),
    .Y(_08788_));
 TAPCELL_ASAP7_75t_R TAP_668 ();
 OAI22x1_ASAP7_75t_R _27043_ (.A1(_00285_),
    .A2(_05768_),
    .B1(_08771_),
    .B2(_01357_),
    .Y(_08790_));
 AND2x4_ASAP7_75t_R _27044_ (.A(_01873_),
    .B(_13527_),
    .Y(_08791_));
 OAI22x1_ASAP7_75t_R _27045_ (.A1(_14936_),
    .A2(_08788_),
    .B1(_08790_),
    .B2(_08791_),
    .Y(_08792_));
 OA211x2_ASAP7_75t_R _27046_ (.A1(_01727_),
    .A2(_08785_),
    .B(_08786_),
    .C(_08792_),
    .Y(_08793_));
 NOR2x1_ASAP7_75t_R _27047_ (.A(_08780_),
    .B(_08793_),
    .Y(_02694_));
 OA211x2_ASAP7_75t_R _27048_ (.A1(_01320_),
    .A2(_08750_),
    .B(_08598_),
    .C(_01331_),
    .Y(_08794_));
 AND2x2_ASAP7_75t_R _27049_ (.A(_00674_),
    .B(_08607_),
    .Y(_08795_));
 AO21x1_ASAP7_75t_R _27050_ (.A1(_00676_),
    .A2(_08614_),
    .B(_08795_),
    .Y(_08796_));
 AO21x1_ASAP7_75t_R _27051_ (.A1(_08610_),
    .A2(_08796_),
    .B(_01727_),
    .Y(_08797_));
 OA21x2_ASAP7_75t_R _27052_ (.A1(_00285_),
    .A2(_00676_),
    .B(_08695_),
    .Y(_08798_));
 OA21x2_ASAP7_75t_R _27053_ (.A1(_01357_),
    .A2(_08782_),
    .B(_08798_),
    .Y(_08799_));
 OA21x2_ASAP7_75t_R _27054_ (.A1(_08794_),
    .A2(_08797_),
    .B(_08799_),
    .Y(_08800_));
 NOR2x2_ASAP7_75t_R _27055_ (.A(_08576_),
    .B(_08598_),
    .Y(_08801_));
 AND2x2_ASAP7_75t_R _27056_ (.A(_05745_),
    .B(_08801_),
    .Y(_08802_));
 AO21x1_ASAP7_75t_R _27057_ (.A1(_06710_),
    .A2(_08802_),
    .B(_07653_),
    .Y(_08803_));
 OR3x1_ASAP7_75t_R _27058_ (.A(_08590_),
    .B(_08800_),
    .C(_08803_),
    .Y(_08804_));
 OAI21x1_ASAP7_75t_R _27059_ (.A1(_00674_),
    .A2(_08591_),
    .B(_08804_),
    .Y(_02695_));
 AND2x2_ASAP7_75t_R _27060_ (.A(_05773_),
    .B(_08614_),
    .Y(_08805_));
 AO21x1_ASAP7_75t_R _27061_ (.A1(_00677_),
    .A2(_08607_),
    .B(_08805_),
    .Y(_08806_));
 NAND2x2_ASAP7_75t_R _27062_ (.A(_01318_),
    .B(_08746_),
    .Y(_08807_));
 OR3x4_ASAP7_75t_R _27063_ (.A(_08747_),
    .B(_08607_),
    .C(_08807_),
    .Y(_08808_));
 OA211x2_ASAP7_75t_R _27064_ (.A1(_01321_),
    .A2(_08808_),
    .B(_08598_),
    .C(_01332_),
    .Y(_08809_));
 AO21x1_ASAP7_75t_R _27065_ (.A1(_08610_),
    .A2(_08806_),
    .B(_08809_),
    .Y(_08810_));
 OA21x2_ASAP7_75t_R _27066_ (.A1(_00285_),
    .A2(_05773_),
    .B(_08695_),
    .Y(_08811_));
 OA211x2_ASAP7_75t_R _27067_ (.A1(_01357_),
    .A2(_08796_),
    .B(_08811_),
    .C(_08591_),
    .Y(_08812_));
 OAI21x1_ASAP7_75t_R _27068_ (.A1(_01727_),
    .A2(_08810_),
    .B(_08812_),
    .Y(_08813_));
 INVx1_ASAP7_75t_R _27069_ (.A(_14626_),
    .Y(_08814_));
 OA33x2_ASAP7_75t_R _27070_ (.A1(_02235_),
    .A2(_08814_),
    .A3(_07437_),
    .B1(_08590_),
    .B2(_08600_),
    .B3(_15042_),
    .Y(_08815_));
 NAND2x1_ASAP7_75t_R _27071_ (.A(_00677_),
    .B(_08779_),
    .Y(_08816_));
 AND3x1_ASAP7_75t_R _27072_ (.A(_08813_),
    .B(_08815_),
    .C(_08816_),
    .Y(_02696_));
 AND2x2_ASAP7_75t_R _27073_ (.A(_06350_),
    .B(_08614_),
    .Y(_08817_));
 AO21x1_ASAP7_75t_R _27074_ (.A1(_00680_),
    .A2(_08607_),
    .B(_08817_),
    .Y(_08818_));
 NAND2x2_ASAP7_75t_R _27075_ (.A(_17607_),
    .B(_08614_),
    .Y(_08819_));
 OR3x1_ASAP7_75t_R _27076_ (.A(_01322_),
    .B(_05752_),
    .C(_08819_),
    .Y(_08820_));
 AND2x2_ASAP7_75t_R _27077_ (.A(_01333_),
    .B(_08738_),
    .Y(_08821_));
 AO221x1_ASAP7_75t_R _27078_ (.A1(_08610_),
    .A2(_08818_),
    .B1(_08820_),
    .B2(_08821_),
    .C(_01727_),
    .Y(_08822_));
 OA21x2_ASAP7_75t_R _27079_ (.A1(_00285_),
    .A2(_06350_),
    .B(_08695_),
    .Y(_08823_));
 OA211x2_ASAP7_75t_R _27080_ (.A1(_01357_),
    .A2(_08806_),
    .B(_08822_),
    .C(_08823_),
    .Y(_08824_));
 AND2x2_ASAP7_75t_R _27081_ (.A(_07077_),
    .B(_07759_),
    .Y(_08825_));
 AO21x1_ASAP7_75t_R _27082_ (.A1(_00680_),
    .A2(_07079_),
    .B(_08825_),
    .Y(_08826_));
 NOR2x1_ASAP7_75t_R _27083_ (.A(_15096_),
    .B(_08600_),
    .Y(_08827_));
 AO21x1_ASAP7_75t_R _27084_ (.A1(_07076_),
    .A2(_08826_),
    .B(_08827_),
    .Y(_08828_));
 OR3x1_ASAP7_75t_R _27085_ (.A(_08590_),
    .B(_08824_),
    .C(_08828_),
    .Y(_08829_));
 OAI21x1_ASAP7_75t_R _27086_ (.A1(_00680_),
    .A2(_08591_),
    .B(_08829_),
    .Y(_02697_));
 AND2x2_ASAP7_75t_R _27087_ (.A(_05772_),
    .B(_08614_),
    .Y(_08830_));
 AO21x1_ASAP7_75t_R _27088_ (.A1(_00682_),
    .A2(_08607_),
    .B(_08830_),
    .Y(_08831_));
 OA211x2_ASAP7_75t_R _27089_ (.A1(_01326_),
    .A2(_08808_),
    .B(_08738_),
    .C(_01334_),
    .Y(_08832_));
 AO21x1_ASAP7_75t_R _27090_ (.A1(_08610_),
    .A2(_08831_),
    .B(_08832_),
    .Y(_08833_));
 OA21x2_ASAP7_75t_R _27091_ (.A1(_00285_),
    .A2(_05772_),
    .B(_08695_),
    .Y(_08834_));
 OA21x2_ASAP7_75t_R _27092_ (.A1(_01357_),
    .A2(_08818_),
    .B(_08834_),
    .Y(_08835_));
 OA21x2_ASAP7_75t_R _27093_ (.A1(_01727_),
    .A2(_08833_),
    .B(_08835_),
    .Y(_08836_));
 OR2x2_ASAP7_75t_R _27094_ (.A(_00682_),
    .B(_07077_),
    .Y(_08837_));
 OA211x2_ASAP7_75t_R _27095_ (.A1(_07790_),
    .A2(_07079_),
    .B(_08837_),
    .C(_07076_),
    .Y(_08838_));
 NOR2x1_ASAP7_75t_R _27096_ (.A(_15157_),
    .B(_08600_),
    .Y(_08839_));
 OR5x1_ASAP7_75t_R _27097_ (.A(_13318_),
    .B(_08590_),
    .C(_08836_),
    .D(_08838_),
    .E(_08839_),
    .Y(_08840_));
 OAI21x1_ASAP7_75t_R _27098_ (.A1(_00682_),
    .A2(_08591_),
    .B(_08840_),
    .Y(_02698_));
 AND2x2_ASAP7_75t_R _27099_ (.A(_06368_),
    .B(_08614_),
    .Y(_08841_));
 AO21x1_ASAP7_75t_R _27100_ (.A1(_00684_),
    .A2(_08607_),
    .B(_08841_),
    .Y(_08842_));
 OA211x2_ASAP7_75t_R _27101_ (.A1(_01320_),
    .A2(_08808_),
    .B(_08738_),
    .C(_01335_),
    .Y(_08843_));
 AO21x1_ASAP7_75t_R _27102_ (.A1(_08610_),
    .A2(_08842_),
    .B(_08843_),
    .Y(_08844_));
 OA21x2_ASAP7_75t_R _27103_ (.A1(_00285_),
    .A2(_06368_),
    .B(_08695_),
    .Y(_08845_));
 OA21x2_ASAP7_75t_R _27104_ (.A1(_01357_),
    .A2(_08831_),
    .B(_08845_),
    .Y(_08846_));
 OA21x2_ASAP7_75t_R _27105_ (.A1(_01727_),
    .A2(_08844_),
    .B(_08846_),
    .Y(_08847_));
 NOR2x1_ASAP7_75t_R _27106_ (.A(_14574_),
    .B(_08600_),
    .Y(_08848_));
 OR4x1_ASAP7_75t_R _27107_ (.A(_07827_),
    .B(_08590_),
    .C(_08847_),
    .D(_08848_),
    .Y(_08849_));
 OAI21x1_ASAP7_75t_R _27108_ (.A1(_00684_),
    .A2(_08591_),
    .B(_08849_),
    .Y(_02699_));
 AO32x1_ASAP7_75t_R _27109_ (.A1(_07872_),
    .A2(_14626_),
    .A3(_07078_),
    .B1(_08779_),
    .B2(_00686_),
    .Y(_08850_));
 AND2x2_ASAP7_75t_R _27110_ (.A(_05771_),
    .B(_08614_),
    .Y(_08851_));
 AO21x1_ASAP7_75t_R _27111_ (.A1(_00686_),
    .A2(_08607_),
    .B(_08851_),
    .Y(_08852_));
 OR3x1_ASAP7_75t_R _27112_ (.A(_01321_),
    .B(_08748_),
    .C(_08807_),
    .Y(_08853_));
 AND3x1_ASAP7_75t_R _27113_ (.A(_01336_),
    .B(_08738_),
    .C(_08853_),
    .Y(_08854_));
 AO21x1_ASAP7_75t_R _27114_ (.A1(_08610_),
    .A2(_08852_),
    .B(_08854_),
    .Y(_08855_));
 OA21x2_ASAP7_75t_R _27115_ (.A1(_00285_),
    .A2(_05771_),
    .B(_08576_),
    .Y(_08856_));
 OA21x2_ASAP7_75t_R _27116_ (.A1(_01357_),
    .A2(_08842_),
    .B(_08856_),
    .Y(_08857_));
 AO21x1_ASAP7_75t_R _27117_ (.A1(_13878_),
    .A2(_08801_),
    .B(_08857_),
    .Y(_08858_));
 OA211x2_ASAP7_75t_R _27118_ (.A1(_01727_),
    .A2(_08855_),
    .B(_08858_),
    .C(_08786_),
    .Y(_08859_));
 NOR2x1_ASAP7_75t_R _27119_ (.A(_08850_),
    .B(_08859_),
    .Y(_02700_));
 OR3x1_ASAP7_75t_R _27120_ (.A(_01322_),
    .B(_05752_),
    .C(_08748_),
    .Y(_08860_));
 AND3x4_ASAP7_75t_R _27121_ (.A(_00282_),
    .B(_13317_),
    .C(_05743_),
    .Y(_08861_));
 AND2x2_ASAP7_75t_R _27122_ (.A(_06384_),
    .B(_08614_),
    .Y(_08862_));
 AO21x1_ASAP7_75t_R _27123_ (.A1(_00718_),
    .A2(_08607_),
    .B(_08862_),
    .Y(_08863_));
 AO32x1_ASAP7_75t_R _27124_ (.A1(_01337_),
    .A2(_08860_),
    .A3(_08861_),
    .B1(_08610_),
    .B2(_08863_),
    .Y(_08864_));
 OA21x2_ASAP7_75t_R _27125_ (.A1(_00285_),
    .A2(_06384_),
    .B(_08695_),
    .Y(_08865_));
 OA21x2_ASAP7_75t_R _27126_ (.A1(_01357_),
    .A2(_08852_),
    .B(_08865_),
    .Y(_08866_));
 OA21x2_ASAP7_75t_R _27127_ (.A1(_01727_),
    .A2(_08864_),
    .B(_08866_),
    .Y(_08867_));
 NOR2x1_ASAP7_75t_R _27128_ (.A(_15401_),
    .B(_08600_),
    .Y(_08868_));
 OR4x1_ASAP7_75t_R _27129_ (.A(_07920_),
    .B(_08590_),
    .C(_08867_),
    .D(_08868_),
    .Y(_08869_));
 OAI21x1_ASAP7_75t_R _27130_ (.A1(_00718_),
    .A2(_08591_),
    .B(_08869_),
    .Y(_02701_));
 NAND2x1_ASAP7_75t_R _27131_ (.A(_06787_),
    .B(_07079_),
    .Y(_08870_));
 NAND2x1_ASAP7_75t_R _27132_ (.A(_02241_),
    .B(_07077_),
    .Y(_08871_));
 AO32x1_ASAP7_75t_R _27133_ (.A1(_07076_),
    .A2(_08870_),
    .A3(_08871_),
    .B1(_08802_),
    .B2(_15555_),
    .Y(_08872_));
 OR3x4_ASAP7_75t_R _27134_ (.A(_17607_),
    .B(_08607_),
    .C(_08807_),
    .Y(_08873_));
 OA211x2_ASAP7_75t_R _27135_ (.A1(_01326_),
    .A2(_08873_),
    .B(_08861_),
    .C(_01338_),
    .Y(_08874_));
 AND2x2_ASAP7_75t_R _27136_ (.A(_15557_),
    .B(_08614_),
    .Y(_08875_));
 AO21x1_ASAP7_75t_R _27137_ (.A1(_00750_),
    .A2(_08607_),
    .B(_08875_),
    .Y(_08876_));
 AO21x1_ASAP7_75t_R _27138_ (.A1(_08610_),
    .A2(_08876_),
    .B(_01727_),
    .Y(_08877_));
 OA21x2_ASAP7_75t_R _27139_ (.A1(_00285_),
    .A2(_15557_),
    .B(_08695_),
    .Y(_08878_));
 OA21x2_ASAP7_75t_R _27140_ (.A1(_01357_),
    .A2(_08863_),
    .B(_08878_),
    .Y(_08879_));
 OA21x2_ASAP7_75t_R _27141_ (.A1(_08874_),
    .A2(_08877_),
    .B(_08879_),
    .Y(_08880_));
 OR3x1_ASAP7_75t_R _27142_ (.A(_08590_),
    .B(_08872_),
    .C(_08880_),
    .Y(_08881_));
 OAI21x1_ASAP7_75t_R _27143_ (.A1(_00750_),
    .A2(_08591_),
    .B(_08881_),
    .Y(_02702_));
 OA211x2_ASAP7_75t_R _27144_ (.A1(_01320_),
    .A2(_08873_),
    .B(_08738_),
    .C(_01339_),
    .Y(_08882_));
 AND2x2_ASAP7_75t_R _27145_ (.A(_00783_),
    .B(_08607_),
    .Y(_08883_));
 AO21x1_ASAP7_75t_R _27146_ (.A1(_00785_),
    .A2(_08614_),
    .B(_08883_),
    .Y(_08884_));
 AO21x1_ASAP7_75t_R _27147_ (.A1(_08610_),
    .A2(_08884_),
    .B(_01727_),
    .Y(_08885_));
 OA21x2_ASAP7_75t_R _27148_ (.A1(_00285_),
    .A2(_00785_),
    .B(_08695_),
    .Y(_08886_));
 OA21x2_ASAP7_75t_R _27149_ (.A1(_01357_),
    .A2(_08876_),
    .B(_08886_),
    .Y(_08887_));
 OAI21x1_ASAP7_75t_R _27150_ (.A1(_08882_),
    .A2(_08885_),
    .B(_08887_),
    .Y(_08888_));
 OA211x2_ASAP7_75t_R _27151_ (.A1(_15665_),
    .A2(_08600_),
    .B(_08004_),
    .C(_13576_),
    .Y(_08889_));
 AND3x1_ASAP7_75t_R _27152_ (.A(_08591_),
    .B(_08888_),
    .C(_08889_),
    .Y(_08890_));
 AO21x1_ASAP7_75t_R _27153_ (.A1(_06789_),
    .A2(_08590_),
    .B(_08890_),
    .Y(_02703_));
 NAND2x1_ASAP7_75t_R _27154_ (.A(_00816_),
    .B(_08590_),
    .Y(_08891_));
 AND2x2_ASAP7_75t_R _27155_ (.A(_05770_),
    .B(_08614_),
    .Y(_08892_));
 AO21x1_ASAP7_75t_R _27156_ (.A1(_00816_),
    .A2(_08607_),
    .B(_08892_),
    .Y(_08893_));
 OR3x4_ASAP7_75t_R _27157_ (.A(_01318_),
    .B(_05750_),
    .C(_08607_),
    .Y(_08894_));
 OA211x2_ASAP7_75t_R _27158_ (.A1(_01321_),
    .A2(_08894_),
    .B(_08861_),
    .C(_01340_),
    .Y(_08895_));
 AOI211x1_ASAP7_75t_R _27159_ (.A1(_08610_),
    .A2(_08893_),
    .B(_08895_),
    .C(_01727_),
    .Y(_08896_));
 OA21x2_ASAP7_75t_R _27160_ (.A1(_00285_),
    .A2(_05770_),
    .B(_08576_),
    .Y(_08897_));
 OAI21x1_ASAP7_75t_R _27161_ (.A1(_01357_),
    .A2(_08884_),
    .B(_08897_),
    .Y(_08898_));
 OA21x2_ASAP7_75t_R _27162_ (.A1(_06792_),
    .A2(_08788_),
    .B(_08898_),
    .Y(_08899_));
 OR4x1_ASAP7_75t_R _27163_ (.A(_07076_),
    .B(_08590_),
    .C(_08896_),
    .D(_08899_),
    .Y(_08900_));
 OA211x2_ASAP7_75t_R _27164_ (.A1(_08052_),
    .A2(_08590_),
    .B(_08891_),
    .C(_08900_),
    .Y(_02704_));
 INVx1_ASAP7_75t_R _27165_ (.A(_00849_),
    .Y(_08901_));
 OR4x1_ASAP7_75t_R _27166_ (.A(_01319_),
    .B(_01318_),
    .C(_05750_),
    .D(_08607_),
    .Y(_08902_));
 AND2x2_ASAP7_75t_R _27167_ (.A(_06412_),
    .B(_08614_),
    .Y(_08903_));
 AO21x1_ASAP7_75t_R _27168_ (.A1(_00849_),
    .A2(_08607_),
    .B(_08903_),
    .Y(_08904_));
 AO32x1_ASAP7_75t_R _27169_ (.A1(_01341_),
    .A2(_08598_),
    .A3(_08902_),
    .B1(_08904_),
    .B2(_08610_),
    .Y(_08905_));
 OA21x2_ASAP7_75t_R _27170_ (.A1(_00285_),
    .A2(_06412_),
    .B(_08695_),
    .Y(_08906_));
 OA21x2_ASAP7_75t_R _27171_ (.A1(_01357_),
    .A2(_08893_),
    .B(_08906_),
    .Y(_08907_));
 OAI21x1_ASAP7_75t_R _27172_ (.A1(_01727_),
    .A2(_08905_),
    .B(_08907_),
    .Y(_08908_));
 OA211x2_ASAP7_75t_R _27173_ (.A1(_15890_),
    .A2(_08600_),
    .B(_08089_),
    .C(_13576_),
    .Y(_08909_));
 AND3x1_ASAP7_75t_R _27174_ (.A(_08591_),
    .B(_08908_),
    .C(_08909_),
    .Y(_08910_));
 AO21x1_ASAP7_75t_R _27175_ (.A1(_08901_),
    .A2(_08590_),
    .B(_08910_),
    .Y(_02705_));
 AND2x2_ASAP7_75t_R _27176_ (.A(_16020_),
    .B(_08614_),
    .Y(_08911_));
 AO21x1_ASAP7_75t_R _27177_ (.A1(_00881_),
    .A2(_08607_),
    .B(_08911_),
    .Y(_08912_));
 OA211x2_ASAP7_75t_R _27178_ (.A1(_01326_),
    .A2(_08894_),
    .B(_08738_),
    .C(_01342_),
    .Y(_08913_));
 AO21x1_ASAP7_75t_R _27179_ (.A1(_08610_),
    .A2(_08912_),
    .B(_08913_),
    .Y(_08914_));
 OA21x2_ASAP7_75t_R _27180_ (.A1(_00285_),
    .A2(_16020_),
    .B(_08695_),
    .Y(_08915_));
 OA21x2_ASAP7_75t_R _27181_ (.A1(_01357_),
    .A2(_08904_),
    .B(_08915_),
    .Y(_08916_));
 OA21x2_ASAP7_75t_R _27182_ (.A1(_01727_),
    .A2(_08914_),
    .B(_08916_),
    .Y(_08917_));
 AO21x1_ASAP7_75t_R _27183_ (.A1(_16018_),
    .A2(_08802_),
    .B(_08121_),
    .Y(_08918_));
 OR3x1_ASAP7_75t_R _27184_ (.A(_08590_),
    .B(_08917_),
    .C(_08918_),
    .Y(_08919_));
 OAI21x1_ASAP7_75t_R _27185_ (.A1(_00881_),
    .A2(_08591_),
    .B(_08919_),
    .Y(_02706_));
 OA211x2_ASAP7_75t_R _27186_ (.A1(_01320_),
    .A2(_08894_),
    .B(_08598_),
    .C(_01343_),
    .Y(_08920_));
 AND2x2_ASAP7_75t_R _27187_ (.A(_06426_),
    .B(_08614_),
    .Y(_08921_));
 AO21x1_ASAP7_75t_R _27188_ (.A1(_00914_),
    .A2(_08607_),
    .B(_08921_),
    .Y(_08922_));
 AO21x1_ASAP7_75t_R _27189_ (.A1(_08610_),
    .A2(_08922_),
    .B(_01727_),
    .Y(_08923_));
 OA21x2_ASAP7_75t_R _27190_ (.A1(_00285_),
    .A2(_06426_),
    .B(_08695_),
    .Y(_08924_));
 OA21x2_ASAP7_75t_R _27191_ (.A1(_01357_),
    .A2(_08912_),
    .B(_08924_),
    .Y(_08925_));
 OAI21x1_ASAP7_75t_R _27192_ (.A1(_08920_),
    .A2(_08923_),
    .B(_08925_),
    .Y(_08926_));
 OA211x2_ASAP7_75t_R _27193_ (.A1(_16132_),
    .A2(_08600_),
    .B(_08163_),
    .C(_13576_),
    .Y(_08927_));
 AND3x1_ASAP7_75t_R _27194_ (.A(_08591_),
    .B(_08926_),
    .C(_08927_),
    .Y(_08928_));
 AO21x1_ASAP7_75t_R _27195_ (.A1(_16087_),
    .A2(_08590_),
    .B(_08928_),
    .Y(_02707_));
 NAND2x1_ASAP7_75t_R _27196_ (.A(_08203_),
    .B(_08591_),
    .Y(_08929_));
 OA21x2_ASAP7_75t_R _27197_ (.A1(_00946_),
    .A2(_08591_),
    .B(_08929_),
    .Y(_08930_));
 AND2x2_ASAP7_75t_R _27198_ (.A(_16260_),
    .B(_08614_),
    .Y(_08931_));
 AO21x1_ASAP7_75t_R _27199_ (.A1(_00946_),
    .A2(_08607_),
    .B(_08931_),
    .Y(_08932_));
 NAND2x2_ASAP7_75t_R _27200_ (.A(_05751_),
    .B(_01322_),
    .Y(_08933_));
 OR3x1_ASAP7_75t_R _27201_ (.A(_01321_),
    .B(_08748_),
    .C(_08933_),
    .Y(_08934_));
 AO21x1_ASAP7_75t_R _27202_ (.A1(_01344_),
    .A2(_08934_),
    .B(_08610_),
    .Y(_08935_));
 OA21x2_ASAP7_75t_R _27203_ (.A1(_08738_),
    .A2(_08932_),
    .B(_08935_),
    .Y(_08936_));
 OA21x2_ASAP7_75t_R _27204_ (.A1(_00285_),
    .A2(_16260_),
    .B(_08576_),
    .Y(_08937_));
 OA21x2_ASAP7_75t_R _27205_ (.A1(_01357_),
    .A2(_08922_),
    .B(_08937_),
    .Y(_08938_));
 AO21x1_ASAP7_75t_R _27206_ (.A1(_06799_),
    .A2(_08801_),
    .B(_08938_),
    .Y(_08939_));
 OA211x2_ASAP7_75t_R _27207_ (.A1(_01727_),
    .A2(_08936_),
    .B(_08939_),
    .C(_08786_),
    .Y(_08940_));
 NOR2x1_ASAP7_75t_R _27208_ (.A(_08930_),
    .B(_08940_),
    .Y(_02708_));
 OA21x2_ASAP7_75t_R _27209_ (.A1(_00285_),
    .A2(_06440_),
    .B(_08576_),
    .Y(_08941_));
 OAI21x1_ASAP7_75t_R _27210_ (.A1(_01357_),
    .A2(_08932_),
    .B(_08941_),
    .Y(_08942_));
 OA21x2_ASAP7_75t_R _27211_ (.A1(_16372_),
    .A2(_08788_),
    .B(_08942_),
    .Y(_08943_));
 OR5x1_ASAP7_75t_R _27212_ (.A(_01319_),
    .B(_01318_),
    .C(_08746_),
    .D(_17607_),
    .E(_08607_),
    .Y(_08944_));
 AND3x1_ASAP7_75t_R _27213_ (.A(_01345_),
    .B(_08598_),
    .C(_08944_),
    .Y(_08945_));
 INVx1_ASAP7_75t_R _27214_ (.A(_08945_),
    .Y(_08946_));
 AND2x2_ASAP7_75t_R _27215_ (.A(_06737_),
    .B(_08607_),
    .Y(_08947_));
 AO21x1_ASAP7_75t_R _27216_ (.A1(net162),
    .A2(_08614_),
    .B(_08947_),
    .Y(_08948_));
 INVx1_ASAP7_75t_R _27217_ (.A(_01727_),
    .Y(_08949_));
 OA21x2_ASAP7_75t_R _27218_ (.A1(_08738_),
    .A2(_08948_),
    .B(_08949_),
    .Y(_08950_));
 AO21x1_ASAP7_75t_R _27219_ (.A1(_08946_),
    .A2(_08950_),
    .B(_07076_),
    .Y(_08951_));
 OA211x2_ASAP7_75t_R _27220_ (.A1(_08943_),
    .A2(_08951_),
    .B(_08230_),
    .C(_08591_),
    .Y(_08952_));
 AO21x1_ASAP7_75t_R _27221_ (.A1(_06737_),
    .A2(_08590_),
    .B(_08952_),
    .Y(_02709_));
 OR3x4_ASAP7_75t_R _27222_ (.A(_17607_),
    .B(_08607_),
    .C(_08933_),
    .Y(_08953_));
 OA211x2_ASAP7_75t_R _27223_ (.A1(_01326_),
    .A2(_08953_),
    .B(_08861_),
    .C(_01346_),
    .Y(_08954_));
 AND2x2_ASAP7_75t_R _27224_ (.A(_05760_),
    .B(_08614_),
    .Y(_08955_));
 AO21x1_ASAP7_75t_R _27225_ (.A1(_01011_),
    .A2(_08607_),
    .B(_08955_),
    .Y(_08956_));
 AO21x1_ASAP7_75t_R _27226_ (.A1(_08610_),
    .A2(_08956_),
    .B(_01727_),
    .Y(_08957_));
 OAI21x1_ASAP7_75t_R _27227_ (.A1(_08954_),
    .A2(_08957_),
    .B(_05745_),
    .Y(_08958_));
 AO221x1_ASAP7_75t_R _27228_ (.A1(_13530_),
    .A2(net163),
    .B1(_08948_),
    .B2(_05741_),
    .C(_08791_),
    .Y(_08959_));
 OA21x2_ASAP7_75t_R _27229_ (.A1(_05849_),
    .A2(_08788_),
    .B(_08959_),
    .Y(_08960_));
 OA211x2_ASAP7_75t_R _27230_ (.A1(_05745_),
    .A2(_08280_),
    .B(_08591_),
    .C(_13576_),
    .Y(_08961_));
 OA21x2_ASAP7_75t_R _27231_ (.A1(_08958_),
    .A2(_08960_),
    .B(_08961_),
    .Y(_08962_));
 AO21x1_ASAP7_75t_R _27232_ (.A1(_06806_),
    .A2(_08590_),
    .B(_08962_),
    .Y(_02710_));
 INVx1_ASAP7_75t_R _27233_ (.A(_01045_),
    .Y(_08963_));
 OA21x2_ASAP7_75t_R _27234_ (.A1(_00285_),
    .A2(_06452_),
    .B(_08695_),
    .Y(_08964_));
 OAI21x1_ASAP7_75t_R _27235_ (.A1(_01357_),
    .A2(_08956_),
    .B(_08964_),
    .Y(_08965_));
 AND2x2_ASAP7_75t_R _27236_ (.A(_06452_),
    .B(_08614_),
    .Y(_08966_));
 AO21x1_ASAP7_75t_R _27237_ (.A1(_01045_),
    .A2(_08607_),
    .B(_08966_),
    .Y(_08967_));
 OA211x2_ASAP7_75t_R _27238_ (.A1(_01320_),
    .A2(_08953_),
    .B(_08861_),
    .C(_01347_),
    .Y(_08968_));
 AOI211x1_ASAP7_75t_R _27239_ (.A1(_08610_),
    .A2(_08967_),
    .B(_08968_),
    .C(_01727_),
    .Y(_08969_));
 OA21x2_ASAP7_75t_R _27240_ (.A1(_04595_),
    .A2(_08600_),
    .B(_08302_),
    .Y(_08970_));
 OA211x2_ASAP7_75t_R _27241_ (.A1(_08965_),
    .A2(_08969_),
    .B(_08970_),
    .C(_08591_),
    .Y(_08971_));
 AO21x1_ASAP7_75t_R _27242_ (.A1(_08963_),
    .A2(_08590_),
    .B(_08971_),
    .Y(_02711_));
 OR3x1_ASAP7_75t_R _27243_ (.A(_04715_),
    .B(_08590_),
    .C(_08600_),
    .Y(_08972_));
 INVx1_ASAP7_75t_R _27244_ (.A(_08972_),
    .Y(_08973_));
 AO221x1_ASAP7_75t_R _27245_ (.A1(_14626_),
    .A2(_08350_),
    .B1(_08590_),
    .B2(_01077_),
    .C(_08973_),
    .Y(_08974_));
 OR3x4_ASAP7_75t_R _27246_ (.A(_01318_),
    .B(_01322_),
    .C(_08819_),
    .Y(_08975_));
 OA211x2_ASAP7_75t_R _27247_ (.A1(_01321_),
    .A2(_08975_),
    .B(_08598_),
    .C(_01348_),
    .Y(_08976_));
 AND2x2_ASAP7_75t_R _27248_ (.A(_04719_),
    .B(_08614_),
    .Y(_08977_));
 AO21x1_ASAP7_75t_R _27249_ (.A1(_01077_),
    .A2(_08607_),
    .B(_08977_),
    .Y(_08978_));
 AO21x1_ASAP7_75t_R _27250_ (.A1(_08610_),
    .A2(_08978_),
    .B(_01727_),
    .Y(_08979_));
 OA211x2_ASAP7_75t_R _27251_ (.A1(_00285_),
    .A2(_04719_),
    .B(_08576_),
    .C(_08786_),
    .Y(_08980_));
 OA21x2_ASAP7_75t_R _27252_ (.A1(_01357_),
    .A2(_08967_),
    .B(_08980_),
    .Y(_08981_));
 OA21x2_ASAP7_75t_R _27253_ (.A1(_08976_),
    .A2(_08979_),
    .B(_08981_),
    .Y(_08982_));
 NOR2x1_ASAP7_75t_R _27254_ (.A(_08974_),
    .B(_08982_),
    .Y(_02712_));
 NAND2x1_ASAP7_75t_R _27255_ (.A(_06750_),
    .B(_08607_),
    .Y(_08983_));
 OA21x2_ASAP7_75t_R _27256_ (.A1(_06464_),
    .A2(_08607_),
    .B(_08983_),
    .Y(_08984_));
 OR3x2_ASAP7_75t_R _27257_ (.A(_01319_),
    .B(_01318_),
    .C(_01322_),
    .Y(_08985_));
 OA211x2_ASAP7_75t_R _27258_ (.A1(_08819_),
    .A2(_08985_),
    .B(_01349_),
    .C(_08738_),
    .Y(_08986_));
 AO21x1_ASAP7_75t_R _27259_ (.A1(_08610_),
    .A2(_08984_),
    .B(_08986_),
    .Y(_08987_));
 OA21x2_ASAP7_75t_R _27260_ (.A1(_00285_),
    .A2(_06464_),
    .B(_08695_),
    .Y(_08988_));
 OA21x2_ASAP7_75t_R _27261_ (.A1(_01357_),
    .A2(_08978_),
    .B(_08988_),
    .Y(_08989_));
 OAI21x1_ASAP7_75t_R _27262_ (.A1(_01727_),
    .A2(_08987_),
    .B(_08989_),
    .Y(_08990_));
 OA21x2_ASAP7_75t_R _27263_ (.A1(_04828_),
    .A2(_08600_),
    .B(_08371_),
    .Y(_08991_));
 AO21x1_ASAP7_75t_R _27264_ (.A1(_08990_),
    .A2(_08991_),
    .B(_08590_),
    .Y(_08992_));
 OA21x2_ASAP7_75t_R _27265_ (.A1(_06750_),
    .A2(_08591_),
    .B(_08992_),
    .Y(_02713_));
 OA211x2_ASAP7_75t_R _27266_ (.A1(_01326_),
    .A2(_08975_),
    .B(_08738_),
    .C(_01350_),
    .Y(_08993_));
 AND2x2_ASAP7_75t_R _27267_ (.A(_04937_),
    .B(_08614_),
    .Y(_08994_));
 AO21x1_ASAP7_75t_R _27268_ (.A1(_01142_),
    .A2(_08607_),
    .B(_08994_),
    .Y(_08995_));
 AO21x1_ASAP7_75t_R _27269_ (.A1(_08610_),
    .A2(_08995_),
    .B(_01727_),
    .Y(_08996_));
 OA21x2_ASAP7_75t_R _27270_ (.A1(_00285_),
    .A2(_04937_),
    .B(_08695_),
    .Y(_08997_));
 OA21x2_ASAP7_75t_R _27271_ (.A1(_01357_),
    .A2(_08984_),
    .B(_08997_),
    .Y(_08998_));
 OAI21x1_ASAP7_75t_R _27272_ (.A1(_08993_),
    .A2(_08996_),
    .B(_08998_),
    .Y(_08999_));
 AO21x1_ASAP7_75t_R _27273_ (.A1(_04910_),
    .A2(_04934_),
    .B(_08600_),
    .Y(_09000_));
 AND5x1_ASAP7_75t_R _27274_ (.A(_13576_),
    .B(_08398_),
    .C(_08591_),
    .D(_08999_),
    .E(_09000_),
    .Y(_09001_));
 AO21x1_ASAP7_75t_R _27275_ (.A1(_06813_),
    .A2(_08590_),
    .B(_09001_),
    .Y(_02714_));
 OA211x2_ASAP7_75t_R _27276_ (.A1(_01320_),
    .A2(_08975_),
    .B(_08598_),
    .C(_01351_),
    .Y(_09002_));
 AND2x2_ASAP7_75t_R _27277_ (.A(_06477_),
    .B(_08614_),
    .Y(_09003_));
 AO21x1_ASAP7_75t_R _27278_ (.A1(_01176_),
    .A2(_08607_),
    .B(_09003_),
    .Y(_09004_));
 AO21x1_ASAP7_75t_R _27279_ (.A1(_08610_),
    .A2(_09004_),
    .B(_01727_),
    .Y(_09005_));
 OA21x2_ASAP7_75t_R _27280_ (.A1(_00285_),
    .A2(_06477_),
    .B(_08695_),
    .Y(_09006_));
 OA21x2_ASAP7_75t_R _27281_ (.A1(_01357_),
    .A2(_08995_),
    .B(_09006_),
    .Y(_09007_));
 OAI21x1_ASAP7_75t_R _27282_ (.A1(_09002_),
    .A2(_09005_),
    .B(_09007_),
    .Y(_09008_));
 OA211x2_ASAP7_75t_R _27283_ (.A1(_05044_),
    .A2(_08600_),
    .B(_08430_),
    .C(_13576_),
    .Y(_09009_));
 AND3x1_ASAP7_75t_R _27284_ (.A(_08591_),
    .B(_09008_),
    .C(_09009_),
    .Y(_09010_));
 AO21x1_ASAP7_75t_R _27285_ (.A1(_06815_),
    .A2(_08590_),
    .B(_09010_),
    .Y(_02715_));
 AND2x2_ASAP7_75t_R _27286_ (.A(_05154_),
    .B(_08614_),
    .Y(_09011_));
 AO21x1_ASAP7_75t_R _27287_ (.A1(_01208_),
    .A2(_08607_),
    .B(_09011_),
    .Y(_09012_));
 OR3x4_ASAP7_75t_R _27288_ (.A(_01318_),
    .B(_01322_),
    .C(_08748_),
    .Y(_09013_));
 OA211x2_ASAP7_75t_R _27289_ (.A1(_01321_),
    .A2(_09013_),
    .B(_08738_),
    .C(_01352_),
    .Y(_09014_));
 AO21x1_ASAP7_75t_R _27290_ (.A1(_08610_),
    .A2(_09012_),
    .B(_09014_),
    .Y(_09015_));
 OA21x2_ASAP7_75t_R _27291_ (.A1(_00285_),
    .A2(_05154_),
    .B(_08576_),
    .Y(_09016_));
 OAI21x1_ASAP7_75t_R _27292_ (.A1(_01357_),
    .A2(_09004_),
    .B(_09016_),
    .Y(_09017_));
 OAI21x1_ASAP7_75t_R _27293_ (.A1(_05891_),
    .A2(_08788_),
    .B(_09017_),
    .Y(_09018_));
 OA211x2_ASAP7_75t_R _27294_ (.A1(_01727_),
    .A2(_09015_),
    .B(_09018_),
    .C(_08786_),
    .Y(_09019_));
 AOI221x1_ASAP7_75t_R _27295_ (.A1(_14626_),
    .A2(_08457_),
    .B1(_08590_),
    .B2(_01208_),
    .C(_09019_),
    .Y(_02716_));
 OR3x1_ASAP7_75t_R _27296_ (.A(_17607_),
    .B(_08607_),
    .C(_08985_),
    .Y(_09020_));
 AND2x2_ASAP7_75t_R _27297_ (.A(_06491_),
    .B(_08614_),
    .Y(_09021_));
 AO21x1_ASAP7_75t_R _27298_ (.A1(_01242_),
    .A2(_08607_),
    .B(_09021_),
    .Y(_09022_));
 AO32x1_ASAP7_75t_R _27299_ (.A1(_01353_),
    .A2(_08598_),
    .A3(_09020_),
    .B1(_09022_),
    .B2(_08610_),
    .Y(_09023_));
 OA21x2_ASAP7_75t_R _27300_ (.A1(_00285_),
    .A2(_06491_),
    .B(_08576_),
    .Y(_09024_));
 OA21x2_ASAP7_75t_R _27301_ (.A1(_01357_),
    .A2(_09012_),
    .B(_09024_),
    .Y(_09025_));
 AO21x1_ASAP7_75t_R _27302_ (.A1(_05261_),
    .A2(_08801_),
    .B(_09025_),
    .Y(_09026_));
 OA211x2_ASAP7_75t_R _27303_ (.A1(_01727_),
    .A2(_09023_),
    .B(_09026_),
    .C(_08786_),
    .Y(_09027_));
 AND2x2_ASAP7_75t_R _27304_ (.A(_08495_),
    .B(_08591_),
    .Y(_09028_));
 AOI211x1_ASAP7_75t_R _27305_ (.A1(_01242_),
    .A2(_08590_),
    .B(_09027_),
    .C(_09028_),
    .Y(_02717_));
 OA211x2_ASAP7_75t_R _27306_ (.A1(_01326_),
    .A2(_09013_),
    .B(_08861_),
    .C(_01354_),
    .Y(_09029_));
 AND2x2_ASAP7_75t_R _27307_ (.A(_05372_),
    .B(_08614_),
    .Y(_09030_));
 AO21x1_ASAP7_75t_R _27308_ (.A1(_01274_),
    .A2(_08607_),
    .B(_09030_),
    .Y(_09031_));
 AO21x1_ASAP7_75t_R _27309_ (.A1(_08610_),
    .A2(_09031_),
    .B(_01727_),
    .Y(_09032_));
 OAI22x1_ASAP7_75t_R _27310_ (.A1(_00285_),
    .A2(_05372_),
    .B1(_09022_),
    .B2(_01357_),
    .Y(_09033_));
 OAI22x1_ASAP7_75t_R _27311_ (.A1(_05369_),
    .A2(_08788_),
    .B1(_09033_),
    .B2(_08791_),
    .Y(_09034_));
 OA211x2_ASAP7_75t_R _27312_ (.A1(_09029_),
    .A2(_09032_),
    .B(_09034_),
    .C(_08786_),
    .Y(_09035_));
 AOI221x1_ASAP7_75t_R _27313_ (.A1(_14626_),
    .A2(_08519_),
    .B1(_08590_),
    .B2(_01274_),
    .C(_09035_),
    .Y(_02718_));
 OA211x2_ASAP7_75t_R _27314_ (.A1(_01320_),
    .A2(_09013_),
    .B(_08598_),
    .C(_01355_),
    .Y(_09036_));
 AO21x1_ASAP7_75t_R _27315_ (.A1(_05503_),
    .A2(net173),
    .B(_08738_),
    .Y(_09037_));
 NAND2x1_ASAP7_75t_R _27316_ (.A(_08949_),
    .B(_09037_),
    .Y(_09038_));
 OA21x2_ASAP7_75t_R _27317_ (.A1(_00285_),
    .A2(_05512_),
    .B(_08576_),
    .Y(_09039_));
 OA21x2_ASAP7_75t_R _27318_ (.A1(_01357_),
    .A2(_09031_),
    .B(_09039_),
    .Y(_09040_));
 OAI21x1_ASAP7_75t_R _27319_ (.A1(_09036_),
    .A2(_09038_),
    .B(_09040_),
    .Y(_09041_));
 TAPCELL_ASAP7_75t_R TAP_667 ();
 OA21x2_ASAP7_75t_R _27321_ (.A1(_05474_),
    .A2(_08788_),
    .B(_08786_),
    .Y(_09043_));
 AND2x2_ASAP7_75t_R _27322_ (.A(_08549_),
    .B(_08591_),
    .Y(_09044_));
 AO221x1_ASAP7_75t_R _27323_ (.A1(_05503_),
    .A2(_08590_),
    .B1(_09041_),
    .B2(_09043_),
    .C(_09044_),
    .Y(_02719_));
 INVx1_ASAP7_75t_R _27324_ (.A(_01677_),
    .Y(_09045_));
 AO32x1_ASAP7_75t_R _27325_ (.A1(_05503_),
    .A2(_05741_),
    .A3(net173),
    .B1(_08791_),
    .B2(_08598_),
    .Y(_09046_));
 AO221x1_ASAP7_75t_R _27326_ (.A1(_02261_),
    .A2(_07078_),
    .B1(_09046_),
    .B2(_05745_),
    .C(_08590_),
    .Y(_09047_));
 OA21x2_ASAP7_75t_R _27327_ (.A1(_09045_),
    .A2(_08591_),
    .B(_09047_),
    .Y(_02720_));
 INVx1_ASAP7_75t_R _27328_ (.A(_00034_),
    .Y(_09048_));
 XNOR2x1_ASAP7_75t_R _27329_ (.B(_02256_),
    .Y(_09049_),
    .A(_00070_));
 XNOR2x1_ASAP7_75t_R _27330_ (.B(_17526_),
    .Y(_09050_),
    .A(_00069_));
 XNOR2x1_ASAP7_75t_R _27331_ (.B(_09050_),
    .Y(_09051_),
    .A(_09049_));
 XNOR2x1_ASAP7_75t_R _27332_ (.B(_17502_),
    .Y(_09052_),
    .A(_00068_));
 XNOR2x1_ASAP7_75t_R _27333_ (.B(_09052_),
    .Y(_09053_),
    .A(_09051_));
 XOR2x2_ASAP7_75t_R _27334_ (.A(_00051_),
    .B(_02352_),
    .Y(_09054_));
 XNOR2x1_ASAP7_75t_R _27335_ (.B(_00071_),
    .Y(_09055_),
    .A(_17471_));
 XNOR2x1_ASAP7_75t_R _27336_ (.B(_09055_),
    .Y(_09056_),
    .A(_09054_));
 XNOR2x1_ASAP7_75t_R _27337_ (.B(_02260_),
    .Y(_09057_),
    .A(_02259_));
 XNOR2x1_ASAP7_75t_R _27338_ (.B(_02258_),
    .Y(_09058_),
    .A(_02257_));
 XNOR2x1_ASAP7_75t_R _27339_ (.B(_09058_),
    .Y(_09059_),
    .A(_09057_));
 XNOR2x1_ASAP7_75t_R _27340_ (.B(_09059_),
    .Y(_09060_),
    .A(_09056_));
 XNOR2x1_ASAP7_75t_R _27341_ (.B(_09060_),
    .Y(_09061_),
    .A(_09053_));
 OA21x2_ASAP7_75t_R _27342_ (.A1(_00034_),
    .A2(_05519_),
    .B(_05931_),
    .Y(_09062_));
 XNOR2x1_ASAP7_75t_R _27343_ (.B(_09062_),
    .Y(_09063_),
    .A(_09061_));
 NAND2x1_ASAP7_75t_R _27344_ (.A(_17494_),
    .B(_17518_),
    .Y(_09064_));
 XNOR2x1_ASAP7_75t_R _27345_ (.B(_09064_),
    .Y(_09065_),
    .A(_09063_));
 AO221x1_ASAP7_75t_R _27346_ (.A1(_08791_),
    .A2(_08598_),
    .B1(_09065_),
    .B2(_07078_),
    .C(_08590_),
    .Y(_09066_));
 OA21x2_ASAP7_75t_R _27347_ (.A1(_09048_),
    .A2(_08591_),
    .B(_09066_),
    .Y(_02721_));
 NAND2x2_ASAP7_75t_R _27348_ (.A(_06705_),
    .B(_05757_),
    .Y(_09067_));
 TAPCELL_ASAP7_75t_R TAP_666 ();
 TAPCELL_ASAP7_75t_R TAP_665 ();
 TAPCELL_ASAP7_75t_R TAP_664 ();
 AND2x6_ASAP7_75t_R _27352_ (.A(_06705_),
    .B(_05757_),
    .Y(_09071_));
 TAPCELL_ASAP7_75t_R TAP_663 ();
 TAPCELL_ASAP7_75t_R TAP_662 ();
 NAND2x1_ASAP7_75t_R _27355_ (.A(_13758_),
    .B(_08582_),
    .Y(_09074_));
 OA211x2_ASAP7_75t_R _27356_ (.A1(_16503_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09074_),
    .Y(_09075_));
 AOI21x1_ASAP7_75t_R _27357_ (.A1(_01676_),
    .A2(_09067_),
    .B(_09075_),
    .Y(_02722_));
 AND3x1_ASAP7_75t_R _27358_ (.A(\ex_block_i.alu_adder_result_ex_o[1] ),
    .B(_05474_),
    .C(_05915_),
    .Y(_09076_));
 AO21x1_ASAP7_75t_R _27359_ (.A1(_13523_),
    .A2(_08582_),
    .B(_09076_),
    .Y(_09077_));
 OR2x2_ASAP7_75t_R _27360_ (.A(_09067_),
    .B(_09077_),
    .Y(_09078_));
 OA21x2_ASAP7_75t_R _27361_ (.A1(_08625_),
    .A2(_09071_),
    .B(_09078_),
    .Y(_02723_));
 NAND2x1_ASAP7_75t_R _27362_ (.A(_14684_),
    .B(_08582_),
    .Y(_09079_));
 OA211x2_ASAP7_75t_R _27363_ (.A1(_05767_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09079_),
    .Y(_09080_));
 AOI21x1_ASAP7_75t_R _27364_ (.A1(_01674_),
    .A2(_09067_),
    .B(_09080_),
    .Y(_02724_));
 INVx1_ASAP7_75t_R _27365_ (.A(_01673_),
    .Y(_09081_));
 TAPCELL_ASAP7_75t_R TAP_661 ();
 TAPCELL_ASAP7_75t_R TAP_660 ();
 TAPCELL_ASAP7_75t_R TAP_659 ();
 TAPCELL_ASAP7_75t_R TAP_658 ();
 AO21x1_ASAP7_75t_R _27370_ (.A1(_05474_),
    .A2(_05915_),
    .B(_14752_),
    .Y(_09086_));
 OA211x2_ASAP7_75t_R _27371_ (.A1(net174),
    .A2(_08582_),
    .B(_09071_),
    .C(_09086_),
    .Y(_09087_));
 AO21x1_ASAP7_75t_R _27372_ (.A1(_09081_),
    .A2(_09067_),
    .B(_09087_),
    .Y(_02725_));
 NAND2x1_ASAP7_75t_R _27373_ (.A(_14820_),
    .B(_08582_),
    .Y(_09088_));
 OA211x2_ASAP7_75t_R _27374_ (.A1(_05766_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09088_),
    .Y(_09089_));
 AOI21x1_ASAP7_75t_R _27375_ (.A1(_01672_),
    .A2(_09067_),
    .B(_09089_),
    .Y(_02726_));
 AO21x1_ASAP7_75t_R _27376_ (.A1(_05474_),
    .A2(_05915_),
    .B(_14873_),
    .Y(_09090_));
 OA211x2_ASAP7_75t_R _27377_ (.A1(net176),
    .A2(_08582_),
    .B(_09071_),
    .C(_09090_),
    .Y(_09091_));
 AO21x1_ASAP7_75t_R _27378_ (.A1(_08643_),
    .A2(_09067_),
    .B(_09091_),
    .Y(_02727_));
 NAND2x1_ASAP7_75t_R _27379_ (.A(_14936_),
    .B(_08582_),
    .Y(_09092_));
 OA211x2_ASAP7_75t_R _27380_ (.A1(_05768_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09092_),
    .Y(_09093_));
 AOI21x1_ASAP7_75t_R _27381_ (.A1(_01670_),
    .A2(_09067_),
    .B(_09093_),
    .Y(_02728_));
 OR2x2_ASAP7_75t_R _27382_ (.A(_06710_),
    .B(_08577_),
    .Y(_09094_));
 OA211x2_ASAP7_75t_R _27383_ (.A1(_00676_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09094_),
    .Y(_09095_));
 AOI21x1_ASAP7_75t_R _27384_ (.A1(_01669_),
    .A2(_09067_),
    .B(_09095_),
    .Y(_02729_));
 INVx1_ASAP7_75t_R _27385_ (.A(_01668_),
    .Y(_09096_));
 AO21x1_ASAP7_75t_R _27386_ (.A1(_05474_),
    .A2(_05915_),
    .B(_15042_),
    .Y(_09097_));
 OA211x2_ASAP7_75t_R _27387_ (.A1(net179),
    .A2(_08582_),
    .B(_09071_),
    .C(_09097_),
    .Y(_09098_));
 AO21x1_ASAP7_75t_R _27388_ (.A1(_09096_),
    .A2(_09067_),
    .B(_09098_),
    .Y(_02730_));
 AO21x1_ASAP7_75t_R _27389_ (.A1(_05474_),
    .A2(_05915_),
    .B(_15096_),
    .Y(_09099_));
 OA211x2_ASAP7_75t_R _27390_ (.A1(net180),
    .A2(_08582_),
    .B(_09071_),
    .C(_09099_),
    .Y(_09100_));
 AO21x1_ASAP7_75t_R _27391_ (.A1(_08633_),
    .A2(_09067_),
    .B(_09100_),
    .Y(_02731_));
 NAND2x1_ASAP7_75t_R _27392_ (.A(_15157_),
    .B(_08582_),
    .Y(_09101_));
 OA211x2_ASAP7_75t_R _27393_ (.A1(_05772_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09101_),
    .Y(_09102_));
 AOI21x1_ASAP7_75t_R _27394_ (.A1(_01666_),
    .A2(_09067_),
    .B(_09102_),
    .Y(_02732_));
 INVx1_ASAP7_75t_R _27395_ (.A(_01665_),
    .Y(_09103_));
 TAPCELL_ASAP7_75t_R TAP_657 ();
 AO21x1_ASAP7_75t_R _27397_ (.A1(_05474_),
    .A2(_05915_),
    .B(_14574_),
    .Y(_09105_));
 OA211x2_ASAP7_75t_R _27398_ (.A1(net152),
    .A2(_08582_),
    .B(_09071_),
    .C(_09105_),
    .Y(_09106_));
 AO21x1_ASAP7_75t_R _27399_ (.A1(_09103_),
    .A2(_09067_),
    .B(_09106_),
    .Y(_02733_));
 OR2x2_ASAP7_75t_R _27400_ (.A(_13878_),
    .B(_08577_),
    .Y(_09107_));
 OA211x2_ASAP7_75t_R _27401_ (.A1(_05771_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09107_),
    .Y(_09108_));
 AOI21x1_ASAP7_75t_R _27402_ (.A1(_01664_),
    .A2(_09067_),
    .B(_09108_),
    .Y(_02734_));
 TAPCELL_ASAP7_75t_R TAP_656 ();
 AO21x1_ASAP7_75t_R _27404_ (.A1(_05474_),
    .A2(_05915_),
    .B(_15401_),
    .Y(_09110_));
 OA211x2_ASAP7_75t_R _27405_ (.A1(net154),
    .A2(_08582_),
    .B(_09071_),
    .C(_09110_),
    .Y(_09111_));
 AO21x1_ASAP7_75t_R _27406_ (.A1(_08650_),
    .A2(_09067_),
    .B(_09111_),
    .Y(_02735_));
 AO21x1_ASAP7_75t_R _27407_ (.A1(_05474_),
    .A2(_05915_),
    .B(_15555_),
    .Y(_09112_));
 OA211x2_ASAP7_75t_R _27408_ (.A1(_15557_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09112_),
    .Y(_09113_));
 AOI21x1_ASAP7_75t_R _27409_ (.A1(_01662_),
    .A2(_09067_),
    .B(_09113_),
    .Y(_02736_));
 INVx1_ASAP7_75t_R _27410_ (.A(_01661_),
    .Y(_09114_));
 AO21x1_ASAP7_75t_R _27411_ (.A1(_05474_),
    .A2(_05915_),
    .B(_15665_),
    .Y(_09115_));
 OA211x2_ASAP7_75t_R _27412_ (.A1(net156),
    .A2(_08582_),
    .B(_09071_),
    .C(_09115_),
    .Y(_09116_));
 AO21x1_ASAP7_75t_R _27413_ (.A1(_09114_),
    .A2(_09067_),
    .B(_09116_),
    .Y(_02737_));
 NAND2x1_ASAP7_75t_R _27414_ (.A(_05770_),
    .B(_08577_),
    .Y(_09117_));
 OA211x2_ASAP7_75t_R _27415_ (.A1(_06792_),
    .A2(_08577_),
    .B(_09071_),
    .C(_09117_),
    .Y(_09118_));
 AO21x1_ASAP7_75t_R _27416_ (.A1(_08662_),
    .A2(_09067_),
    .B(_09118_),
    .Y(_02738_));
 AO21x1_ASAP7_75t_R _27417_ (.A1(_05474_),
    .A2(_05915_),
    .B(_15890_),
    .Y(_09119_));
 OA211x2_ASAP7_75t_R _27418_ (.A1(net158),
    .A2(_08582_),
    .B(_09071_),
    .C(_09119_),
    .Y(_09120_));
 AO21x1_ASAP7_75t_R _27419_ (.A1(_08665_),
    .A2(_09067_),
    .B(_09120_),
    .Y(_02739_));
 OR2x2_ASAP7_75t_R _27420_ (.A(_16018_),
    .B(_08577_),
    .Y(_09121_));
 OA211x2_ASAP7_75t_R _27421_ (.A1(_16020_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09121_),
    .Y(_09122_));
 AOI21x1_ASAP7_75t_R _27422_ (.A1(_01658_),
    .A2(_09067_),
    .B(_09122_),
    .Y(_02740_));
 INVx1_ASAP7_75t_R _27423_ (.A(_01657_),
    .Y(_09123_));
 AO21x1_ASAP7_75t_R _27424_ (.A1(_05474_),
    .A2(_05915_),
    .B(_16132_),
    .Y(_09124_));
 OA211x2_ASAP7_75t_R _27425_ (.A1(net257),
    .A2(_08582_),
    .B(_09071_),
    .C(_09124_),
    .Y(_09125_));
 AO21x1_ASAP7_75t_R _27426_ (.A1(_09123_),
    .A2(_09067_),
    .B(_09125_),
    .Y(_02741_));
 NAND2x1_ASAP7_75t_R _27427_ (.A(_16256_),
    .B(_08582_),
    .Y(_09126_));
 OA211x2_ASAP7_75t_R _27428_ (.A1(_16260_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09126_),
    .Y(_09127_));
 AOI21x1_ASAP7_75t_R _27429_ (.A1(_01656_),
    .A2(_09067_),
    .B(_09127_),
    .Y(_02742_));
 AO21x1_ASAP7_75t_R _27430_ (.A1(_05474_),
    .A2(_05915_),
    .B(_16372_),
    .Y(_09128_));
 OA211x2_ASAP7_75t_R _27431_ (.A1(net162),
    .A2(_08582_),
    .B(_09071_),
    .C(_09128_),
    .Y(_09129_));
 AO21x1_ASAP7_75t_R _27432_ (.A1(_08687_),
    .A2(_09067_),
    .B(_09129_),
    .Y(_02743_));
 AO21x1_ASAP7_75t_R _27433_ (.A1(_05474_),
    .A2(_05915_),
    .B(_05849_),
    .Y(_09130_));
 OA211x2_ASAP7_75t_R _27434_ (.A1(net163),
    .A2(_08582_),
    .B(_09071_),
    .C(_09130_),
    .Y(_09131_));
 AO21x1_ASAP7_75t_R _27435_ (.A1(_08684_),
    .A2(_09067_),
    .B(_09131_),
    .Y(_02744_));
 NAND2x1_ASAP7_75t_R _27436_ (.A(_04595_),
    .B(_08582_),
    .Y(_09132_));
 OA211x2_ASAP7_75t_R _27437_ (.A1(_06452_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09132_),
    .Y(_09133_));
 AOI21x1_ASAP7_75t_R _27438_ (.A1(_01653_),
    .A2(_09067_),
    .B(_09133_),
    .Y(_02745_));
 NAND2x1_ASAP7_75t_R _27439_ (.A(_04715_),
    .B(_08582_),
    .Y(_09134_));
 OA211x2_ASAP7_75t_R _27440_ (.A1(_04719_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09134_),
    .Y(_09135_));
 AOI21x1_ASAP7_75t_R _27441_ (.A1(_01652_),
    .A2(_09067_),
    .B(_09135_),
    .Y(_02746_));
 AO21x1_ASAP7_75t_R _27442_ (.A1(_05474_),
    .A2(_05915_),
    .B(_04828_),
    .Y(_09136_));
 OA211x2_ASAP7_75t_R _27443_ (.A1(net166),
    .A2(_08582_),
    .B(_09071_),
    .C(_09136_),
    .Y(_09137_));
 AO21x1_ASAP7_75t_R _27444_ (.A1(_08672_),
    .A2(_09067_),
    .B(_09137_),
    .Y(_02747_));
 OR2x2_ASAP7_75t_R _27445_ (.A(_04935_),
    .B(_08577_),
    .Y(_09138_));
 OA211x2_ASAP7_75t_R _27446_ (.A1(_04937_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09138_),
    .Y(_09139_));
 AOI21x1_ASAP7_75t_R _27447_ (.A1(_01650_),
    .A2(_09067_),
    .B(_09139_),
    .Y(_02748_));
 NAND2x1_ASAP7_75t_R _27448_ (.A(_05044_),
    .B(_08582_),
    .Y(_09140_));
 OA211x2_ASAP7_75t_R _27449_ (.A1(_06477_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09140_),
    .Y(_09141_));
 AOI21x1_ASAP7_75t_R _27450_ (.A1(_01649_),
    .A2(_09067_),
    .B(_09141_),
    .Y(_02749_));
 AO21x1_ASAP7_75t_R _27451_ (.A1(_05474_),
    .A2(_05915_),
    .B(_05891_),
    .Y(_09142_));
 OA211x2_ASAP7_75t_R _27452_ (.A1(net169),
    .A2(_08582_),
    .B(_09071_),
    .C(_09142_),
    .Y(_09143_));
 AO21x1_ASAP7_75t_R _27453_ (.A1(_08680_),
    .A2(_09067_),
    .B(_09143_),
    .Y(_02750_));
 OR2x2_ASAP7_75t_R _27454_ (.A(_05261_),
    .B(_08577_),
    .Y(_09144_));
 OA211x2_ASAP7_75t_R _27455_ (.A1(_06491_),
    .A2(_08582_),
    .B(_09071_),
    .C(_09144_),
    .Y(_09145_));
 AOI21x1_ASAP7_75t_R _27456_ (.A1(_01647_),
    .A2(_09067_),
    .B(_09145_),
    .Y(_02751_));
 INVx1_ASAP7_75t_R _27457_ (.A(_01646_),
    .Y(_09146_));
 AO21x1_ASAP7_75t_R _27458_ (.A1(_05474_),
    .A2(_05915_),
    .B(_05369_),
    .Y(_09147_));
 OA211x2_ASAP7_75t_R _27459_ (.A1(net172),
    .A2(_08582_),
    .B(_09071_),
    .C(_09147_),
    .Y(_09148_));
 AO21x1_ASAP7_75t_R _27460_ (.A1(_09146_),
    .A2(_09067_),
    .B(_09148_),
    .Y(_02752_));
 OA211x2_ASAP7_75t_R _27461_ (.A1(net173),
    .A2(_05930_),
    .B(_09071_),
    .C(_05474_),
    .Y(_09149_));
 AO21x1_ASAP7_75t_R _27462_ (.A1(_08677_),
    .A2(_09067_),
    .B(_09149_),
    .Y(_02753_));
 AND3x4_ASAP7_75t_R _27463_ (.A(_06705_),
    .B(_01357_),
    .C(_05757_),
    .Y(_09150_));
 TAPCELL_ASAP7_75t_R TAP_655 ();
 TAPCELL_ASAP7_75t_R TAP_654 ();
 NAND2x2_ASAP7_75t_R _27466_ (.A(_05741_),
    .B(_05757_),
    .Y(_09153_));
 OR2x4_ASAP7_75t_R _27467_ (.A(_01321_),
    .B(_09153_),
    .Y(_09154_));
 OA21x2_ASAP7_75t_R _27468_ (.A1(_08608_),
    .A2(_09154_),
    .B(_01323_),
    .Y(_09155_));
 NOR2x1_ASAP7_75t_R _27469_ (.A(_09150_),
    .B(_09155_),
    .Y(_02754_));
 TAPCELL_ASAP7_75t_R TAP_653 ();
 OA21x2_ASAP7_75t_R _27471_ (.A1(_08708_),
    .A2(_09153_),
    .B(_01324_),
    .Y(_09157_));
 NOR2x1_ASAP7_75t_R _27472_ (.A(_09150_),
    .B(_09157_),
    .Y(_02755_));
 OR2x6_ASAP7_75t_R _27473_ (.A(_01326_),
    .B(_09153_),
    .Y(_09158_));
 TAPCELL_ASAP7_75t_R TAP_652 ();
 OA21x2_ASAP7_75t_R _27475_ (.A1(_08608_),
    .A2(_09158_),
    .B(_01325_),
    .Y(_09160_));
 NOR2x1_ASAP7_75t_R _27476_ (.A(_09150_),
    .B(_09160_),
    .Y(_02756_));
 TAPCELL_ASAP7_75t_R TAP_651 ();
 OR2x6_ASAP7_75t_R _27478_ (.A(_01320_),
    .B(_09153_),
    .Y(_09162_));
 TAPCELL_ASAP7_75t_R TAP_650 ();
 OAI22x1_ASAP7_75t_R _27480_ (.A1(_01327_),
    .A2(_09150_),
    .B1(_09162_),
    .B2(_08608_),
    .Y(_02757_));
 OA21x2_ASAP7_75t_R _27481_ (.A1(_08750_),
    .A2(_09154_),
    .B(_01328_),
    .Y(_09164_));
 NOR2x1_ASAP7_75t_R _27482_ (.A(_09150_),
    .B(_09164_),
    .Y(_02758_));
 OR4x1_ASAP7_75t_R _27483_ (.A(_08746_),
    .B(_05752_),
    .C(_08748_),
    .D(_09153_),
    .Y(_09165_));
 AOI21x1_ASAP7_75t_R _27484_ (.A1(_01329_),
    .A2(_09165_),
    .B(_09150_),
    .Y(_02759_));
 OAI22x1_ASAP7_75t_R _27485_ (.A1(_01330_),
    .A2(_09150_),
    .B1(_09158_),
    .B2(_08750_),
    .Y(_02760_));
 OAI22x1_ASAP7_75t_R _27486_ (.A1(_01331_),
    .A2(_09150_),
    .B1(_09162_),
    .B2(_08750_),
    .Y(_02761_));
 OA21x2_ASAP7_75t_R _27487_ (.A1(_08808_),
    .A2(_09154_),
    .B(_01332_),
    .Y(_09166_));
 NOR2x1_ASAP7_75t_R _27488_ (.A(_09150_),
    .B(_09166_),
    .Y(_02762_));
 OA21x2_ASAP7_75t_R _27489_ (.A1(_08820_),
    .A2(_09153_),
    .B(_01333_),
    .Y(_09167_));
 NOR2x1_ASAP7_75t_R _27490_ (.A(_09150_),
    .B(_09167_),
    .Y(_02763_));
 TAPCELL_ASAP7_75t_R TAP_649 ();
 OAI22x1_ASAP7_75t_R _27492_ (.A1(_01334_),
    .A2(_09150_),
    .B1(_09158_),
    .B2(_08808_),
    .Y(_02764_));
 OAI22x1_ASAP7_75t_R _27493_ (.A1(_01335_),
    .A2(_09150_),
    .B1(_09162_),
    .B2(_08808_),
    .Y(_02765_));
 OR3x2_ASAP7_75t_R _27494_ (.A(_01321_),
    .B(_08748_),
    .C(_09153_),
    .Y(_09169_));
 OAI22x1_ASAP7_75t_R _27495_ (.A1(_01336_),
    .A2(_09150_),
    .B1(_09169_),
    .B2(_08807_),
    .Y(_02766_));
 OR4x1_ASAP7_75t_R _27496_ (.A(_01322_),
    .B(_05752_),
    .C(_08748_),
    .D(_09153_),
    .Y(_09170_));
 AOI21x1_ASAP7_75t_R _27497_ (.A1(_01337_),
    .A2(_09170_),
    .B(_09150_),
    .Y(_02767_));
 OAI22x1_ASAP7_75t_R _27498_ (.A1(_01338_),
    .A2(_09150_),
    .B1(_09158_),
    .B2(_08873_),
    .Y(_02768_));
 OAI22x1_ASAP7_75t_R _27499_ (.A1(_01339_),
    .A2(_09150_),
    .B1(_09162_),
    .B2(_08873_),
    .Y(_02769_));
 OAI22x1_ASAP7_75t_R _27500_ (.A1(_01340_),
    .A2(_09150_),
    .B1(_09154_),
    .B2(_08894_),
    .Y(_02770_));
 OR5x1_ASAP7_75t_R _27501_ (.A(_01319_),
    .B(_01318_),
    .C(_05750_),
    .D(_08607_),
    .E(_09153_),
    .Y(_09171_));
 AOI21x1_ASAP7_75t_R _27502_ (.A1(_01341_),
    .A2(_09171_),
    .B(_09150_),
    .Y(_02771_));
 OAI22x1_ASAP7_75t_R _27503_ (.A1(_01342_),
    .A2(_09150_),
    .B1(_09158_),
    .B2(_08894_),
    .Y(_02772_));
 OAI22x1_ASAP7_75t_R _27504_ (.A1(_01343_),
    .A2(_09150_),
    .B1(_09162_),
    .B2(_08894_),
    .Y(_02773_));
 OAI22x1_ASAP7_75t_R _27505_ (.A1(_01344_),
    .A2(_09150_),
    .B1(_09169_),
    .B2(_08933_),
    .Y(_02774_));
 OR5x1_ASAP7_75t_R _27506_ (.A(_01319_),
    .B(_01318_),
    .C(_08746_),
    .D(_08748_),
    .E(_09153_),
    .Y(_09172_));
 OAI21x1_ASAP7_75t_R _27507_ (.A1(_01345_),
    .A2(_09150_),
    .B(_09172_),
    .Y(_02775_));
 OAI22x1_ASAP7_75t_R _27508_ (.A1(_01346_),
    .A2(_09150_),
    .B1(_09158_),
    .B2(_08953_),
    .Y(_02776_));
 OAI22x1_ASAP7_75t_R _27509_ (.A1(_01347_),
    .A2(_09150_),
    .B1(_09162_),
    .B2(_08953_),
    .Y(_02777_));
 OAI22x1_ASAP7_75t_R _27510_ (.A1(_01348_),
    .A2(_09150_),
    .B1(_09154_),
    .B2(_08975_),
    .Y(_02778_));
 OR3x1_ASAP7_75t_R _27511_ (.A(_08819_),
    .B(_08985_),
    .C(_09153_),
    .Y(_09173_));
 AOI21x1_ASAP7_75t_R _27512_ (.A1(_01349_),
    .A2(_09173_),
    .B(_09150_),
    .Y(_02779_));
 OAI22x1_ASAP7_75t_R _27513_ (.A1(_01350_),
    .A2(_09150_),
    .B1(_09158_),
    .B2(_08975_),
    .Y(_02780_));
 OAI22x1_ASAP7_75t_R _27514_ (.A1(_01351_),
    .A2(_09150_),
    .B1(_09162_),
    .B2(_08975_),
    .Y(_02781_));
 OR3x1_ASAP7_75t_R _27515_ (.A(_01318_),
    .B(_01322_),
    .C(_09169_),
    .Y(_09174_));
 OAI21x1_ASAP7_75t_R _27516_ (.A1(_01352_),
    .A2(_09150_),
    .B(_09174_),
    .Y(_02782_));
 OR3x1_ASAP7_75t_R _27517_ (.A(_08748_),
    .B(_08985_),
    .C(_09153_),
    .Y(_09175_));
 AOI21x1_ASAP7_75t_R _27518_ (.A1(_01353_),
    .A2(_09175_),
    .B(_09150_),
    .Y(_02783_));
 OAI22x1_ASAP7_75t_R _27519_ (.A1(_01354_),
    .A2(_09150_),
    .B1(_09158_),
    .B2(_09013_),
    .Y(_02784_));
 OAI22x1_ASAP7_75t_R _27520_ (.A1(_01355_),
    .A2(_09150_),
    .B1(_09162_),
    .B2(_09013_),
    .Y(_02785_));
 AND3x4_ASAP7_75t_R _27521_ (.A(_00284_),
    .B(_01872_),
    .C(_01873_),
    .Y(_09176_));
 AND3x1_ASAP7_75t_R _27522_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_05757_),
    .C(_09176_),
    .Y(_09177_));
 AOI21x1_ASAP7_75t_R _27523_ (.A1(_17600_),
    .A2(_05747_),
    .B(_09177_),
    .Y(_02786_));
 AND3x1_ASAP7_75t_R _27524_ (.A(_08621_),
    .B(_05757_),
    .C(_09176_),
    .Y(_09178_));
 AOI21x1_ASAP7_75t_R _27525_ (.A1(_17601_),
    .A2(_05747_),
    .B(_09178_),
    .Y(_02787_));
 AND3x1_ASAP7_75t_R _27526_ (.A(_08660_),
    .B(_05757_),
    .C(_09176_),
    .Y(_09179_));
 AOI21x1_ASAP7_75t_R _27527_ (.A1(_17607_),
    .A2(_05747_),
    .B(_09179_),
    .Y(_02788_));
 AND3x1_ASAP7_75t_R _27528_ (.A(_05757_),
    .B(_08629_),
    .C(_09176_),
    .Y(_09180_));
 AOI21x1_ASAP7_75t_R _27529_ (.A1(_01322_),
    .A2(_05747_),
    .B(_09180_),
    .Y(_02789_));
 OA21x2_ASAP7_75t_R _27530_ (.A1(_02291_),
    .A2(_05750_),
    .B(_09176_),
    .Y(_09181_));
 OA21x2_ASAP7_75t_R _27531_ (.A1(_05747_),
    .A2(_09181_),
    .B(_01318_),
    .Y(_09182_));
 AND4x1_ASAP7_75t_R _27532_ (.A(_05751_),
    .B(_05757_),
    .C(_08657_),
    .D(_09176_),
    .Y(_09183_));
 NOR2x1_ASAP7_75t_R _27533_ (.A(_09182_),
    .B(_09183_),
    .Y(_02790_));
 NAND2x1_ASAP7_75t_R _27534_ (.A(_01316_),
    .B(_05733_),
    .Y(_09184_));
 OA21x2_ASAP7_75t_R _27535_ (.A1(_05733_),
    .A2(net218),
    .B(_09184_),
    .Y(_02791_));
 INVx1_ASAP7_75t_R _27536_ (.A(_01644_),
    .Y(_09185_));
 AND4x1_ASAP7_75t_R _27537_ (.A(_00279_),
    .B(_00175_),
    .C(_14615_),
    .D(_05734_),
    .Y(_09186_));
 AO21x1_ASAP7_75t_R _27538_ (.A1(_09185_),
    .A2(_05733_),
    .B(_09186_),
    .Y(_02792_));
 OR2x2_ASAP7_75t_R _27539_ (.A(\ex_block_i.alu_adder_result_ex_o[0] ),
    .B(_05733_),
    .Y(_09187_));
 OA21x2_ASAP7_75t_R _27540_ (.A1(_07135_),
    .A2(_05734_),
    .B(_09187_),
    .Y(_02793_));
 OR2x2_ASAP7_75t_R _27541_ (.A(net279),
    .B(_05733_),
    .Y(_09188_));
 OA21x2_ASAP7_75t_R _27542_ (.A1(_07120_),
    .A2(_05734_),
    .B(_09188_),
    .Y(_02794_));
 INVx1_ASAP7_75t_R _27543_ (.A(_01607_),
    .Y(_09189_));
 AO21x1_ASAP7_75t_R _27544_ (.A1(_09189_),
    .A2(_13284_),
    .B(_01609_),
    .Y(_09190_));
 NAND2x1_ASAP7_75t_R _27545_ (.A(_05731_),
    .B(_09190_),
    .Y(_09191_));
 AND3x1_ASAP7_75t_R _27546_ (.A(net59),
    .B(_05523_),
    .C(_01609_),
    .Y(_09192_));
 NOR2x1_ASAP7_75t_R _27547_ (.A(_01608_),
    .B(_05732_),
    .Y(_09193_));
 AO21x1_ASAP7_75t_R _27548_ (.A1(_13221_),
    .A2(_01608_),
    .B(_09193_),
    .Y(_09194_));
 AO32x2_ASAP7_75t_R _27549_ (.A1(_00277_),
    .A2(net26),
    .A3(_09191_),
    .B1(_09192_),
    .B2(_09194_),
    .Y(_09195_));
 TAPCELL_ASAP7_75t_R TAP_648 ();
 TAPCELL_ASAP7_75t_R TAP_647 ();
 TAPCELL_ASAP7_75t_R TAP_646 ();
 NOR2x1_ASAP7_75t_R _27553_ (.A(_01641_),
    .B(_09195_),
    .Y(_09199_));
 AO21x1_ASAP7_75t_R _27554_ (.A1(\ex_block_i.alu_adder_result_ex_o[0] ),
    .A2(_09195_),
    .B(_09199_),
    .Y(_02795_));
 NOR2x1_ASAP7_75t_R _27555_ (.A(_01640_),
    .B(_09195_),
    .Y(_09200_));
 AO21x1_ASAP7_75t_R _27556_ (.A1(net279),
    .A2(_09195_),
    .B(_09200_),
    .Y(_02796_));
 TAPCELL_ASAP7_75t_R TAP_645 ();
 NOR2x1_ASAP7_75t_R _27558_ (.A(_01639_),
    .B(_09195_),
    .Y(_09202_));
 AO21x1_ASAP7_75t_R _27559_ (.A1(net171),
    .A2(_09195_),
    .B(_09202_),
    .Y(_02797_));
 NOR2x1_ASAP7_75t_R _27560_ (.A(_01638_),
    .B(_09195_),
    .Y(_09203_));
 AO21x1_ASAP7_75t_R _27561_ (.A1(net275),
    .A2(_09195_),
    .B(_09203_),
    .Y(_02798_));
 NOR2x1_ASAP7_75t_R _27562_ (.A(_01637_),
    .B(_09195_),
    .Y(_09204_));
 AO21x1_ASAP7_75t_R _27563_ (.A1(net175),
    .A2(_09195_),
    .B(_09204_),
    .Y(_02799_));
 NOR2x1_ASAP7_75t_R _27564_ (.A(_01636_),
    .B(_09195_),
    .Y(_09205_));
 AO21x1_ASAP7_75t_R _27565_ (.A1(net176),
    .A2(_09195_),
    .B(_09205_),
    .Y(_02800_));
 NOR2x1_ASAP7_75t_R _27566_ (.A(_01635_),
    .B(_09195_),
    .Y(_09206_));
 AO21x1_ASAP7_75t_R _27567_ (.A1(net177),
    .A2(_09195_),
    .B(_09206_),
    .Y(_02801_));
 TAPCELL_ASAP7_75t_R TAP_644 ();
 NAND2x1_ASAP7_75t_R _27569_ (.A(_00676_),
    .B(_09195_),
    .Y(_09208_));
 OA21x2_ASAP7_75t_R _27570_ (.A1(_14991_),
    .A2(_09195_),
    .B(_09208_),
    .Y(_02802_));
 NAND2x1_ASAP7_75t_R _27571_ (.A(_05773_),
    .B(_09195_),
    .Y(_09209_));
 OA21x2_ASAP7_75t_R _27572_ (.A1(_14995_),
    .A2(_09195_),
    .B(_09209_),
    .Y(_02803_));
 NOR2x1_ASAP7_75t_R _27573_ (.A(_01632_),
    .B(_09195_),
    .Y(_09210_));
 AO21x1_ASAP7_75t_R _27574_ (.A1(net180),
    .A2(_09195_),
    .B(_09210_),
    .Y(_02804_));
 NOR2x1_ASAP7_75t_R _27575_ (.A(_01631_),
    .B(_09195_),
    .Y(_09211_));
 AO21x1_ASAP7_75t_R _27576_ (.A1(net151),
    .A2(_09195_),
    .B(_09211_),
    .Y(_02805_));
 NOR2x1_ASAP7_75t_R _27577_ (.A(_01630_),
    .B(_09195_),
    .Y(_09212_));
 AO21x1_ASAP7_75t_R _27578_ (.A1(net152),
    .A2(_09195_),
    .B(_09212_),
    .Y(_02806_));
 TAPCELL_ASAP7_75t_R TAP_643 ();
 NOR2x1_ASAP7_75t_R _27580_ (.A(_01629_),
    .B(_09195_),
    .Y(_09214_));
 AO21x1_ASAP7_75t_R _27581_ (.A1(net153),
    .A2(_09195_),
    .B(_09214_),
    .Y(_02807_));
 NOR2x1_ASAP7_75t_R _27582_ (.A(_01628_),
    .B(_09195_),
    .Y(_09215_));
 AO21x1_ASAP7_75t_R _27583_ (.A1(net154),
    .A2(_09195_),
    .B(_09215_),
    .Y(_02808_));
 TAPCELL_ASAP7_75t_R TAP_642 ();
 NOR2x1_ASAP7_75t_R _27585_ (.A(_01627_),
    .B(_09195_),
    .Y(_09217_));
 AO21x1_ASAP7_75t_R _27586_ (.A1(net155),
    .A2(_09195_),
    .B(_09217_),
    .Y(_02809_));
 NAND2x1_ASAP7_75t_R _27587_ (.A(net256),
    .B(_09195_),
    .Y(_09218_));
 OA21x2_ASAP7_75t_R _27588_ (.A1(_15621_),
    .A2(_09195_),
    .B(_09218_),
    .Y(_02810_));
 NAND2x1_ASAP7_75t_R _27589_ (.A(_05770_),
    .B(_09195_),
    .Y(_09219_));
 OA21x2_ASAP7_75t_R _27590_ (.A1(_15733_),
    .A2(_09195_),
    .B(_09219_),
    .Y(_02811_));
 NOR2x1_ASAP7_75t_R _27591_ (.A(_01624_),
    .B(_09195_),
    .Y(_09220_));
 AO21x1_ASAP7_75t_R _27592_ (.A1(net158),
    .A2(_09195_),
    .B(_09220_),
    .Y(_02812_));
 NOR2x1_ASAP7_75t_R _27593_ (.A(_01623_),
    .B(_09195_),
    .Y(_09221_));
 AO21x1_ASAP7_75t_R _27594_ (.A1(net159),
    .A2(_09195_),
    .B(_09221_),
    .Y(_02813_));
 NOR2x1_ASAP7_75t_R _27595_ (.A(_01622_),
    .B(_09195_),
    .Y(_09222_));
 AO21x1_ASAP7_75t_R _27596_ (.A1(net257),
    .A2(_09195_),
    .B(_09222_),
    .Y(_02814_));
 NOR2x1_ASAP7_75t_R _27597_ (.A(_01621_),
    .B(_09195_),
    .Y(_09223_));
 AO21x1_ASAP7_75t_R _27598_ (.A1(net161),
    .A2(_09195_),
    .B(_09223_),
    .Y(_02815_));
 NOR2x1_ASAP7_75t_R _27599_ (.A(_01620_),
    .B(_09195_),
    .Y(_09224_));
 AO21x1_ASAP7_75t_R _27600_ (.A1(net255),
    .A2(_09195_),
    .B(_09224_),
    .Y(_02816_));
 INVx1_ASAP7_75t_R _27601_ (.A(_01619_),
    .Y(_09225_));
 NAND2x1_ASAP7_75t_R _27602_ (.A(_05760_),
    .B(_09195_),
    .Y(_09226_));
 OA21x2_ASAP7_75t_R _27603_ (.A1(_09225_),
    .A2(_09195_),
    .B(_09226_),
    .Y(_02817_));
 NOR2x1_ASAP7_75t_R _27604_ (.A(_01618_),
    .B(_09195_),
    .Y(_09227_));
 AO21x1_ASAP7_75t_R _27605_ (.A1(net164),
    .A2(_09195_),
    .B(_09227_),
    .Y(_02818_));
 NOR2x1_ASAP7_75t_R _27606_ (.A(_01617_),
    .B(_09195_),
    .Y(_09228_));
 AO21x1_ASAP7_75t_R _27607_ (.A1(net165),
    .A2(_09195_),
    .B(_09228_),
    .Y(_02819_));
 NOR2x1_ASAP7_75t_R _27608_ (.A(_01616_),
    .B(_09195_),
    .Y(_09229_));
 AO21x1_ASAP7_75t_R _27609_ (.A1(net166),
    .A2(_09195_),
    .B(_09229_),
    .Y(_02820_));
 INVx1_ASAP7_75t_R _27610_ (.A(_01615_),
    .Y(_09230_));
 NAND2x1_ASAP7_75t_R _27611_ (.A(_04937_),
    .B(_09195_),
    .Y(_09231_));
 OA21x2_ASAP7_75t_R _27612_ (.A1(_09230_),
    .A2(_09195_),
    .B(_09231_),
    .Y(_02821_));
 NOR2x1_ASAP7_75t_R _27613_ (.A(_01614_),
    .B(_09195_),
    .Y(_09232_));
 AO21x1_ASAP7_75t_R _27614_ (.A1(net168),
    .A2(_09195_),
    .B(_09232_),
    .Y(_02822_));
 INVx1_ASAP7_75t_R _27615_ (.A(_01613_),
    .Y(_09233_));
 NAND2x1_ASAP7_75t_R _27616_ (.A(_05154_),
    .B(_09195_),
    .Y(_09234_));
 OA21x2_ASAP7_75t_R _27617_ (.A1(_09233_),
    .A2(_09195_),
    .B(_09234_),
    .Y(_02823_));
 NOR2x1_ASAP7_75t_R _27618_ (.A(_01612_),
    .B(_09195_),
    .Y(_09235_));
 AO21x1_ASAP7_75t_R _27619_ (.A1(net2116),
    .A2(_09195_),
    .B(_09235_),
    .Y(_02824_));
 NAND2x1_ASAP7_75t_R _27620_ (.A(_05372_),
    .B(_09195_),
    .Y(_09236_));
 OA21x2_ASAP7_75t_R _27621_ (.A1(_05326_),
    .A2(_09195_),
    .B(_09236_),
    .Y(_02825_));
 NOR2x1_ASAP7_75t_R _27622_ (.A(_01610_),
    .B(_09195_),
    .Y(_09237_));
 AO21x1_ASAP7_75t_R _27623_ (.A1(net173),
    .A2(_09195_),
    .B(_09237_),
    .Y(_02826_));
 INVx1_ASAP7_75t_R _27624_ (.A(net59),
    .Y(_09238_));
 OAI21x1_ASAP7_75t_R _27625_ (.A1(_09238_),
    .A2(_01608_),
    .B(_05731_),
    .Y(_09239_));
 INVx1_ASAP7_75t_R _27626_ (.A(net26),
    .Y(_09240_));
 OA211x2_ASAP7_75t_R _27627_ (.A1(_13220_),
    .A2(_09239_),
    .B(_00277_),
    .C(_09240_),
    .Y(_02827_));
 INVx1_ASAP7_75t_R _27628_ (.A(_05730_),
    .Y(_09241_));
 OA21x2_ASAP7_75t_R _27629_ (.A1(_00281_),
    .A2(_02537_),
    .B(_05739_),
    .Y(_09242_));
 AO21x1_ASAP7_75t_R _27630_ (.A1(_06070_),
    .A2(_06148_),
    .B(_09242_),
    .Y(_09243_));
 NAND2x1_ASAP7_75t_R _27631_ (.A(_01609_),
    .B(_09243_),
    .Y(_09244_));
 OA21x2_ASAP7_75t_R _27632_ (.A1(_09241_),
    .A2(_09244_),
    .B(_01608_),
    .Y(_09245_));
 NOR2x1_ASAP7_75t_R _27633_ (.A(net26),
    .B(_09245_),
    .Y(_09246_));
 AND3x1_ASAP7_75t_R _27634_ (.A(net26),
    .B(_01608_),
    .C(_09244_),
    .Y(_09247_));
 OA21x2_ASAP7_75t_R _27635_ (.A1(_13220_),
    .A2(_05730_),
    .B(_09247_),
    .Y(_09248_));
 OA21x2_ASAP7_75t_R _27636_ (.A1(_09246_),
    .A2(_09248_),
    .B(_00277_),
    .Y(_02828_));
 AND3x1_ASAP7_75t_R _27637_ (.A(_09238_),
    .B(_01609_),
    .C(_09194_),
    .Y(_02829_));
 AND3x1_ASAP7_75t_R _27638_ (.A(_13221_),
    .B(net59),
    .C(_01608_),
    .Y(_09249_));
 AO21x1_ASAP7_75t_R _27639_ (.A1(_00277_),
    .A2(_09239_),
    .B(_09249_),
    .Y(_09250_));
 NAND2x1_ASAP7_75t_R _27640_ (.A(_01609_),
    .B(_09250_),
    .Y(_09251_));
 AND4x1_ASAP7_75t_R _27641_ (.A(net25),
    .B(_01609_),
    .C(_13645_),
    .D(_09250_),
    .Y(_09252_));
 AO21x1_ASAP7_75t_R _27642_ (.A1(_09189_),
    .A2(_09251_),
    .B(_09252_),
    .Y(_02830_));
 AO32x1_ASAP7_75t_R _27643_ (.A1(net59),
    .A2(_13284_),
    .A3(_01609_),
    .B1(_06161_),
    .B2(net26),
    .Y(_09253_));
 AO21x1_ASAP7_75t_R _27644_ (.A1(_00277_),
    .A2(_09253_),
    .B(_13283_),
    .Y(_09254_));
 OA21x2_ASAP7_75t_R _27645_ (.A1(_05732_),
    .A2(_09245_),
    .B(_09254_),
    .Y(_02831_));
 OA222x2_ASAP7_75t_R _27646_ (.A1(_16499_),
    .A2(_06266_),
    .B1(_06262_),
    .B2(_01944_),
    .C1(_06258_),
    .C2(_00658_),
    .Y(_09255_));
 AND2x2_ASAP7_75t_R _27647_ (.A(_06536_),
    .B(_06540_),
    .Y(_09256_));
 AND3x4_ASAP7_75t_R _27648_ (.A(_06558_),
    .B(_06606_),
    .C(_06625_),
    .Y(_09257_));
 TAPCELL_ASAP7_75t_R TAP_641 ();
 TAPCELL_ASAP7_75t_R TAP_640 ();
 TAPCELL_ASAP7_75t_R TAP_639 ();
 TAPCELL_ASAP7_75t_R TAP_638 ();
 TAPCELL_ASAP7_75t_R TAP_637 ();
 AO21x1_ASAP7_75t_R _27654_ (.A1(_09256_),
    .A2(_09257_),
    .B(_00662_),
    .Y(_09263_));
 TAPCELL_ASAP7_75t_R TAP_636 ();
 TAPCELL_ASAP7_75t_R TAP_635 ();
 AOI21x1_ASAP7_75t_R _27657_ (.A1(_06664_),
    .A2(_09257_),
    .B(_06254_),
    .Y(_09266_));
 AOI22x1_ASAP7_75t_R _27658_ (.A1(_06254_),
    .A2(_09255_),
    .B1(_09263_),
    .B2(_09266_),
    .Y(_02832_));
 NAND2x1_ASAP7_75t_R _27659_ (.A(_00241_),
    .B(_09257_),
    .Y(_09267_));
 OA211x2_ASAP7_75t_R _27660_ (.A1(_17536_),
    .A2(_09257_),
    .B(_09267_),
    .C(net287),
    .Y(_09268_));
 NOR2x1_ASAP7_75t_R _27661_ (.A(_06271_),
    .B(_09268_),
    .Y(_02833_));
 TAPCELL_ASAP7_75t_R TAP_634 ();
 OR3x4_ASAP7_75t_R _27663_ (.A(_06655_),
    .B(_06656_),
    .C(_06624_),
    .Y(_09270_));
 TAPCELL_ASAP7_75t_R TAP_633 ();
 TAPCELL_ASAP7_75t_R TAP_632 ();
 TAPCELL_ASAP7_75t_R TAP_631 ();
 TAPCELL_ASAP7_75t_R TAP_630 ();
 AND2x2_ASAP7_75t_R _27668_ (.A(_02539_),
    .B(_09257_),
    .Y(_09275_));
 AO21x1_ASAP7_75t_R _27669_ (.A1(_01606_),
    .A2(_09270_),
    .B(_09275_),
    .Y(_09276_));
 AOI21x1_ASAP7_75t_R _27670_ (.A1(net287),
    .A2(_09276_),
    .B(_06291_),
    .Y(_02834_));
 OR2x2_ASAP7_75t_R _27671_ (.A(_02538_),
    .B(_09270_),
    .Y(_09277_));
 XNOR2x1_ASAP7_75t_R _27672_ (.B(_09277_),
    .Y(_09278_),
    .A(_01605_));
 AOI21x1_ASAP7_75t_R _27673_ (.A1(net287),
    .A2(_09278_),
    .B(_06302_),
    .Y(_02835_));
 AND2x2_ASAP7_75t_R _27674_ (.A(_02541_),
    .B(_09257_),
    .Y(_09279_));
 AO21x1_ASAP7_75t_R _27675_ (.A1(_01604_),
    .A2(_09270_),
    .B(_09279_),
    .Y(_09280_));
 AOI21x1_ASAP7_75t_R _27676_ (.A1(net287),
    .A2(_09280_),
    .B(_06310_),
    .Y(_02836_));
 OR2x2_ASAP7_75t_R _27677_ (.A(_02540_),
    .B(_09270_),
    .Y(_09281_));
 XNOR2x1_ASAP7_75t_R _27678_ (.B(_09281_),
    .Y(_09282_),
    .A(_01603_));
 AOI21x1_ASAP7_75t_R _27679_ (.A1(net287),
    .A2(_09282_),
    .B(_06320_),
    .Y(_02837_));
 AND2x2_ASAP7_75t_R _27680_ (.A(_02543_),
    .B(_09257_),
    .Y(_09283_));
 AO21x1_ASAP7_75t_R _27681_ (.A1(_01602_),
    .A2(_09270_),
    .B(_09283_),
    .Y(_09284_));
 AOI21x1_ASAP7_75t_R _27682_ (.A1(net287),
    .A2(_09284_),
    .B(_06333_),
    .Y(_02838_));
 NOR2x1_ASAP7_75t_R _27683_ (.A(_02542_),
    .B(_09270_),
    .Y(_09285_));
 XNOR2x1_ASAP7_75t_R _27684_ (.B(_09285_),
    .Y(_09286_),
    .A(_01601_));
 AO21x1_ASAP7_75t_R _27685_ (.A1(net287),
    .A2(_09286_),
    .B(_06347_),
    .Y(_02839_));
 TAPCELL_ASAP7_75t_R TAP_629 ();
 NAND2x1_ASAP7_75t_R _27687_ (.A(_02545_),
    .B(_09257_),
    .Y(_09288_));
 OA21x2_ASAP7_75t_R _27688_ (.A1(\cs_registers_i.pc_if_i[9] ),
    .A2(_09257_),
    .B(_09288_),
    .Y(_09289_));
 AO21x1_ASAP7_75t_R _27689_ (.A1(net287),
    .A2(_09289_),
    .B(_06355_),
    .Y(_02840_));
 OR2x2_ASAP7_75t_R _27690_ (.A(_02544_),
    .B(_09270_),
    .Y(_09290_));
 XNOR2x1_ASAP7_75t_R _27691_ (.B(_09290_),
    .Y(_09291_),
    .A(_01599_));
 AOI21x1_ASAP7_75t_R _27692_ (.A1(net287),
    .A2(_09291_),
    .B(_06362_),
    .Y(_02841_));
 TAPCELL_ASAP7_75t_R TAP_628 ();
 AND2x2_ASAP7_75t_R _27694_ (.A(_02547_),
    .B(_09257_),
    .Y(_09293_));
 AO21x1_ASAP7_75t_R _27695_ (.A1(_01598_),
    .A2(_09270_),
    .B(_09293_),
    .Y(_09294_));
 OAI21x1_ASAP7_75t_R _27696_ (.A1(_06254_),
    .A2(_09294_),
    .B(_06375_),
    .Y(_02842_));
 OR2x2_ASAP7_75t_R _27697_ (.A(_02546_),
    .B(_09270_),
    .Y(_09295_));
 XNOR2x1_ASAP7_75t_R _27698_ (.B(_09295_),
    .Y(_09296_),
    .A(_01597_));
 AOI21x1_ASAP7_75t_R _27699_ (.A1(net287),
    .A2(_09296_),
    .B(_06381_),
    .Y(_02843_));
 NAND2x1_ASAP7_75t_R _27700_ (.A(_02549_),
    .B(_09257_),
    .Y(_09297_));
 OA21x2_ASAP7_75t_R _27701_ (.A1(\cs_registers_i.pc_if_i[13] ),
    .A2(_09257_),
    .B(_09297_),
    .Y(_09298_));
 AO21x1_ASAP7_75t_R _27702_ (.A1(net287),
    .A2(_09298_),
    .B(_06389_),
    .Y(_02844_));
 OR2x2_ASAP7_75t_R _27703_ (.A(_02548_),
    .B(_09270_),
    .Y(_09299_));
 XNOR2x1_ASAP7_75t_R _27704_ (.B(_09299_),
    .Y(_09300_),
    .A(_01595_));
 AOI21x1_ASAP7_75t_R _27705_ (.A1(net287),
    .A2(_09300_),
    .B(_06395_),
    .Y(_02845_));
 AND2x2_ASAP7_75t_R _27706_ (.A(_02551_),
    .B(_09257_),
    .Y(_09301_));
 AO21x1_ASAP7_75t_R _27707_ (.A1(_01594_),
    .A2(_09270_),
    .B(_09301_),
    .Y(_09302_));
 AOI21x1_ASAP7_75t_R _27708_ (.A1(net286),
    .A2(_09302_),
    .B(_06400_),
    .Y(_02846_));
 OR2x2_ASAP7_75t_R _27709_ (.A(_02550_),
    .B(_09270_),
    .Y(_09303_));
 XNOR2x1_ASAP7_75t_R _27710_ (.B(_09303_),
    .Y(_09304_),
    .A(_01593_));
 AOI21x1_ASAP7_75t_R _27711_ (.A1(net286),
    .A2(_09304_),
    .B(_06409_),
    .Y(_02847_));
 TAPCELL_ASAP7_75t_R TAP_627 ();
 AND2x2_ASAP7_75t_R _27713_ (.A(_02553_),
    .B(_09257_),
    .Y(_09306_));
 AO21x1_ASAP7_75t_R _27714_ (.A1(_01592_),
    .A2(_09270_),
    .B(_09306_),
    .Y(_09307_));
 AOI21x1_ASAP7_75t_R _27715_ (.A1(net286),
    .A2(_09307_),
    .B(_06415_),
    .Y(_02848_));
 TAPCELL_ASAP7_75t_R TAP_626 ();
 OAI21x1_ASAP7_75t_R _27717_ (.A1(_02552_),
    .A2(_09270_),
    .B(_01591_),
    .Y(_09309_));
 OR3x1_ASAP7_75t_R _27718_ (.A(_01591_),
    .B(_02552_),
    .C(_09270_),
    .Y(_09310_));
 AND3x1_ASAP7_75t_R _27719_ (.A(net286),
    .B(_09309_),
    .C(_09310_),
    .Y(_09311_));
 AO21x1_ASAP7_75t_R _27720_ (.A1(_06254_),
    .A2(_06422_),
    .B(_09311_),
    .Y(_02849_));
 AND2x2_ASAP7_75t_R _27721_ (.A(_02555_),
    .B(_09257_),
    .Y(_09312_));
 AO21x1_ASAP7_75t_R _27722_ (.A1(_01590_),
    .A2(_09270_),
    .B(_09312_),
    .Y(_09313_));
 AOI21x1_ASAP7_75t_R _27723_ (.A1(net286),
    .A2(_09313_),
    .B(_06429_),
    .Y(_02850_));
 OR2x2_ASAP7_75t_R _27724_ (.A(_02554_),
    .B(_09270_),
    .Y(_09314_));
 XNOR2x1_ASAP7_75t_R _27725_ (.B(_09314_),
    .Y(_09315_),
    .A(_01589_));
 AOI21x1_ASAP7_75t_R _27726_ (.A1(net286),
    .A2(_09315_),
    .B(_06436_),
    .Y(_02851_));
 AND2x2_ASAP7_75t_R _27727_ (.A(_02557_),
    .B(_09257_),
    .Y(_09316_));
 AO21x1_ASAP7_75t_R _27728_ (.A1(_01588_),
    .A2(_09270_),
    .B(_09316_),
    .Y(_09317_));
 AOI21x1_ASAP7_75t_R _27729_ (.A1(net286),
    .A2(_09317_),
    .B(_06443_),
    .Y(_02852_));
 OR2x2_ASAP7_75t_R _27730_ (.A(_02556_),
    .B(_09270_),
    .Y(_09318_));
 XNOR2x1_ASAP7_75t_R _27731_ (.B(_09318_),
    .Y(_09319_),
    .A(_01587_));
 AOI21x1_ASAP7_75t_R _27732_ (.A1(net286),
    .A2(_09319_),
    .B(_06449_),
    .Y(_02853_));
 AND2x2_ASAP7_75t_R _27733_ (.A(_02559_),
    .B(_09257_),
    .Y(_09320_));
 AO21x1_ASAP7_75t_R _27734_ (.A1(_01586_),
    .A2(_09270_),
    .B(_09320_),
    .Y(_09321_));
 AOI21x1_ASAP7_75t_R _27735_ (.A1(net286),
    .A2(_09321_),
    .B(_06455_),
    .Y(_02854_));
 OR2x2_ASAP7_75t_R _27736_ (.A(_02558_),
    .B(_09270_),
    .Y(_09322_));
 XNOR2x1_ASAP7_75t_R _27737_ (.B(_09322_),
    .Y(_09323_),
    .A(_01585_));
 AOI21x1_ASAP7_75t_R _27738_ (.A1(net286),
    .A2(_09323_),
    .B(_06461_),
    .Y(_02855_));
 AND2x2_ASAP7_75t_R _27739_ (.A(_02561_),
    .B(_09257_),
    .Y(_09324_));
 AO21x1_ASAP7_75t_R _27740_ (.A1(_01584_),
    .A2(_09270_),
    .B(_09324_),
    .Y(_09325_));
 AOI21x1_ASAP7_75t_R _27741_ (.A1(net286),
    .A2(_09325_),
    .B(_06468_),
    .Y(_02856_));
 OR2x2_ASAP7_75t_R _27742_ (.A(_02560_),
    .B(_09270_),
    .Y(_09326_));
 XNOR2x1_ASAP7_75t_R _27743_ (.B(_09326_),
    .Y(_09327_),
    .A(_01583_));
 AOI21x1_ASAP7_75t_R _27744_ (.A1(net286),
    .A2(_09327_),
    .B(_06474_),
    .Y(_02857_));
 AND2x2_ASAP7_75t_R _27745_ (.A(_02563_),
    .B(_09257_),
    .Y(_09328_));
 AO21x1_ASAP7_75t_R _27746_ (.A1(_01582_),
    .A2(_09270_),
    .B(_09328_),
    .Y(_09329_));
 AOI21x1_ASAP7_75t_R _27747_ (.A1(net286),
    .A2(_09329_),
    .B(_06481_),
    .Y(_02858_));
 OR2x2_ASAP7_75t_R _27748_ (.A(_02562_),
    .B(_09270_),
    .Y(_09330_));
 XNOR2x1_ASAP7_75t_R _27749_ (.B(_09330_),
    .Y(_09331_),
    .A(_01581_));
 AOI21x1_ASAP7_75t_R _27750_ (.A1(net286),
    .A2(_09331_),
    .B(_06488_),
    .Y(_02859_));
 AND2x2_ASAP7_75t_R _27751_ (.A(_02565_),
    .B(_09257_),
    .Y(_09332_));
 AO21x1_ASAP7_75t_R _27752_ (.A1(_01580_),
    .A2(_09270_),
    .B(_09332_),
    .Y(_09333_));
 AOI21x1_ASAP7_75t_R _27753_ (.A1(net286),
    .A2(_09333_),
    .B(_06494_),
    .Y(_02860_));
 OR2x2_ASAP7_75t_R _27754_ (.A(_02564_),
    .B(_09270_),
    .Y(_09334_));
 XNOR2x1_ASAP7_75t_R _27755_ (.B(_09334_),
    .Y(_09335_),
    .A(_01579_));
 AOI21x1_ASAP7_75t_R _27756_ (.A1(net286),
    .A2(_09335_),
    .B(_06500_),
    .Y(_02861_));
 TAPCELL_ASAP7_75t_R TAP_625 ();
 TAPCELL_ASAP7_75t_R TAP_624 ();
 OR3x1_ASAP7_75t_R _27759_ (.A(_01579_),
    .B(_01580_),
    .C(_06553_),
    .Y(_09338_));
 AO22x1_ASAP7_75t_R _27760_ (.A1(net286),
    .A2(_09270_),
    .B1(_09338_),
    .B2(_06505_),
    .Y(_09339_));
 OR3x1_ASAP7_75t_R _27761_ (.A(_01578_),
    .B(_09270_),
    .C(_09338_),
    .Y(_09340_));
 NAND2x1_ASAP7_75t_R _27762_ (.A(net286),
    .B(_09340_),
    .Y(_09341_));
 AOI22x1_ASAP7_75t_R _27763_ (.A1(_01578_),
    .A2(_09339_),
    .B1(_09341_),
    .B2(_06505_),
    .Y(_02862_));
 INVx1_ASAP7_75t_R _27764_ (.A(_07305_),
    .Y(_09342_));
 AO32x1_ASAP7_75t_R _27765_ (.A1(_05677_),
    .A2(_05624_),
    .A3(_05679_),
    .B1(_05662_),
    .B2(_06894_),
    .Y(_09343_));
 OR4x1_ASAP7_75t_R _27766_ (.A(_06884_),
    .B(_07155_),
    .C(_06886_),
    .D(_09343_),
    .Y(_09344_));
 NAND2x1_ASAP7_75t_R _27767_ (.A(_14140_),
    .B(_07513_),
    .Y(_09345_));
 NAND2x1_ASAP7_75t_R _27768_ (.A(_14139_),
    .B(_06908_),
    .Y(_09346_));
 AND4x1_ASAP7_75t_R _27769_ (.A(_14083_),
    .B(_05538_),
    .C(_09345_),
    .D(_09346_),
    .Y(_09347_));
 OA211x2_ASAP7_75t_R _27770_ (.A1(_05541_),
    .A2(_06899_),
    .B(_05571_),
    .C(_05538_),
    .Y(_09348_));
 OR3x1_ASAP7_75t_R _27771_ (.A(_05628_),
    .B(_05659_),
    .C(_09348_),
    .Y(_09349_));
 OR4x1_ASAP7_75t_R _27772_ (.A(_09347_),
    .B(_06898_),
    .C(_06912_),
    .D(_09349_),
    .Y(_09350_));
 AND4x2_ASAP7_75t_R _27773_ (.A(_02288_),
    .B(_14585_),
    .C(_05535_),
    .D(_06914_),
    .Y(_09351_));
 TAPCELL_ASAP7_75t_R TAP_623 ();
 OA21x2_ASAP7_75t_R _27775_ (.A1(_09344_),
    .A2(_09350_),
    .B(_09351_),
    .Y(_09353_));
 NAND2x2_ASAP7_75t_R _27776_ (.A(_09342_),
    .B(_09353_),
    .Y(_09354_));
 CKINVDCx8_ASAP7_75t_R _27777_ (.A(_09354_),
    .Y(_09355_));
 TAPCELL_ASAP7_75t_R TAP_622 ();
 TAPCELL_ASAP7_75t_R TAP_621 ();
 TAPCELL_ASAP7_75t_R TAP_620 ();
 TAPCELL_ASAP7_75t_R TAP_619 ();
 AND2x2_ASAP7_75t_R _27782_ (.A(_13573_),
    .B(_14501_),
    .Y(_09360_));
 AO21x1_ASAP7_75t_R _27783_ (.A1(_02289_),
    .A2(_18114_),
    .B(_09360_),
    .Y(_09361_));
 AND2x2_ASAP7_75t_R _27784_ (.A(net292),
    .B(_09361_),
    .Y(_09362_));
 AOI21x1_ASAP7_75t_R _27785_ (.A1(_18114_),
    .A2(_07311_),
    .B(_09362_),
    .Y(_09363_));
 OR3x4_ASAP7_75t_R _27786_ (.A(_06896_),
    .B(_06905_),
    .C(_06913_),
    .Y(_09364_));
 AND2x6_ASAP7_75t_R _27787_ (.A(_09364_),
    .B(_09351_),
    .Y(_09365_));
 AND3x4_ASAP7_75t_R _27788_ (.A(_06892_),
    .B(_07515_),
    .C(_09365_),
    .Y(_09366_));
 OR2x6_ASAP7_75t_R _27789_ (.A(_06880_),
    .B(_09366_),
    .Y(_09367_));
 TAPCELL_ASAP7_75t_R TAP_618 ();
 TAPCELL_ASAP7_75t_R TAP_617 ();
 OAI21x1_ASAP7_75t_R _27792_ (.A1(_06184_),
    .A2(_06876_),
    .B(_06224_),
    .Y(_09370_));
 TAPCELL_ASAP7_75t_R TAP_616 ();
 OA21x2_ASAP7_75t_R _27794_ (.A1(_06184_),
    .A2(_06876_),
    .B(_06224_),
    .Y(_09372_));
 TAPCELL_ASAP7_75t_R TAP_615 ();
 AND2x2_ASAP7_75t_R _27796_ (.A(_01720_),
    .B(_09372_),
    .Y(_09374_));
 AO21x1_ASAP7_75t_R _27797_ (.A1(_00662_),
    .A2(_09370_),
    .B(_09374_),
    .Y(_09375_));
 OAI22x1_ASAP7_75t_R _27798_ (.A1(_00658_),
    .A2(_09367_),
    .B1(_09375_),
    .B2(_06873_),
    .Y(_09376_));
 AO21x1_ASAP7_75t_R _27799_ (.A1(_09355_),
    .A2(_09363_),
    .B(_09376_),
    .Y(_02865_));
 TAPCELL_ASAP7_75t_R TAP_614 ();
 TAPCELL_ASAP7_75t_R TAP_613 ();
 AND2x2_ASAP7_75t_R _27802_ (.A(_00162_),
    .B(_09372_),
    .Y(_09379_));
 AO21x2_ASAP7_75t_R _27803_ (.A1(_17536_),
    .A2(_09370_),
    .B(_09379_),
    .Y(_09380_));
 AND2x2_ASAP7_75t_R _27804_ (.A(_02027_),
    .B(_13658_),
    .Y(_09381_));
 AO21x1_ASAP7_75t_R _27805_ (.A1(_01911_),
    .A2(net289),
    .B(_09381_),
    .Y(_09382_));
 OR5x1_ASAP7_75t_R _27806_ (.A(_13301_),
    .B(_13954_),
    .C(_05560_),
    .D(_07507_),
    .E(_09382_),
    .Y(_09383_));
 OA211x2_ASAP7_75t_R _27807_ (.A1(_01993_),
    .A2(_07145_),
    .B(_09383_),
    .C(_14688_),
    .Y(_09384_));
 OA211x2_ASAP7_75t_R _27808_ (.A1(_02137_),
    .A2(_07508_),
    .B(_07364_),
    .C(_09384_),
    .Y(_09385_));
 TAPCELL_ASAP7_75t_R TAP_612 ();
 NOR2x1_ASAP7_75t_R _27810_ (.A(_14502_),
    .B(_14688_),
    .Y(_09387_));
 AO21x1_ASAP7_75t_R _27811_ (.A1(_02289_),
    .A2(_14688_),
    .B(_09387_),
    .Y(_09388_));
 TAPCELL_ASAP7_75t_R TAP_611 ();
 AOI22x1_ASAP7_75t_R _27813_ (.A1(_07383_),
    .A2(_09385_),
    .B1(_09388_),
    .B2(net292),
    .Y(_09390_));
 INVx1_ASAP7_75t_R _27814_ (.A(_09390_),
    .Y(_09391_));
 TAPCELL_ASAP7_75t_R TAP_610 ();
 AOI22x1_ASAP7_75t_R _27816_ (.A1(_06880_),
    .A2(_09380_),
    .B1(_09391_),
    .B2(_09366_),
    .Y(_09393_));
 OA21x2_ASAP7_75t_R _27817_ (.A1(_07376_),
    .A2(_09367_),
    .B(_09393_),
    .Y(_02866_));
 AND2x2_ASAP7_75t_R _27818_ (.A(_14501_),
    .B(_14761_),
    .Y(_09394_));
 AO21x1_ASAP7_75t_R _27819_ (.A1(_02289_),
    .A2(_18121_),
    .B(_09394_),
    .Y(_09395_));
 NAND2x1_ASAP7_75t_R _27820_ (.A(_02286_),
    .B(_09395_),
    .Y(_09396_));
 OA21x2_ASAP7_75t_R _27821_ (.A1(_14761_),
    .A2(_07459_),
    .B(_09396_),
    .Y(_09397_));
 TAPCELL_ASAP7_75t_R TAP_609 ();
 AND2x2_ASAP7_75t_R _27823_ (.A(_00170_),
    .B(_09372_),
    .Y(_09399_));
 AO21x1_ASAP7_75t_R _27824_ (.A1(_01606_),
    .A2(_09370_),
    .B(_09399_),
    .Y(_09400_));
 OAI22x1_ASAP7_75t_R _27825_ (.A1(_00081_),
    .A2(_09367_),
    .B1(_09400_),
    .B2(_06873_),
    .Y(_09401_));
 AO21x1_ASAP7_75t_R _27826_ (.A1(_09355_),
    .A2(_09397_),
    .B(_09401_),
    .Y(_02867_));
 INVx1_ASAP7_75t_R _27827_ (.A(_00084_),
    .Y(_09402_));
 NOR2x2_ASAP7_75t_R _27828_ (.A(_06880_),
    .B(_09366_),
    .Y(_09403_));
 TAPCELL_ASAP7_75t_R TAP_608 ();
 NOR2x1_ASAP7_75t_R _27830_ (.A(_14502_),
    .B(_14822_),
    .Y(_09405_));
 AO21x1_ASAP7_75t_R _27831_ (.A1(_02289_),
    .A2(_14822_),
    .B(_09405_),
    .Y(_09406_));
 TAPCELL_ASAP7_75t_R TAP_607 ();
 AOI22x1_ASAP7_75t_R _27833_ (.A1(_14822_),
    .A2(_07530_),
    .B1(_09406_),
    .B2(net292),
    .Y(_09408_));
 TAPCELL_ASAP7_75t_R TAP_606 ();
 TAPCELL_ASAP7_75t_R TAP_605 ();
 AND2x2_ASAP7_75t_R _27836_ (.A(_00174_),
    .B(_09372_),
    .Y(_09411_));
 AO21x2_ASAP7_75t_R _27837_ (.A1(_01605_),
    .A2(_09370_),
    .B(_09411_),
    .Y(_09412_));
 NOR2x1_ASAP7_75t_R _27838_ (.A(_06873_),
    .B(_09412_),
    .Y(_09413_));
 AO221x1_ASAP7_75t_R _27839_ (.A1(_09402_),
    .A2(_09403_),
    .B1(_09408_),
    .B2(_09366_),
    .C(_09413_),
    .Y(_02868_));
 INVx1_ASAP7_75t_R _27840_ (.A(_00087_),
    .Y(_09414_));
 NOR2x1_ASAP7_75t_R _27841_ (.A(_14502_),
    .B(_18133_),
    .Y(_09415_));
 AO21x1_ASAP7_75t_R _27842_ (.A1(_02289_),
    .A2(_18133_),
    .B(_09415_),
    .Y(_09416_));
 AOI22x1_ASAP7_75t_R _27843_ (.A1(_18133_),
    .A2(_07578_),
    .B1(_09416_),
    .B2(net292),
    .Y(_09417_));
 TAPCELL_ASAP7_75t_R TAP_604 ();
 TAPCELL_ASAP7_75t_R TAP_603 ();
 AND2x2_ASAP7_75t_R _27846_ (.A(_00177_),
    .B(_09372_),
    .Y(_09420_));
 AO21x2_ASAP7_75t_R _27847_ (.A1(_01604_),
    .A2(_09370_),
    .B(_09420_),
    .Y(_09421_));
 NOR2x1_ASAP7_75t_R _27848_ (.A(_06873_),
    .B(_09421_),
    .Y(_09422_));
 AO221x1_ASAP7_75t_R _27849_ (.A1(_09414_),
    .A2(_09403_),
    .B1(_09417_),
    .B2(_09366_),
    .C(_09422_),
    .Y(_02869_));
 INVx1_ASAP7_75t_R _27850_ (.A(_00090_),
    .Y(_09423_));
 AND2x2_ASAP7_75t_R _27851_ (.A(_14501_),
    .B(_14938_),
    .Y(_09424_));
 AO21x1_ASAP7_75t_R _27852_ (.A1(net291),
    .A2(_18138_),
    .B(_09424_),
    .Y(_09425_));
 AOI22x1_ASAP7_75t_R _27853_ (.A1(_18138_),
    .A2(_07609_),
    .B1(_09425_),
    .B2(net293),
    .Y(_09426_));
 AND2x2_ASAP7_75t_R _27854_ (.A(_00180_),
    .B(_09372_),
    .Y(_09427_));
 AO21x1_ASAP7_75t_R _27855_ (.A1(_01603_),
    .A2(_09370_),
    .B(_09427_),
    .Y(_09428_));
 NOR2x1_ASAP7_75t_R _27856_ (.A(_06873_),
    .B(_09428_),
    .Y(_09429_));
 AO221x1_ASAP7_75t_R _27857_ (.A1(_09423_),
    .A2(_09403_),
    .B1(_09426_),
    .B2(_09366_),
    .C(_09429_),
    .Y(_02870_));
 NOR2x1_ASAP7_75t_R _27858_ (.A(_14502_),
    .B(_18143_),
    .Y(_09430_));
 AO21x1_ASAP7_75t_R _27859_ (.A1(_02289_),
    .A2(_18143_),
    .B(_09430_),
    .Y(_09431_));
 AOI22x1_ASAP7_75t_R _27860_ (.A1(_18143_),
    .A2(_07672_),
    .B1(_09431_),
    .B2(net292),
    .Y(_09432_));
 AND2x2_ASAP7_75t_R _27861_ (.A(_00182_),
    .B(_09372_),
    .Y(_09433_));
 AO21x2_ASAP7_75t_R _27862_ (.A1(_01602_),
    .A2(_09370_),
    .B(_09433_),
    .Y(_09434_));
 OAI22x1_ASAP7_75t_R _27863_ (.A1(_01574_),
    .A2(_09367_),
    .B1(_09434_),
    .B2(_06873_),
    .Y(_09435_));
 AO21x1_ASAP7_75t_R _27864_ (.A1(_09366_),
    .A2(_09432_),
    .B(_09435_),
    .Y(_02871_));
 NOR2x1_ASAP7_75t_R _27865_ (.A(_14502_),
    .B(_18148_),
    .Y(_09436_));
 AO21x1_ASAP7_75t_R _27866_ (.A1(_02289_),
    .A2(_18148_),
    .B(_09436_),
    .Y(_09437_));
 AOI22x1_ASAP7_75t_R _27867_ (.A1(_18148_),
    .A2(_07710_),
    .B1(_09437_),
    .B2(net292),
    .Y(_09438_));
 AND2x2_ASAP7_75t_R _27868_ (.A(_00186_),
    .B(_09372_),
    .Y(_09439_));
 AO21x1_ASAP7_75t_R _27869_ (.A1(_01601_),
    .A2(_09370_),
    .B(_09439_),
    .Y(_09440_));
 OAI22x1_ASAP7_75t_R _27870_ (.A1(_01573_),
    .A2(_09367_),
    .B1(_09440_),
    .B2(_06873_),
    .Y(_09441_));
 AO21x1_ASAP7_75t_R _27871_ (.A1(_09355_),
    .A2(_09438_),
    .B(_09441_),
    .Y(_02872_));
 INVx1_ASAP7_75t_R _27872_ (.A(_01572_),
    .Y(_09442_));
 AND2x2_ASAP7_75t_R _27873_ (.A(_14501_),
    .B(_15104_),
    .Y(_09443_));
 AO21x1_ASAP7_75t_R _27874_ (.A1(net291),
    .A2(_18153_),
    .B(_09443_),
    .Y(_09444_));
 AOI22x1_ASAP7_75t_R _27875_ (.A1(_18153_),
    .A2(_07777_),
    .B1(_09444_),
    .B2(net293),
    .Y(_09445_));
 AND2x2_ASAP7_75t_R _27876_ (.A(_00189_),
    .B(_09372_),
    .Y(_09446_));
 AO21x1_ASAP7_75t_R _27877_ (.A1(_01600_),
    .A2(_09370_),
    .B(_09446_),
    .Y(_09447_));
 NOR2x1_ASAP7_75t_R _27878_ (.A(_06873_),
    .B(_09447_),
    .Y(_09448_));
 AO221x1_ASAP7_75t_R _27879_ (.A1(_09442_),
    .A2(_09403_),
    .B1(_09445_),
    .B2(_09366_),
    .C(_09448_),
    .Y(_02873_));
 INVx1_ASAP7_75t_R _27880_ (.A(_01571_),
    .Y(_09449_));
 AND2x2_ASAP7_75t_R _27881_ (.A(_14501_),
    .B(_15159_),
    .Y(_09450_));
 AO21x1_ASAP7_75t_R _27882_ (.A1(net291),
    .A2(_18158_),
    .B(_09450_),
    .Y(_09451_));
 AOI22x1_ASAP7_75t_R _27883_ (.A1(_18158_),
    .A2(_07801_),
    .B1(_09451_),
    .B2(net293),
    .Y(_09452_));
 AND2x2_ASAP7_75t_R _27884_ (.A(_00193_),
    .B(_09372_),
    .Y(_09453_));
 AO21x1_ASAP7_75t_R _27885_ (.A1(_01599_),
    .A2(_09370_),
    .B(_09453_),
    .Y(_09454_));
 NOR2x1_ASAP7_75t_R _27886_ (.A(_06873_),
    .B(_09454_),
    .Y(_09455_));
 AO221x1_ASAP7_75t_R _27887_ (.A1(_09449_),
    .A2(_09403_),
    .B1(_09452_),
    .B2(_09366_),
    .C(_09455_),
    .Y(_02874_));
 NOR2x1_ASAP7_75t_R _27888_ (.A(_14502_),
    .B(_14576_),
    .Y(_09456_));
 AO21x1_ASAP7_75t_R _27889_ (.A1(_02289_),
    .A2(_14576_),
    .B(_09456_),
    .Y(_09457_));
 AOI22x1_ASAP7_75t_R _27890_ (.A1(_14576_),
    .A2(_07849_),
    .B1(_09457_),
    .B2(net292),
    .Y(_09458_));
 TAPCELL_ASAP7_75t_R TAP_602 ();
 AND2x2_ASAP7_75t_R _27892_ (.A(_00196_),
    .B(_09372_),
    .Y(_09460_));
 AO21x2_ASAP7_75t_R _27893_ (.A1(_01598_),
    .A2(_09370_),
    .B(_09460_),
    .Y(_09461_));
 OAI22x1_ASAP7_75t_R _27894_ (.A1(_01570_),
    .A2(_09367_),
    .B1(_09461_),
    .B2(_06873_),
    .Y(_09462_));
 AO21x1_ASAP7_75t_R _27895_ (.A1(_09366_),
    .A2(_09458_),
    .B(_09462_),
    .Y(_02875_));
 AND2x2_ASAP7_75t_R _27896_ (.A(_18165_),
    .B(_14501_),
    .Y(_09463_));
 AO21x1_ASAP7_75t_R _27897_ (.A1(_02289_),
    .A2(_18167_),
    .B(_09463_),
    .Y(_09464_));
 AOI22x1_ASAP7_75t_R _27898_ (.A1(_18167_),
    .A2(_07894_),
    .B1(_09464_),
    .B2(net292),
    .Y(_09465_));
 TAPCELL_ASAP7_75t_R TAP_601 ();
 AND2x2_ASAP7_75t_R _27900_ (.A(_00199_),
    .B(_09372_),
    .Y(_09467_));
 AO21x1_ASAP7_75t_R _27901_ (.A1(_01597_),
    .A2(_09370_),
    .B(_09467_),
    .Y(_09468_));
 OAI22x1_ASAP7_75t_R _27902_ (.A1(_01569_),
    .A2(_09367_),
    .B1(_09468_),
    .B2(_06873_),
    .Y(_09469_));
 AO21x1_ASAP7_75t_R _27903_ (.A1(_09366_),
    .A2(_09465_),
    .B(_09469_),
    .Y(_02876_));
 INVx1_ASAP7_75t_R _27904_ (.A(_01568_),
    .Y(_09470_));
 NOR2x1_ASAP7_75t_R _27905_ (.A(_14502_),
    .B(_15407_),
    .Y(_09471_));
 AO21x1_ASAP7_75t_R _27906_ (.A1(_02289_),
    .A2(_15407_),
    .B(_09471_),
    .Y(_09472_));
 AOI22x1_ASAP7_75t_R _27907_ (.A1(_15407_),
    .A2(_07932_),
    .B1(_09472_),
    .B2(net292),
    .Y(_09473_));
 TAPCELL_ASAP7_75t_R TAP_600 ();
 AND2x2_ASAP7_75t_R _27909_ (.A(_00201_),
    .B(_09372_),
    .Y(_09475_));
 AO21x2_ASAP7_75t_R _27910_ (.A1(_01596_),
    .A2(_09370_),
    .B(_09475_),
    .Y(_09476_));
 NOR2x1_ASAP7_75t_R _27911_ (.A(_06873_),
    .B(_09476_),
    .Y(_09477_));
 AO221x1_ASAP7_75t_R _27912_ (.A1(_09470_),
    .A2(_09403_),
    .B1(_09473_),
    .B2(_09366_),
    .C(_09477_),
    .Y(_02877_));
 INVx1_ASAP7_75t_R _27913_ (.A(_01567_),
    .Y(_09478_));
 NOR2x1_ASAP7_75t_R _27914_ (.A(_14502_),
    .B(_15556_),
    .Y(_09479_));
 AO21x1_ASAP7_75t_R _27915_ (.A1(_02289_),
    .A2(_15556_),
    .B(_09479_),
    .Y(_09480_));
 AOI22x1_ASAP7_75t_R _27916_ (.A1(_15556_),
    .A2(_07970_),
    .B1(_09480_),
    .B2(net292),
    .Y(_09481_));
 AND2x2_ASAP7_75t_R _27917_ (.A(_00204_),
    .B(_09372_),
    .Y(_09482_));
 AO21x2_ASAP7_75t_R _27918_ (.A1(_01595_),
    .A2(_09370_),
    .B(_09482_),
    .Y(_09483_));
 NOR2x1_ASAP7_75t_R _27919_ (.A(_06873_),
    .B(_09483_),
    .Y(_09484_));
 AO221x1_ASAP7_75t_R _27920_ (.A1(_09478_),
    .A2(_09403_),
    .B1(_09481_),
    .B2(_09366_),
    .C(_09484_),
    .Y(_02878_));
 INVx1_ASAP7_75t_R _27921_ (.A(_01566_),
    .Y(_09485_));
 AND2x2_ASAP7_75t_R _27922_ (.A(_14501_),
    .B(_15668_),
    .Y(_09486_));
 AO21x1_ASAP7_75t_R _27923_ (.A1(_02289_),
    .A2(_18182_),
    .B(_09486_),
    .Y(_09487_));
 AOI22x1_ASAP7_75t_R _27924_ (.A1(_18182_),
    .A2(_08017_),
    .B1(_09487_),
    .B2(_02286_),
    .Y(_09488_));
 TAPCELL_ASAP7_75t_R TAP_599 ();
 AND2x2_ASAP7_75t_R _27926_ (.A(_00206_),
    .B(_09372_),
    .Y(_09490_));
 AO21x2_ASAP7_75t_R _27927_ (.A1(_01594_),
    .A2(_09370_),
    .B(_09490_),
    .Y(_09491_));
 NOR2x1_ASAP7_75t_R _27928_ (.A(_06873_),
    .B(_09491_),
    .Y(_09492_));
 AO221x1_ASAP7_75t_R _27929_ (.A1(_09485_),
    .A2(_09403_),
    .B1(_09488_),
    .B2(_09366_),
    .C(_09492_),
    .Y(_02879_));
 NAND2x1_ASAP7_75t_R _27930_ (.A(_02289_),
    .B(_18186_),
    .Y(_09493_));
 OA21x2_ASAP7_75t_R _27931_ (.A1(_14502_),
    .A2(_18186_),
    .B(_09493_),
    .Y(_09494_));
 INVx1_ASAP7_75t_R _27932_ (.A(net293),
    .Y(_09495_));
 OA22x2_ASAP7_75t_R _27933_ (.A1(_15781_),
    .A2(_08068_),
    .B1(_09494_),
    .B2(_09495_),
    .Y(_09496_));
 TAPCELL_ASAP7_75t_R TAP_598 ();
 AND2x2_ASAP7_75t_R _27935_ (.A(_00208_),
    .B(_09372_),
    .Y(_09498_));
 AO21x1_ASAP7_75t_R _27936_ (.A1(_01593_),
    .A2(_09370_),
    .B(_09498_),
    .Y(_09499_));
 OAI22x1_ASAP7_75t_R _27937_ (.A1(_01565_),
    .A2(_09367_),
    .B1(_09499_),
    .B2(_06873_),
    .Y(_09500_));
 AO21x1_ASAP7_75t_R _27938_ (.A1(_09355_),
    .A2(_09496_),
    .B(_09500_),
    .Y(_02880_));
 NOR2x1_ASAP7_75t_R _27939_ (.A(_14502_),
    .B(_15897_),
    .Y(_09501_));
 AO21x1_ASAP7_75t_R _27940_ (.A1(_02289_),
    .A2(_15897_),
    .B(_09501_),
    .Y(_09502_));
 AOI22x1_ASAP7_75t_R _27941_ (.A1(_15897_),
    .A2(_08106_),
    .B1(_09502_),
    .B2(net292),
    .Y(_09503_));
 TAPCELL_ASAP7_75t_R TAP_597 ();
 AND2x2_ASAP7_75t_R _27943_ (.A(_00209_),
    .B(_09372_),
    .Y(_09505_));
 AO21x2_ASAP7_75t_R _27944_ (.A1(_01592_),
    .A2(_09370_),
    .B(_09505_),
    .Y(_09506_));
 TAPCELL_ASAP7_75t_R TAP_596 ();
 OAI22x1_ASAP7_75t_R _27946_ (.A1(_01564_),
    .A2(_09367_),
    .B1(_09506_),
    .B2(_06873_),
    .Y(_09508_));
 AO21x1_ASAP7_75t_R _27947_ (.A1(_09366_),
    .A2(_09503_),
    .B(_09508_),
    .Y(_02881_));
 AND2x2_ASAP7_75t_R _27948_ (.A(_14501_),
    .B(_18198_),
    .Y(_09509_));
 AO21x1_ASAP7_75t_R _27949_ (.A1(net291),
    .A2(_18196_),
    .B(_09509_),
    .Y(_09510_));
 AND2x2_ASAP7_75t_R _27950_ (.A(net293),
    .B(_09510_),
    .Y(_09511_));
 AOI21x1_ASAP7_75t_R _27951_ (.A1(_18196_),
    .A2(_08133_),
    .B(_09511_),
    .Y(_09512_));
 TAPCELL_ASAP7_75t_R TAP_595 ();
 AND2x2_ASAP7_75t_R _27953_ (.A(_00211_),
    .B(_09372_),
    .Y(_09514_));
 AO21x1_ASAP7_75t_R _27954_ (.A1(_01591_),
    .A2(_09370_),
    .B(_09514_),
    .Y(_09515_));
 OAI22x1_ASAP7_75t_R _27955_ (.A1(_01563_),
    .A2(_09367_),
    .B1(_09515_),
    .B2(_06873_),
    .Y(_09516_));
 AO21x1_ASAP7_75t_R _27956_ (.A1(_09355_),
    .A2(_09512_),
    .B(_09516_),
    .Y(_02882_));
 NOR2x1_ASAP7_75t_R _27957_ (.A(_14502_),
    .B(_16137_),
    .Y(_09517_));
 AO21x1_ASAP7_75t_R _27958_ (.A1(net291),
    .A2(_16137_),
    .B(_09517_),
    .Y(_09518_));
 AOI22x1_ASAP7_75t_R _27959_ (.A1(_16137_),
    .A2(_08178_),
    .B1(_09518_),
    .B2(net293),
    .Y(_09519_));
 TAPCELL_ASAP7_75t_R TAP_594 ();
 AND2x2_ASAP7_75t_R _27961_ (.A(_00212_),
    .B(_09372_),
    .Y(_09521_));
 AO21x1_ASAP7_75t_R _27962_ (.A1(_01590_),
    .A2(_09370_),
    .B(_09521_),
    .Y(_09522_));
 OAI22x1_ASAP7_75t_R _27963_ (.A1(_01562_),
    .A2(_09367_),
    .B1(_09522_),
    .B2(_06873_),
    .Y(_09523_));
 AO21x1_ASAP7_75t_R _27964_ (.A1(_09355_),
    .A2(_09519_),
    .B(_09523_),
    .Y(_02883_));
 AND2x2_ASAP7_75t_R _27965_ (.A(_14501_),
    .B(_16259_),
    .Y(_09524_));
 AO21x1_ASAP7_75t_R _27966_ (.A1(net291),
    .A2(_18206_),
    .B(_09524_),
    .Y(_09525_));
 AOI22x1_ASAP7_75t_R _27967_ (.A1(_18206_),
    .A2(_08215_),
    .B1(_09525_),
    .B2(net293),
    .Y(_09526_));
 AND2x2_ASAP7_75t_R _27968_ (.A(_00214_),
    .B(_09372_),
    .Y(_09527_));
 AO21x1_ASAP7_75t_R _27969_ (.A1(_01589_),
    .A2(_09370_),
    .B(_09527_),
    .Y(_09528_));
 OAI22x1_ASAP7_75t_R _27970_ (.A1(_01561_),
    .A2(_09367_),
    .B1(_09528_),
    .B2(_06873_),
    .Y(_09529_));
 AO21x1_ASAP7_75t_R _27971_ (.A1(_09366_),
    .A2(_09526_),
    .B(_09529_),
    .Y(_02884_));
 NOR2x1_ASAP7_75t_R _27972_ (.A(_14502_),
    .B(_18211_),
    .Y(_09530_));
 AO21x1_ASAP7_75t_R _27973_ (.A1(_02289_),
    .A2(_18211_),
    .B(_09530_),
    .Y(_09531_));
 AOI22x1_ASAP7_75t_R _27974_ (.A1(_18211_),
    .A2(_08244_),
    .B1(_09531_),
    .B2(net292),
    .Y(_09532_));
 TAPCELL_ASAP7_75t_R TAP_593 ();
 AND2x2_ASAP7_75t_R _27976_ (.A(_00215_),
    .B(_09372_),
    .Y(_09534_));
 AO21x1_ASAP7_75t_R _27977_ (.A1(_01588_),
    .A2(_09370_),
    .B(_09534_),
    .Y(_09535_));
 OAI22x1_ASAP7_75t_R _27978_ (.A1(_01560_),
    .A2(_09367_),
    .B1(_09535_),
    .B2(_06873_),
    .Y(_09536_));
 AO21x1_ASAP7_75t_R _27979_ (.A1(_09366_),
    .A2(_09532_),
    .B(_09536_),
    .Y(_02885_));
 NOR2x1_ASAP7_75t_R _27980_ (.A(_14502_),
    .B(_16480_),
    .Y(_09537_));
 AO21x1_ASAP7_75t_R _27981_ (.A1(_02289_),
    .A2(_16480_),
    .B(_09537_),
    .Y(_09538_));
 AOI22x1_ASAP7_75t_R _27982_ (.A1(_16480_),
    .A2(_08273_),
    .B1(_09538_),
    .B2(net292),
    .Y(_09539_));
 AND2x2_ASAP7_75t_R _27983_ (.A(_00217_),
    .B(_09372_),
    .Y(_09540_));
 AO21x1_ASAP7_75t_R _27984_ (.A1(_01587_),
    .A2(_09370_),
    .B(_09540_),
    .Y(_09541_));
 OAI22x1_ASAP7_75t_R _27985_ (.A1(_01559_),
    .A2(_09367_),
    .B1(_09541_),
    .B2(_06873_),
    .Y(_09542_));
 AO21x1_ASAP7_75t_R _27986_ (.A1(_09355_),
    .A2(_09539_),
    .B(_09542_),
    .Y(_02886_));
 AND2x2_ASAP7_75t_R _27987_ (.A(_14501_),
    .B(_04603_),
    .Y(_09543_));
 AO21x1_ASAP7_75t_R _27988_ (.A1(net291),
    .A2(_18222_),
    .B(_09543_),
    .Y(_09544_));
 AOI22x1_ASAP7_75t_R _27989_ (.A1(_18222_),
    .A2(_08315_),
    .B1(_09544_),
    .B2(net293),
    .Y(_09545_));
 TAPCELL_ASAP7_75t_R TAP_592 ();
 AND2x2_ASAP7_75t_R _27991_ (.A(_00218_),
    .B(_09372_),
    .Y(_09547_));
 AO21x1_ASAP7_75t_R _27992_ (.A1(_01586_),
    .A2(_09370_),
    .B(_09547_),
    .Y(_09548_));
 OAI22x1_ASAP7_75t_R _27993_ (.A1(_01558_),
    .A2(_09367_),
    .B1(_09548_),
    .B2(_06873_),
    .Y(_09549_));
 AO21x1_ASAP7_75t_R _27994_ (.A1(_09355_),
    .A2(_09545_),
    .B(_09549_),
    .Y(_02887_));
 AND2x2_ASAP7_75t_R _27995_ (.A(_00220_),
    .B(_09372_),
    .Y(_09550_));
 AO21x1_ASAP7_75t_R _27996_ (.A1(_01585_),
    .A2(_09370_),
    .B(_09550_),
    .Y(_09551_));
 AND2x2_ASAP7_75t_R _27997_ (.A(_14501_),
    .B(_04718_),
    .Y(_09552_));
 AO21x1_ASAP7_75t_R _27998_ (.A1(_02289_),
    .A2(_18226_),
    .B(_09552_),
    .Y(_09553_));
 INVx1_ASAP7_75t_R _27999_ (.A(_08347_),
    .Y(_09554_));
 OAI22x1_ASAP7_75t_R _28000_ (.A1(_01955_),
    .A2(_07659_),
    .B1(_07150_),
    .B2(_00141_),
    .Y(_09555_));
 AO221x1_ASAP7_75t_R _28001_ (.A1(_05538_),
    .A2(_05584_),
    .B1(_07155_),
    .B2(net78),
    .C(_04718_),
    .Y(_09556_));
 AO21x1_ASAP7_75t_R _28002_ (.A1(_05632_),
    .A2(_09555_),
    .B(_09556_),
    .Y(_09557_));
 AOI21x1_ASAP7_75t_R _28003_ (.A1(_06884_),
    .A2(_08348_),
    .B(_09557_),
    .Y(_09558_));
 OA211x2_ASAP7_75t_R _28004_ (.A1(_08338_),
    .A2(_08341_),
    .B(_09554_),
    .C(_09558_),
    .Y(_09559_));
 AO21x2_ASAP7_75t_R _28005_ (.A1(net292),
    .A2(_09553_),
    .B(_09559_),
    .Y(_09560_));
 INVx1_ASAP7_75t_R _28006_ (.A(_09366_),
    .Y(_09561_));
 OA22x2_ASAP7_75t_R _28007_ (.A1(_06873_),
    .A2(_09551_),
    .B1(_09560_),
    .B2(_09561_),
    .Y(_09562_));
 OAI21x1_ASAP7_75t_R _28008_ (.A1(_01557_),
    .A2(_09367_),
    .B(_09562_),
    .Y(_02888_));
 AND2x2_ASAP7_75t_R _28009_ (.A(_14501_),
    .B(_04829_),
    .Y(_09563_));
 AO21x1_ASAP7_75t_R _28010_ (.A1(net291),
    .A2(_18231_),
    .B(_09563_),
    .Y(_09564_));
 AOI22x1_ASAP7_75t_R _28011_ (.A1(_18231_),
    .A2(_08385_),
    .B1(_09564_),
    .B2(net293),
    .Y(_09565_));
 TAPCELL_ASAP7_75t_R TAP_591 ();
 AND2x2_ASAP7_75t_R _28013_ (.A(_00221_),
    .B(_09372_),
    .Y(_09567_));
 AO21x1_ASAP7_75t_R _28014_ (.A1(_01584_),
    .A2(_09370_),
    .B(_09567_),
    .Y(_09568_));
 OAI22x1_ASAP7_75t_R _28015_ (.A1(_01556_),
    .A2(_09367_),
    .B1(_09568_),
    .B2(_06873_),
    .Y(_09569_));
 AO21x1_ASAP7_75t_R _28016_ (.A1(_09355_),
    .A2(_09565_),
    .B(_09569_),
    .Y(_02889_));
 AND2x2_ASAP7_75t_R _28017_ (.A(_14501_),
    .B(_18235_),
    .Y(_09570_));
 AO21x1_ASAP7_75t_R _28018_ (.A1(net291),
    .A2(_18237_),
    .B(_09570_),
    .Y(_09571_));
 AOI22x1_ASAP7_75t_R _28019_ (.A1(_18237_),
    .A2(_08412_),
    .B1(_09571_),
    .B2(net293),
    .Y(_09572_));
 AND2x2_ASAP7_75t_R _28020_ (.A(_00223_),
    .B(_09372_),
    .Y(_09573_));
 AO21x1_ASAP7_75t_R _28021_ (.A1(_01583_),
    .A2(_09370_),
    .B(_09573_),
    .Y(_09574_));
 OAI22x1_ASAP7_75t_R _28022_ (.A1(_01555_),
    .A2(_09367_),
    .B1(_09574_),
    .B2(_06873_),
    .Y(_09575_));
 AO21x1_ASAP7_75t_R _28023_ (.A1(_09355_),
    .A2(_09572_),
    .B(_09575_),
    .Y(_02890_));
 AND2x2_ASAP7_75t_R _28024_ (.A(_14501_),
    .B(_05045_),
    .Y(_09576_));
 AO21x1_ASAP7_75t_R _28025_ (.A1(net291),
    .A2(_18242_),
    .B(_09576_),
    .Y(_09577_));
 AOI22x1_ASAP7_75t_R _28026_ (.A1(_18242_),
    .A2(_08445_),
    .B1(_09577_),
    .B2(net293),
    .Y(_09578_));
 TAPCELL_ASAP7_75t_R TAP_590 ();
 AND2x2_ASAP7_75t_R _28028_ (.A(_00224_),
    .B(_09372_),
    .Y(_09580_));
 AO21x1_ASAP7_75t_R _28029_ (.A1(_01582_),
    .A2(_09370_),
    .B(_09580_),
    .Y(_09581_));
 OAI22x1_ASAP7_75t_R _28030_ (.A1(_01554_),
    .A2(_09367_),
    .B1(_09581_),
    .B2(_06873_),
    .Y(_09582_));
 AO21x1_ASAP7_75t_R _28031_ (.A1(_09355_),
    .A2(_09578_),
    .B(_09582_),
    .Y(_02891_));
 AND2x2_ASAP7_75t_R _28032_ (.A(net291),
    .B(_18246_),
    .Y(_09583_));
 AO21x1_ASAP7_75t_R _28033_ (.A1(_14501_),
    .A2(_18248_),
    .B(_09583_),
    .Y(_09584_));
 AOI22x1_ASAP7_75t_R _28034_ (.A1(_18246_),
    .A2(_08478_),
    .B1(_09584_),
    .B2(net293),
    .Y(_09585_));
 AND2x2_ASAP7_75t_R _28035_ (.A(_00226_),
    .B(_09372_),
    .Y(_09586_));
 AO21x1_ASAP7_75t_R _28036_ (.A1(_01581_),
    .A2(_09370_),
    .B(_09586_),
    .Y(_09587_));
 OAI22x1_ASAP7_75t_R _28037_ (.A1(_01553_),
    .A2(_09367_),
    .B1(_09587_),
    .B2(_06873_),
    .Y(_09588_));
 AO21x1_ASAP7_75t_R _28038_ (.A1(_09355_),
    .A2(_09585_),
    .B(_09588_),
    .Y(_02892_));
 NAND2x1_ASAP7_75t_R _28039_ (.A(net291),
    .B(_18251_),
    .Y(_09589_));
 OA21x2_ASAP7_75t_R _28040_ (.A1(_14502_),
    .A2(_18251_),
    .B(_09589_),
    .Y(_09590_));
 OA22x2_ASAP7_75t_R _28041_ (.A1(_18253_),
    .A2(_08509_),
    .B1(_09590_),
    .B2(_09495_),
    .Y(_09591_));
 TAPCELL_ASAP7_75t_R TAP_589 ();
 AND2x2_ASAP7_75t_R _28043_ (.A(_00227_),
    .B(_09372_),
    .Y(_09593_));
 AO21x2_ASAP7_75t_R _28044_ (.A1(_01580_),
    .A2(_09370_),
    .B(_09593_),
    .Y(_09594_));
 OAI22x1_ASAP7_75t_R _28045_ (.A1(_01552_),
    .A2(_09367_),
    .B1(_09594_),
    .B2(_06873_),
    .Y(_09595_));
 AO21x1_ASAP7_75t_R _28046_ (.A1(_09355_),
    .A2(_09591_),
    .B(_09595_),
    .Y(_02893_));
 AND2x2_ASAP7_75t_R _28047_ (.A(_14501_),
    .B(_05371_),
    .Y(_09596_));
 AO21x1_ASAP7_75t_R _28048_ (.A1(net291),
    .A2(_18256_),
    .B(_09596_),
    .Y(_09597_));
 AOI22x1_ASAP7_75t_R _28049_ (.A1(_18256_),
    .A2(_08542_),
    .B1(_09597_),
    .B2(net293),
    .Y(_09598_));
 AND2x2_ASAP7_75t_R _28050_ (.A(_00229_),
    .B(_09372_),
    .Y(_09599_));
 AO21x1_ASAP7_75t_R _28051_ (.A1(_01579_),
    .A2(_09370_),
    .B(_09599_),
    .Y(_09600_));
 OAI22x1_ASAP7_75t_R _28052_ (.A1(_01551_),
    .A2(_09367_),
    .B1(_09600_),
    .B2(_06873_),
    .Y(_09601_));
 AO21x1_ASAP7_75t_R _28053_ (.A1(_09366_),
    .A2(_09598_),
    .B(_09601_),
    .Y(_02894_));
 INVx1_ASAP7_75t_R _28054_ (.A(_01550_),
    .Y(_09602_));
 AND2x2_ASAP7_75t_R _28055_ (.A(_14501_),
    .B(_05478_),
    .Y(_09603_));
 AO21x1_ASAP7_75t_R _28056_ (.A1(_02289_),
    .A2(_17587_),
    .B(_09603_),
    .Y(_09604_));
 AOI22x1_ASAP7_75t_R _28057_ (.A1(_17587_),
    .A2(_08568_),
    .B1(_09604_),
    .B2(_02286_),
    .Y(_09605_));
 AND2x2_ASAP7_75t_R _28058_ (.A(_00230_),
    .B(_09372_),
    .Y(_09606_));
 AO21x1_ASAP7_75t_R _28059_ (.A1(_01578_),
    .A2(_09370_),
    .B(_09606_),
    .Y(_09607_));
 NOR2x1_ASAP7_75t_R _28060_ (.A(_06873_),
    .B(_09607_),
    .Y(_09608_));
 AO221x1_ASAP7_75t_R _28061_ (.A1(_09602_),
    .A2(_09403_),
    .B1(_09605_),
    .B2(_09366_),
    .C(_09608_),
    .Y(_02895_));
 NAND2x2_ASAP7_75t_R _28062_ (.A(net286),
    .B(_06771_),
    .Y(_09609_));
 TAPCELL_ASAP7_75t_R TAP_588 ();
 AND3x1_ASAP7_75t_R _28064_ (.A(_01549_),
    .B(net287),
    .C(_06771_),
    .Y(_09611_));
 AOI21x1_ASAP7_75t_R _28065_ (.A1(_02596_),
    .A2(_09609_),
    .B(_09611_),
    .Y(_02896_));
 AND3x1_ASAP7_75t_R _28066_ (.A(_01548_),
    .B(net287),
    .C(_06771_),
    .Y(_09612_));
 AOI21x1_ASAP7_75t_R _28067_ (.A1(_02567_),
    .A2(_09609_),
    .B(_09612_),
    .Y(_02897_));
 AND3x1_ASAP7_75t_R _28068_ (.A(_01547_),
    .B(net287),
    .C(_06771_),
    .Y(_09613_));
 AOI21x1_ASAP7_75t_R _28069_ (.A1(_02569_),
    .A2(_09609_),
    .B(_09613_),
    .Y(_02898_));
 TAPCELL_ASAP7_75t_R TAP_587 ();
 XOR2x1_ASAP7_75t_R _28071_ (.A(_02568_),
    .Y(_09615_),
    .B(_06311_));
 TAPCELL_ASAP7_75t_R TAP_586 ();
 NOR2x1_ASAP7_75t_R _28073_ (.A(_01546_),
    .B(_09609_),
    .Y(_09617_));
 AO21x1_ASAP7_75t_R _28074_ (.A1(_09609_),
    .A2(_09615_),
    .B(_09617_),
    .Y(_02899_));
 AND3x1_ASAP7_75t_R _28075_ (.A(_01545_),
    .B(net287),
    .C(_06771_),
    .Y(_09618_));
 AOI21x1_ASAP7_75t_R _28076_ (.A1(_02571_),
    .A2(_09609_),
    .B(_09618_),
    .Y(_02900_));
 XOR2x1_ASAP7_75t_R _28077_ (.A(_02570_),
    .Y(_09619_),
    .B(_06334_));
 NOR2x1_ASAP7_75t_R _28078_ (.A(_01544_),
    .B(_09609_),
    .Y(_09620_));
 AO21x1_ASAP7_75t_R _28079_ (.A1(_09609_),
    .A2(_09619_),
    .B(_09620_),
    .Y(_02901_));
 NAND2x1_ASAP7_75t_R _28080_ (.A(_02573_),
    .B(_09609_),
    .Y(_09621_));
 OA21x2_ASAP7_75t_R _28081_ (.A1(_06336_),
    .A2(_09609_),
    .B(_09621_),
    .Y(_02902_));
 OR3x1_ASAP7_75t_R _28082_ (.A(_06312_),
    .B(_02572_),
    .C(_06516_),
    .Y(_09622_));
 XOR2x1_ASAP7_75t_R _28083_ (.A(_01542_),
    .Y(_09623_),
    .B(_09622_));
 XOR2x1_ASAP7_75t_R _28084_ (.A(_02572_),
    .Y(_09624_),
    .B(_06354_));
 AND2x2_ASAP7_75t_R _28085_ (.A(_06254_),
    .B(_09624_),
    .Y(_09625_));
 AO21x1_ASAP7_75t_R _28086_ (.A1(net287),
    .A2(_09623_),
    .B(_09625_),
    .Y(_02903_));
 AND3x1_ASAP7_75t_R _28087_ (.A(_01541_),
    .B(net287),
    .C(_06771_),
    .Y(_09626_));
 AOI21x1_ASAP7_75t_R _28088_ (.A1(_02575_),
    .A2(_09609_),
    .B(_09626_),
    .Y(_02904_));
 AND2x6_ASAP7_75t_R _28089_ (.A(net286),
    .B(_06771_),
    .Y(_09627_));
 XOR2x1_ASAP7_75t_R _28090_ (.A(_02574_),
    .Y(_09628_),
    .B(_06376_));
 NAND2x1_ASAP7_75t_R _28091_ (.A(_01540_),
    .B(_09627_),
    .Y(_09629_));
 OA21x2_ASAP7_75t_R _28092_ (.A1(_09627_),
    .A2(_09628_),
    .B(_09629_),
    .Y(_02905_));
 AND3x1_ASAP7_75t_R _28093_ (.A(_01539_),
    .B(net287),
    .C(_06771_),
    .Y(_09630_));
 AOI21x1_ASAP7_75t_R _28094_ (.A1(_02577_),
    .A2(_09609_),
    .B(_09630_),
    .Y(_02906_));
 OR3x1_ASAP7_75t_R _28095_ (.A(_06312_),
    .B(_02576_),
    .C(_06516_),
    .Y(_09631_));
 XOR2x1_ASAP7_75t_R _28096_ (.A(_01538_),
    .Y(_09632_),
    .B(_09631_));
 XOR2x1_ASAP7_75t_R _28097_ (.A(_02576_),
    .Y(_09633_),
    .B(_06388_));
 AND2x2_ASAP7_75t_R _28098_ (.A(_06254_),
    .B(_09633_),
    .Y(_09634_));
 AO21x1_ASAP7_75t_R _28099_ (.A1(net287),
    .A2(_09632_),
    .B(_09634_),
    .Y(_02907_));
 AND3x1_ASAP7_75t_R _28100_ (.A(_01537_),
    .B(net287),
    .C(_06771_),
    .Y(_09635_));
 AOI21x1_ASAP7_75t_R _28101_ (.A1(_02579_),
    .A2(_09609_),
    .B(_09635_),
    .Y(_02908_));
 XOR2x1_ASAP7_75t_R _28102_ (.A(_02578_),
    .Y(_09636_),
    .B(_06401_));
 NOR2x1_ASAP7_75t_R _28103_ (.A(_01536_),
    .B(_09609_),
    .Y(_09637_));
 AO21x1_ASAP7_75t_R _28104_ (.A1(_09609_),
    .A2(_09636_),
    .B(_09637_),
    .Y(_02909_));
 AND3x1_ASAP7_75t_R _28105_ (.A(_01535_),
    .B(net286),
    .C(_06771_),
    .Y(_09638_));
 AOI21x1_ASAP7_75t_R _28106_ (.A1(_02581_),
    .A2(_09609_),
    .B(_09638_),
    .Y(_02910_));
 XOR2x1_ASAP7_75t_R _28107_ (.A(_02580_),
    .Y(_09639_),
    .B(_06416_));
 NOR2x1_ASAP7_75t_R _28108_ (.A(_01534_),
    .B(_09609_),
    .Y(_09640_));
 AO21x1_ASAP7_75t_R _28109_ (.A1(_09609_),
    .A2(_09639_),
    .B(_09640_),
    .Y(_02911_));
 AND3x1_ASAP7_75t_R _28110_ (.A(_01533_),
    .B(net286),
    .C(_06771_),
    .Y(_09641_));
 AOI21x1_ASAP7_75t_R _28111_ (.A1(_02583_),
    .A2(_09609_),
    .B(_09641_),
    .Y(_02912_));
 XNOR2x1_ASAP7_75t_R _28112_ (.B(_06430_),
    .Y(_09642_),
    .A(_02582_));
 NOR2x1_ASAP7_75t_R _28113_ (.A(_01532_),
    .B(_09609_),
    .Y(_09643_));
 AO21x1_ASAP7_75t_R _28114_ (.A1(_09609_),
    .A2(_09642_),
    .B(_09643_),
    .Y(_02913_));
 AND3x1_ASAP7_75t_R _28115_ (.A(_01531_),
    .B(net286),
    .C(_06771_),
    .Y(_09644_));
 AOI21x1_ASAP7_75t_R _28116_ (.A1(_02585_),
    .A2(_09609_),
    .B(_09644_),
    .Y(_02914_));
 XNOR2x1_ASAP7_75t_R _28117_ (.B(_06444_),
    .Y(_09645_),
    .A(_02584_));
 NOR2x1_ASAP7_75t_R _28118_ (.A(_01530_),
    .B(_09609_),
    .Y(_09646_));
 AO21x1_ASAP7_75t_R _28119_ (.A1(_09609_),
    .A2(_09645_),
    .B(_09646_),
    .Y(_02915_));
 AND3x1_ASAP7_75t_R _28120_ (.A(_01529_),
    .B(net286),
    .C(_06771_),
    .Y(_09647_));
 AOI21x1_ASAP7_75t_R _28121_ (.A1(_02587_),
    .A2(_09609_),
    .B(_09647_),
    .Y(_02916_));
 XNOR2x1_ASAP7_75t_R _28122_ (.B(_06456_),
    .Y(_09648_),
    .A(_02586_));
 NAND2x1_ASAP7_75t_R _28123_ (.A(_01528_),
    .B(_09627_),
    .Y(_09649_));
 OA21x2_ASAP7_75t_R _28124_ (.A1(_09627_),
    .A2(_09648_),
    .B(_09649_),
    .Y(_02917_));
 AND3x1_ASAP7_75t_R _28125_ (.A(_01527_),
    .B(net286),
    .C(_06771_),
    .Y(_09650_));
 AOI21x1_ASAP7_75t_R _28126_ (.A1(_02589_),
    .A2(_09609_),
    .B(_09650_),
    .Y(_02918_));
 XNOR2x1_ASAP7_75t_R _28127_ (.B(_06469_),
    .Y(_09651_),
    .A(_02588_));
 NAND2x1_ASAP7_75t_R _28128_ (.A(_01526_),
    .B(_09627_),
    .Y(_09652_));
 OA21x2_ASAP7_75t_R _28129_ (.A1(_09627_),
    .A2(_09651_),
    .B(_09652_),
    .Y(_02919_));
 AND3x1_ASAP7_75t_R _28130_ (.A(_01525_),
    .B(net286),
    .C(_06771_),
    .Y(_09653_));
 AOI21x1_ASAP7_75t_R _28131_ (.A1(_02591_),
    .A2(_09609_),
    .B(_09653_),
    .Y(_02920_));
 XNOR2x1_ASAP7_75t_R _28132_ (.B(_06482_),
    .Y(_09654_),
    .A(_02590_));
 NAND2x1_ASAP7_75t_R _28133_ (.A(_01524_),
    .B(_09627_),
    .Y(_09655_));
 OA21x2_ASAP7_75t_R _28134_ (.A1(_09627_),
    .A2(_09654_),
    .B(_09655_),
    .Y(_02921_));
 AND3x1_ASAP7_75t_R _28135_ (.A(_01523_),
    .B(net286),
    .C(_06771_),
    .Y(_09656_));
 AOI21x1_ASAP7_75t_R _28136_ (.A1(_02593_),
    .A2(_09609_),
    .B(_09656_),
    .Y(_02922_));
 XNOR2x1_ASAP7_75t_R _28137_ (.B(_06495_),
    .Y(_09657_),
    .A(_02592_));
 NAND2x1_ASAP7_75t_R _28138_ (.A(_01522_),
    .B(_09627_),
    .Y(_09658_));
 OA21x2_ASAP7_75t_R _28139_ (.A1(_09627_),
    .A2(_09657_),
    .B(_09658_),
    .Y(_02923_));
 AND3x1_ASAP7_75t_R _28140_ (.A(_01521_),
    .B(net286),
    .C(_06771_),
    .Y(_09659_));
 AOI21x1_ASAP7_75t_R _28141_ (.A1(_02595_),
    .A2(_09609_),
    .B(_09659_),
    .Y(_02924_));
 XOR2x1_ASAP7_75t_R _28142_ (.A(_02594_),
    .Y(_09660_),
    .B(_06506_));
 NOR2x1_ASAP7_75t_R _28143_ (.A(_01520_),
    .B(_09609_),
    .Y(_09661_));
 AO21x1_ASAP7_75t_R _28144_ (.A1(_09609_),
    .A2(_09660_),
    .B(_09661_),
    .Y(_02925_));
 TAPCELL_ASAP7_75t_R TAP_585 ();
 AND2x2_ASAP7_75t_R _28146_ (.A(_00323_),
    .B(_05548_),
    .Y(_09663_));
 AND3x2_ASAP7_75t_R _28147_ (.A(_00194_),
    .B(_06922_),
    .C(_09663_),
    .Y(_09664_));
 AND2x6_ASAP7_75t_R _28148_ (.A(_06881_),
    .B(_09664_),
    .Y(_09665_));
 TAPCELL_ASAP7_75t_R TAP_584 ();
 TAPCELL_ASAP7_75t_R TAP_583 ();
 TAPCELL_ASAP7_75t_R TAP_582 ();
 NOR2x1_ASAP7_75t_R _28152_ (.A(_00293_),
    .B(_09665_),
    .Y(_09669_));
 AO21x1_ASAP7_75t_R _28153_ (.A1(_07180_),
    .A2(_09665_),
    .B(_09669_),
    .Y(_02926_));
 TAPCELL_ASAP7_75t_R TAP_581 ();
 NOR2x1_ASAP7_75t_R _28155_ (.A(_00247_),
    .B(_09665_),
    .Y(_09671_));
 AO21x1_ASAP7_75t_R _28156_ (.A1(_07313_),
    .A2(_09665_),
    .B(_09671_),
    .Y(_02927_));
 TAPCELL_ASAP7_75t_R TAP_580 ();
 NOR2x1_ASAP7_75t_R _28158_ (.A(_00355_),
    .B(_09665_),
    .Y(_09673_));
 AO21x1_ASAP7_75t_R _28159_ (.A1(_07398_),
    .A2(_09665_),
    .B(_09673_),
    .Y(_02928_));
 TAPCELL_ASAP7_75t_R TAP_579 ();
 NOR2x1_ASAP7_75t_R _28161_ (.A(_00386_),
    .B(_09665_),
    .Y(_09675_));
 AO21x1_ASAP7_75t_R _28162_ (.A1(_07469_),
    .A2(_09665_),
    .B(_09675_),
    .Y(_02929_));
 TAPCELL_ASAP7_75t_R TAP_578 ();
 NOR2x1_ASAP7_75t_R _28164_ (.A(_00416_),
    .B(_09665_),
    .Y(_09677_));
 AO21x1_ASAP7_75t_R _28165_ (.A1(_07534_),
    .A2(_09665_),
    .B(_09677_),
    .Y(_02930_));
 TAPCELL_ASAP7_75t_R TAP_577 ();
 NOR2x1_ASAP7_75t_R _28167_ (.A(_00446_),
    .B(_09665_),
    .Y(_09679_));
 AO21x1_ASAP7_75t_R _28168_ (.A1(_07581_),
    .A2(_09665_),
    .B(_09679_),
    .Y(_02931_));
 TAPCELL_ASAP7_75t_R TAP_576 ();
 NOR2x1_ASAP7_75t_R _28170_ (.A(_00476_),
    .B(_09665_),
    .Y(_09681_));
 AO21x1_ASAP7_75t_R _28171_ (.A1(net253),
    .A2(_09665_),
    .B(_09681_),
    .Y(_02932_));
 TAPCELL_ASAP7_75t_R TAP_575 ();
 NOR2x1_ASAP7_75t_R _28173_ (.A(_00506_),
    .B(_09665_),
    .Y(_09683_));
 AO21x1_ASAP7_75t_R _28174_ (.A1(_07676_),
    .A2(_09665_),
    .B(_09683_),
    .Y(_02933_));
 TAPCELL_ASAP7_75t_R TAP_574 ();
 TAPCELL_ASAP7_75t_R TAP_573 ();
 NOR2x1_ASAP7_75t_R _28177_ (.A(_00536_),
    .B(_09665_),
    .Y(_09686_));
 AO21x1_ASAP7_75t_R _28178_ (.A1(_07738_),
    .A2(_09665_),
    .B(_09686_),
    .Y(_02934_));
 TAPCELL_ASAP7_75t_R TAP_572 ();
 NOR2x1_ASAP7_75t_R _28180_ (.A(_00566_),
    .B(_09665_),
    .Y(_09688_));
 AO21x1_ASAP7_75t_R _28181_ (.A1(_07780_),
    .A2(_09665_),
    .B(_09688_),
    .Y(_02935_));
 TAPCELL_ASAP7_75t_R TAP_571 ();
 TAPCELL_ASAP7_75t_R TAP_570 ();
 NOR2x1_ASAP7_75t_R _28184_ (.A(_00596_),
    .B(_09665_),
    .Y(_09691_));
 AO21x1_ASAP7_75t_R _28185_ (.A1(_07817_),
    .A2(_09665_),
    .B(_09691_),
    .Y(_02936_));
 TAPCELL_ASAP7_75t_R TAP_569 ();
 NOR2x1_ASAP7_75t_R _28187_ (.A(_00626_),
    .B(_09665_),
    .Y(_09693_));
 AO21x1_ASAP7_75t_R _28188_ (.A1(_07865_),
    .A2(_09665_),
    .B(_09693_),
    .Y(_02937_));
 TAPCELL_ASAP7_75t_R TAP_568 ();
 NOR2x1_ASAP7_75t_R _28190_ (.A(_00325_),
    .B(_09665_),
    .Y(_09695_));
 AO21x1_ASAP7_75t_R _28191_ (.A1(_07908_),
    .A2(_09665_),
    .B(_09695_),
    .Y(_02938_));
 TAPCELL_ASAP7_75t_R TAP_567 ();
 NOR2x1_ASAP7_75t_R _28193_ (.A(_00688_),
    .B(_09665_),
    .Y(_09697_));
 AO21x1_ASAP7_75t_R _28194_ (.A1(_07950_),
    .A2(_09665_),
    .B(_09697_),
    .Y(_02939_));
 TAPCELL_ASAP7_75t_R TAP_566 ();
 NOR2x1_ASAP7_75t_R _28196_ (.A(_00720_),
    .B(_09665_),
    .Y(_09699_));
 AO21x1_ASAP7_75t_R _28197_ (.A1(_07990_),
    .A2(_09665_),
    .B(_09699_),
    .Y(_02940_));
 TAPCELL_ASAP7_75t_R TAP_565 ();
 NOR2x1_ASAP7_75t_R _28199_ (.A(_00753_),
    .B(_09665_),
    .Y(_09701_));
 AO21x1_ASAP7_75t_R _28200_ (.A1(_08034_),
    .A2(_09665_),
    .B(_09701_),
    .Y(_02941_));
 TAPCELL_ASAP7_75t_R TAP_564 ();
 NOR2x1_ASAP7_75t_R _28202_ (.A(_00786_),
    .B(_09665_),
    .Y(_09703_));
 AO21x1_ASAP7_75t_R _28203_ (.A1(_08073_),
    .A2(_09665_),
    .B(_09703_),
    .Y(_02942_));
 TAPCELL_ASAP7_75t_R TAP_563 ();
 NOR2x1_ASAP7_75t_R _28205_ (.A(_00819_),
    .B(_09665_),
    .Y(_09705_));
 AO21x1_ASAP7_75t_R _28206_ (.A1(_08116_),
    .A2(_09665_),
    .B(_09705_),
    .Y(_02943_));
 TAPCELL_ASAP7_75t_R TAP_562 ();
 TAPCELL_ASAP7_75t_R TAP_561 ();
 NOR2x1_ASAP7_75t_R _28209_ (.A(_00851_),
    .B(_09665_),
    .Y(_09708_));
 AO21x1_ASAP7_75t_R _28210_ (.A1(_08150_),
    .A2(_09665_),
    .B(_09708_),
    .Y(_02944_));
 TAPCELL_ASAP7_75t_R TAP_560 ();
 NOR2x1_ASAP7_75t_R _28212_ (.A(_00884_),
    .B(_09665_),
    .Y(_09710_));
 AO21x1_ASAP7_75t_R _28213_ (.A1(_08187_),
    .A2(_09665_),
    .B(_09710_),
    .Y(_02945_));
 TAPCELL_ASAP7_75t_R TAP_559 ();
 TAPCELL_ASAP7_75t_R TAP_558 ();
 NOR2x1_ASAP7_75t_R _28216_ (.A(_00916_),
    .B(_09665_),
    .Y(_09713_));
 AO21x1_ASAP7_75t_R _28217_ (.A1(_08219_),
    .A2(_09665_),
    .B(_09713_),
    .Y(_02946_));
 TAPCELL_ASAP7_75t_R TAP_557 ();
 NOR2x1_ASAP7_75t_R _28219_ (.A(_00949_),
    .B(_09665_),
    .Y(_09715_));
 AO21x1_ASAP7_75t_R _28220_ (.A1(_08254_),
    .A2(_09665_),
    .B(_09715_),
    .Y(_02947_));
 TAPCELL_ASAP7_75t_R TAP_556 ();
 NOR2x1_ASAP7_75t_R _28222_ (.A(_00981_),
    .B(_09665_),
    .Y(_09717_));
 AO21x1_ASAP7_75t_R _28223_ (.A1(_08287_),
    .A2(_09665_),
    .B(_09717_),
    .Y(_02948_));
 TAPCELL_ASAP7_75t_R TAP_555 ();
 NOR2x1_ASAP7_75t_R _28225_ (.A(_01015_),
    .B(_09665_),
    .Y(_09719_));
 AO21x1_ASAP7_75t_R _28226_ (.A1(_08319_),
    .A2(_09665_),
    .B(_09719_),
    .Y(_02949_));
 TAPCELL_ASAP7_75t_R TAP_554 ();
 NOR2x1_ASAP7_75t_R _28228_ (.A(_01047_),
    .B(_09665_),
    .Y(_09721_));
 AO21x1_ASAP7_75t_R _28229_ (.A1(_08357_),
    .A2(_09665_),
    .B(_09721_),
    .Y(_02950_));
 TAPCELL_ASAP7_75t_R TAP_553 ();
 NOR2x1_ASAP7_75t_R _28231_ (.A(_01080_),
    .B(_09665_),
    .Y(_09723_));
 AO21x1_ASAP7_75t_R _28232_ (.A1(_08388_),
    .A2(_09665_),
    .B(_09723_),
    .Y(_02951_));
 TAPCELL_ASAP7_75t_R TAP_552 ();
 NOR2x1_ASAP7_75t_R _28234_ (.A(_01112_),
    .B(_09665_),
    .Y(_09725_));
 AO21x1_ASAP7_75t_R _28235_ (.A1(_08419_),
    .A2(_09665_),
    .B(_09725_),
    .Y(_02952_));
 TAPCELL_ASAP7_75t_R TAP_551 ();
 NOR2x1_ASAP7_75t_R _28237_ (.A(_01146_),
    .B(_09665_),
    .Y(_09727_));
 AO21x1_ASAP7_75t_R _28238_ (.A1(_08451_),
    .A2(_09665_),
    .B(_09727_),
    .Y(_02953_));
 TAPCELL_ASAP7_75t_R TAP_550 ();
 NOR2x1_ASAP7_75t_R _28240_ (.A(_01178_),
    .B(_09665_),
    .Y(_09729_));
 AO21x1_ASAP7_75t_R _28241_ (.A1(_08481_),
    .A2(_09665_),
    .B(_09729_),
    .Y(_02954_));
 TAPCELL_ASAP7_75t_R PHY_549 ();
 NOR2x1_ASAP7_75t_R _28243_ (.A(_01212_),
    .B(_09665_),
    .Y(_09731_));
 AO21x1_ASAP7_75t_R _28244_ (.A1(_08512_),
    .A2(_09665_),
    .B(_09731_),
    .Y(_02955_));
 TAPCELL_ASAP7_75t_R PHY_548 ();
 NOR2x1_ASAP7_75t_R _28246_ (.A(_01244_),
    .B(_09665_),
    .Y(_09733_));
 AO21x1_ASAP7_75t_R _28247_ (.A1(_08545_),
    .A2(_09665_),
    .B(_09733_),
    .Y(_02956_));
 TAPCELL_ASAP7_75t_R PHY_547 ();
 NOR2x1_ASAP7_75t_R _28249_ (.A(_01278_),
    .B(_09665_),
    .Y(_09735_));
 AO21x1_ASAP7_75t_R _28250_ (.A1(_08573_),
    .A2(_09665_),
    .B(_09735_),
    .Y(_02957_));
 NOR2x2_ASAP7_75t_R _28251_ (.A(_00323_),
    .B(_00184_),
    .Y(_09736_));
 AND3x2_ASAP7_75t_R _28252_ (.A(_00194_),
    .B(_06922_),
    .C(_09736_),
    .Y(_09737_));
 AND2x6_ASAP7_75t_R _28253_ (.A(_06881_),
    .B(_09737_),
    .Y(_09738_));
 TAPCELL_ASAP7_75t_R PHY_546 ();
 TAPCELL_ASAP7_75t_R PHY_545 ();
 TAPCELL_ASAP7_75t_R PHY_544 ();
 NOR2x1_ASAP7_75t_R _28257_ (.A(_00294_),
    .B(_09738_),
    .Y(_09742_));
 AO21x1_ASAP7_75t_R _28258_ (.A1(_07180_),
    .A2(_09738_),
    .B(_09742_),
    .Y(_02958_));
 NOR2x1_ASAP7_75t_R _28259_ (.A(_00248_),
    .B(_09738_),
    .Y(_09743_));
 AO21x1_ASAP7_75t_R _28260_ (.A1(_07313_),
    .A2(_09738_),
    .B(_09743_),
    .Y(_02959_));
 NOR2x1_ASAP7_75t_R _28261_ (.A(_00356_),
    .B(_09738_),
    .Y(_09744_));
 AO21x1_ASAP7_75t_R _28262_ (.A1(_07398_),
    .A2(_09738_),
    .B(_09744_),
    .Y(_02960_));
 NOR2x1_ASAP7_75t_R _28263_ (.A(_00387_),
    .B(_09738_),
    .Y(_09745_));
 AO21x1_ASAP7_75t_R _28264_ (.A1(_07469_),
    .A2(_09738_),
    .B(_09745_),
    .Y(_02961_));
 NOR2x1_ASAP7_75t_R _28265_ (.A(_00417_),
    .B(_09738_),
    .Y(_09746_));
 AO21x1_ASAP7_75t_R _28266_ (.A1(_07534_),
    .A2(_09738_),
    .B(_09746_),
    .Y(_02962_));
 NOR2x1_ASAP7_75t_R _28267_ (.A(_00447_),
    .B(_09738_),
    .Y(_09747_));
 AO21x1_ASAP7_75t_R _28268_ (.A1(_07581_),
    .A2(_09738_),
    .B(_09747_),
    .Y(_02963_));
 NOR2x1_ASAP7_75t_R _28269_ (.A(_00477_),
    .B(_09738_),
    .Y(_09748_));
 AO21x1_ASAP7_75t_R _28270_ (.A1(net253),
    .A2(_09738_),
    .B(_09748_),
    .Y(_02964_));
 NOR2x1_ASAP7_75t_R _28271_ (.A(_00507_),
    .B(_09738_),
    .Y(_09749_));
 AO21x1_ASAP7_75t_R _28272_ (.A1(_07676_),
    .A2(_09738_),
    .B(_09749_),
    .Y(_02965_));
 TAPCELL_ASAP7_75t_R PHY_543 ();
 NOR2x1_ASAP7_75t_R _28274_ (.A(_00537_),
    .B(_09738_),
    .Y(_09751_));
 AO21x1_ASAP7_75t_R _28275_ (.A1(net252),
    .A2(_09738_),
    .B(_09751_),
    .Y(_02966_));
 NOR2x1_ASAP7_75t_R _28276_ (.A(_00567_),
    .B(_09738_),
    .Y(_09752_));
 AO21x1_ASAP7_75t_R _28277_ (.A1(_07780_),
    .A2(_09738_),
    .B(_09752_),
    .Y(_02967_));
 TAPCELL_ASAP7_75t_R PHY_542 ();
 NOR2x1_ASAP7_75t_R _28279_ (.A(_00597_),
    .B(_09738_),
    .Y(_09754_));
 AO21x1_ASAP7_75t_R _28280_ (.A1(_07817_),
    .A2(_09738_),
    .B(_09754_),
    .Y(_02968_));
 NOR2x1_ASAP7_75t_R _28281_ (.A(_00627_),
    .B(_09738_),
    .Y(_09755_));
 AO21x1_ASAP7_75t_R _28282_ (.A1(_07865_),
    .A2(_09738_),
    .B(_09755_),
    .Y(_02969_));
 NOR2x1_ASAP7_75t_R _28283_ (.A(_00326_),
    .B(_09738_),
    .Y(_09756_));
 AO21x1_ASAP7_75t_R _28284_ (.A1(_07908_),
    .A2(_09738_),
    .B(_09756_),
    .Y(_02970_));
 NOR2x1_ASAP7_75t_R _28285_ (.A(_00689_),
    .B(_09738_),
    .Y(_09757_));
 AO21x1_ASAP7_75t_R _28286_ (.A1(_07950_),
    .A2(_09738_),
    .B(_09757_),
    .Y(_02971_));
 NOR2x1_ASAP7_75t_R _28287_ (.A(_00721_),
    .B(_09738_),
    .Y(_09758_));
 AO21x1_ASAP7_75t_R _28288_ (.A1(_07990_),
    .A2(_09738_),
    .B(_09758_),
    .Y(_02972_));
 NOR2x1_ASAP7_75t_R _28289_ (.A(_00754_),
    .B(_09738_),
    .Y(_09759_));
 AO21x1_ASAP7_75t_R _28290_ (.A1(_08034_),
    .A2(_09738_),
    .B(_09759_),
    .Y(_02973_));
 NOR2x1_ASAP7_75t_R _28291_ (.A(_00787_),
    .B(_09738_),
    .Y(_09760_));
 AO21x1_ASAP7_75t_R _28292_ (.A1(_08073_),
    .A2(_09738_),
    .B(_09760_),
    .Y(_02974_));
 NOR2x1_ASAP7_75t_R _28293_ (.A(_00820_),
    .B(_09738_),
    .Y(_09761_));
 AO21x1_ASAP7_75t_R _28294_ (.A1(_08116_),
    .A2(_09738_),
    .B(_09761_),
    .Y(_02975_));
 TAPCELL_ASAP7_75t_R PHY_541 ();
 NOR2x1_ASAP7_75t_R _28296_ (.A(_00852_),
    .B(_09738_),
    .Y(_09763_));
 AO21x1_ASAP7_75t_R _28297_ (.A1(_08150_),
    .A2(_09738_),
    .B(_09763_),
    .Y(_02976_));
 NOR2x1_ASAP7_75t_R _28298_ (.A(_00885_),
    .B(_09738_),
    .Y(_09764_));
 AO21x1_ASAP7_75t_R _28299_ (.A1(_08187_),
    .A2(_09738_),
    .B(_09764_),
    .Y(_02977_));
 TAPCELL_ASAP7_75t_R PHY_540 ();
 NOR2x1_ASAP7_75t_R _28301_ (.A(_00917_),
    .B(_09738_),
    .Y(_09766_));
 AO21x1_ASAP7_75t_R _28302_ (.A1(_08219_),
    .A2(_09738_),
    .B(_09766_),
    .Y(_02978_));
 NOR2x1_ASAP7_75t_R _28303_ (.A(_00950_),
    .B(_09738_),
    .Y(_09767_));
 AO21x1_ASAP7_75t_R _28304_ (.A1(_08254_),
    .A2(_09738_),
    .B(_09767_),
    .Y(_02979_));
 NOR2x1_ASAP7_75t_R _28305_ (.A(_00982_),
    .B(_09738_),
    .Y(_09768_));
 AO21x1_ASAP7_75t_R _28306_ (.A1(_08287_),
    .A2(_09738_),
    .B(_09768_),
    .Y(_02980_));
 NOR2x1_ASAP7_75t_R _28307_ (.A(_01016_),
    .B(_09738_),
    .Y(_09769_));
 AO21x1_ASAP7_75t_R _28308_ (.A1(_08319_),
    .A2(_09738_),
    .B(_09769_),
    .Y(_02981_));
 NOR2x1_ASAP7_75t_R _28309_ (.A(_01048_),
    .B(_09738_),
    .Y(_09770_));
 AO21x1_ASAP7_75t_R _28310_ (.A1(_08357_),
    .A2(_09738_),
    .B(_09770_),
    .Y(_02982_));
 NOR2x1_ASAP7_75t_R _28311_ (.A(_01081_),
    .B(_09738_),
    .Y(_09771_));
 AO21x1_ASAP7_75t_R _28312_ (.A1(_08388_),
    .A2(_09738_),
    .B(_09771_),
    .Y(_02983_));
 NOR2x1_ASAP7_75t_R _28313_ (.A(_01113_),
    .B(_09738_),
    .Y(_09772_));
 AO21x1_ASAP7_75t_R _28314_ (.A1(_08419_),
    .A2(_09738_),
    .B(_09772_),
    .Y(_02984_));
 NOR2x1_ASAP7_75t_R _28315_ (.A(_01147_),
    .B(_09738_),
    .Y(_09773_));
 AO21x1_ASAP7_75t_R _28316_ (.A1(_08451_),
    .A2(_09738_),
    .B(_09773_),
    .Y(_02985_));
 NOR2x1_ASAP7_75t_R _28317_ (.A(_01179_),
    .B(_09738_),
    .Y(_09774_));
 AO21x1_ASAP7_75t_R _28318_ (.A1(_08481_),
    .A2(_09738_),
    .B(_09774_),
    .Y(_02986_));
 NOR2x1_ASAP7_75t_R _28319_ (.A(_01213_),
    .B(_09738_),
    .Y(_09775_));
 AO21x1_ASAP7_75t_R _28320_ (.A1(_08512_),
    .A2(_09738_),
    .B(_09775_),
    .Y(_02987_));
 NOR2x1_ASAP7_75t_R _28321_ (.A(_01245_),
    .B(_09738_),
    .Y(_09776_));
 AO21x1_ASAP7_75t_R _28322_ (.A1(_08545_),
    .A2(_09738_),
    .B(_09776_),
    .Y(_02988_));
 NOR2x1_ASAP7_75t_R _28323_ (.A(_01279_),
    .B(_09738_),
    .Y(_09777_));
 AO21x1_ASAP7_75t_R _28324_ (.A1(_08573_),
    .A2(_09738_),
    .B(_09777_),
    .Y(_02989_));
 AND2x2_ASAP7_75t_R _28325_ (.A(_00194_),
    .B(_06922_),
    .Y(_09778_));
 AND2x6_ASAP7_75t_R _28326_ (.A(_13950_),
    .B(_00191_),
    .Y(_09779_));
 AND4x2_ASAP7_75t_R _28327_ (.A(_00323_),
    .B(_00184_),
    .C(_09778_),
    .D(_09779_),
    .Y(_09780_));
 TAPCELL_ASAP7_75t_R PHY_539 ();
 TAPCELL_ASAP7_75t_R PHY_538 ();
 TAPCELL_ASAP7_75t_R PHY_537 ();
 NOR2x1_ASAP7_75t_R _28331_ (.A(_00295_),
    .B(net270),
    .Y(_09784_));
 AO21x1_ASAP7_75t_R _28332_ (.A1(_07180_),
    .A2(net270),
    .B(_09784_),
    .Y(_02990_));
 NOR2x1_ASAP7_75t_R _28333_ (.A(_00249_),
    .B(net270),
    .Y(_09785_));
 AO21x1_ASAP7_75t_R _28334_ (.A1(_07313_),
    .A2(net270),
    .B(_09785_),
    .Y(_02991_));
 NOR2x1_ASAP7_75t_R _28335_ (.A(_00357_),
    .B(net270),
    .Y(_09786_));
 AO21x1_ASAP7_75t_R _28336_ (.A1(_07398_),
    .A2(net270),
    .B(_09786_),
    .Y(_02992_));
 NOR2x1_ASAP7_75t_R _28337_ (.A(_00388_),
    .B(net270),
    .Y(_09787_));
 AO21x1_ASAP7_75t_R _28338_ (.A1(_07469_),
    .A2(net270),
    .B(_09787_),
    .Y(_02993_));
 NOR2x1_ASAP7_75t_R _28339_ (.A(_00418_),
    .B(_09780_),
    .Y(_09788_));
 AO21x1_ASAP7_75t_R _28340_ (.A1(_07534_),
    .A2(_09780_),
    .B(_09788_),
    .Y(_02994_));
 NOR2x1_ASAP7_75t_R _28341_ (.A(_00448_),
    .B(net270),
    .Y(_09789_));
 AO21x1_ASAP7_75t_R _28342_ (.A1(_07581_),
    .A2(net270),
    .B(_09789_),
    .Y(_02995_));
 NOR2x1_ASAP7_75t_R _28343_ (.A(_00478_),
    .B(_09780_),
    .Y(_09790_));
 AO21x1_ASAP7_75t_R _28344_ (.A1(net253),
    .A2(_09780_),
    .B(_09790_),
    .Y(_02996_));
 NOR2x1_ASAP7_75t_R _28345_ (.A(_00508_),
    .B(net270),
    .Y(_09791_));
 AO21x1_ASAP7_75t_R _28346_ (.A1(_07676_),
    .A2(net270),
    .B(_09791_),
    .Y(_02997_));
 TAPCELL_ASAP7_75t_R PHY_536 ();
 NOR2x1_ASAP7_75t_R _28348_ (.A(_00538_),
    .B(_09780_),
    .Y(_09793_));
 AO21x1_ASAP7_75t_R _28349_ (.A1(_07738_),
    .A2(_09780_),
    .B(_09793_),
    .Y(_02998_));
 NOR2x1_ASAP7_75t_R _28350_ (.A(_00568_),
    .B(_09780_),
    .Y(_09794_));
 AO21x1_ASAP7_75t_R _28351_ (.A1(_07780_),
    .A2(_09780_),
    .B(_09794_),
    .Y(_02999_));
 TAPCELL_ASAP7_75t_R PHY_535 ();
 NOR2x1_ASAP7_75t_R _28353_ (.A(_00598_),
    .B(net269),
    .Y(_09796_));
 AO21x1_ASAP7_75t_R _28354_ (.A1(_07817_),
    .A2(net269),
    .B(_09796_),
    .Y(_03000_));
 NOR2x1_ASAP7_75t_R _28355_ (.A(_00628_),
    .B(net270),
    .Y(_09797_));
 AO21x1_ASAP7_75t_R _28356_ (.A1(_07865_),
    .A2(net270),
    .B(_09797_),
    .Y(_03001_));
 NOR2x1_ASAP7_75t_R _28357_ (.A(_00327_),
    .B(net270),
    .Y(_09798_));
 AO21x1_ASAP7_75t_R _28358_ (.A1(_07908_),
    .A2(net270),
    .B(_09798_),
    .Y(_03002_));
 NOR2x1_ASAP7_75t_R _28359_ (.A(_00690_),
    .B(net269),
    .Y(_09799_));
 AO21x1_ASAP7_75t_R _28360_ (.A1(_07950_),
    .A2(net269),
    .B(_09799_),
    .Y(_03003_));
 NOR2x1_ASAP7_75t_R _28361_ (.A(_00722_),
    .B(_09780_),
    .Y(_09800_));
 AO21x1_ASAP7_75t_R _28362_ (.A1(_07990_),
    .A2(_09780_),
    .B(_09800_),
    .Y(_03004_));
 NOR2x1_ASAP7_75t_R _28363_ (.A(_00755_),
    .B(net269),
    .Y(_09801_));
 AO21x1_ASAP7_75t_R _28364_ (.A1(_08034_),
    .A2(net269),
    .B(_09801_),
    .Y(_03005_));
 NOR2x1_ASAP7_75t_R _28365_ (.A(_00788_),
    .B(net269),
    .Y(_09802_));
 AO21x1_ASAP7_75t_R _28366_ (.A1(_08073_),
    .A2(net269),
    .B(_09802_),
    .Y(_03006_));
 NOR2x1_ASAP7_75t_R _28367_ (.A(_00821_),
    .B(net269),
    .Y(_09803_));
 AO21x1_ASAP7_75t_R _28368_ (.A1(_08116_),
    .A2(net269),
    .B(_09803_),
    .Y(_03007_));
 TAPCELL_ASAP7_75t_R PHY_534 ();
 NOR2x1_ASAP7_75t_R _28370_ (.A(_00853_),
    .B(net270),
    .Y(_09805_));
 AO21x1_ASAP7_75t_R _28371_ (.A1(_08150_),
    .A2(net270),
    .B(_09805_),
    .Y(_03008_));
 NOR2x1_ASAP7_75t_R _28372_ (.A(_00886_),
    .B(net269),
    .Y(_09806_));
 AO21x1_ASAP7_75t_R _28373_ (.A1(_08187_),
    .A2(net269),
    .B(_09806_),
    .Y(_03009_));
 TAPCELL_ASAP7_75t_R PHY_533 ();
 NOR2x1_ASAP7_75t_R _28375_ (.A(_00918_),
    .B(net269),
    .Y(_09808_));
 AO21x1_ASAP7_75t_R _28376_ (.A1(_08219_),
    .A2(net269),
    .B(_09808_),
    .Y(_03010_));
 NOR2x1_ASAP7_75t_R _28377_ (.A(_00951_),
    .B(net269),
    .Y(_09809_));
 AO21x1_ASAP7_75t_R _28378_ (.A1(_08254_),
    .A2(net269),
    .B(_09809_),
    .Y(_03011_));
 NOR2x1_ASAP7_75t_R _28379_ (.A(_00983_),
    .B(_09780_),
    .Y(_09810_));
 AO21x1_ASAP7_75t_R _28380_ (.A1(net250),
    .A2(_09780_),
    .B(_09810_),
    .Y(_03012_));
 NOR2x1_ASAP7_75t_R _28381_ (.A(_01017_),
    .B(net270),
    .Y(_09811_));
 AO21x1_ASAP7_75t_R _28382_ (.A1(_08319_),
    .A2(net270),
    .B(_09811_),
    .Y(_03013_));
 NOR2x1_ASAP7_75t_R _28383_ (.A(_01049_),
    .B(net269),
    .Y(_09812_));
 AO21x1_ASAP7_75t_R _28384_ (.A1(_08357_),
    .A2(net269),
    .B(_09812_),
    .Y(_03014_));
 NOR2x1_ASAP7_75t_R _28385_ (.A(_01082_),
    .B(net269),
    .Y(_09813_));
 AO21x1_ASAP7_75t_R _28386_ (.A1(_08388_),
    .A2(net269),
    .B(_09813_),
    .Y(_03015_));
 NOR2x1_ASAP7_75t_R _28387_ (.A(_01114_),
    .B(net269),
    .Y(_09814_));
 AO21x1_ASAP7_75t_R _28388_ (.A1(_08419_),
    .A2(net269),
    .B(_09814_),
    .Y(_03016_));
 NOR2x1_ASAP7_75t_R _28389_ (.A(_01148_),
    .B(net269),
    .Y(_09815_));
 AO21x1_ASAP7_75t_R _28390_ (.A1(_08451_),
    .A2(net269),
    .B(_09815_),
    .Y(_03017_));
 NOR2x1_ASAP7_75t_R _28391_ (.A(_01180_),
    .B(_09780_),
    .Y(_09816_));
 AO21x1_ASAP7_75t_R _28392_ (.A1(_08481_),
    .A2(_09780_),
    .B(_09816_),
    .Y(_03018_));
 NOR2x1_ASAP7_75t_R _28393_ (.A(_01214_),
    .B(net270),
    .Y(_09817_));
 AO21x1_ASAP7_75t_R _28394_ (.A1(_08512_),
    .A2(net270),
    .B(_09817_),
    .Y(_03019_));
 NOR2x1_ASAP7_75t_R _28395_ (.A(_01246_),
    .B(net269),
    .Y(_09818_));
 AO21x1_ASAP7_75t_R _28396_ (.A1(_08545_),
    .A2(net269),
    .B(_09818_),
    .Y(_03020_));
 NOR2x1_ASAP7_75t_R _28397_ (.A(_01280_),
    .B(net270),
    .Y(_09819_));
 AO21x1_ASAP7_75t_R _28398_ (.A1(_08573_),
    .A2(net270),
    .B(_09819_),
    .Y(_03021_));
 AND2x6_ASAP7_75t_R _28399_ (.A(_06923_),
    .B(_09779_),
    .Y(_09820_));
 TAPCELL_ASAP7_75t_R PHY_532 ();
 TAPCELL_ASAP7_75t_R PHY_531 ();
 TAPCELL_ASAP7_75t_R PHY_530 ();
 NOR2x1_ASAP7_75t_R _28403_ (.A(_00296_),
    .B(_09820_),
    .Y(_09824_));
 AO21x1_ASAP7_75t_R _28404_ (.A1(_07180_),
    .A2(_09820_),
    .B(_09824_),
    .Y(_03022_));
 NOR2x1_ASAP7_75t_R _28405_ (.A(_00250_),
    .B(_09820_),
    .Y(_09825_));
 AO21x1_ASAP7_75t_R _28406_ (.A1(_07313_),
    .A2(_09820_),
    .B(_09825_),
    .Y(_03023_));
 NOR2x1_ASAP7_75t_R _28407_ (.A(_00358_),
    .B(_09820_),
    .Y(_09826_));
 AO21x1_ASAP7_75t_R _28408_ (.A1(_07398_),
    .A2(_09820_),
    .B(_09826_),
    .Y(_03024_));
 NOR2x1_ASAP7_75t_R _28409_ (.A(_00389_),
    .B(_09820_),
    .Y(_09827_));
 AO21x1_ASAP7_75t_R _28410_ (.A1(_07469_),
    .A2(_09820_),
    .B(_09827_),
    .Y(_03025_));
 NOR2x1_ASAP7_75t_R _28411_ (.A(_00419_),
    .B(_09820_),
    .Y(_09828_));
 AO21x1_ASAP7_75t_R _28412_ (.A1(_07534_),
    .A2(_09820_),
    .B(_09828_),
    .Y(_03026_));
 NOR2x1_ASAP7_75t_R _28413_ (.A(_00449_),
    .B(_09820_),
    .Y(_09829_));
 AO21x1_ASAP7_75t_R _28414_ (.A1(_07581_),
    .A2(_09820_),
    .B(_09829_),
    .Y(_03027_));
 NOR2x1_ASAP7_75t_R _28415_ (.A(_00479_),
    .B(_09820_),
    .Y(_09830_));
 AO21x1_ASAP7_75t_R _28416_ (.A1(net253),
    .A2(_09820_),
    .B(_09830_),
    .Y(_03028_));
 NOR2x1_ASAP7_75t_R _28417_ (.A(_00509_),
    .B(_09820_),
    .Y(_09831_));
 AO21x1_ASAP7_75t_R _28418_ (.A1(_07676_),
    .A2(_09820_),
    .B(_09831_),
    .Y(_03029_));
 TAPCELL_ASAP7_75t_R PHY_529 ();
 NOR2x1_ASAP7_75t_R _28420_ (.A(_00539_),
    .B(_09820_),
    .Y(_09833_));
 AO21x1_ASAP7_75t_R _28421_ (.A1(_07738_),
    .A2(_09820_),
    .B(_09833_),
    .Y(_03030_));
 NOR2x1_ASAP7_75t_R _28422_ (.A(_00569_),
    .B(_09820_),
    .Y(_09834_));
 AO21x1_ASAP7_75t_R _28423_ (.A1(_07780_),
    .A2(_09820_),
    .B(_09834_),
    .Y(_03031_));
 TAPCELL_ASAP7_75t_R PHY_528 ();
 NOR2x1_ASAP7_75t_R _28425_ (.A(_00599_),
    .B(_09820_),
    .Y(_09836_));
 AO21x1_ASAP7_75t_R _28426_ (.A1(_07817_),
    .A2(_09820_),
    .B(_09836_),
    .Y(_03032_));
 NOR2x1_ASAP7_75t_R _28427_ (.A(_00629_),
    .B(_09820_),
    .Y(_09837_));
 AO21x1_ASAP7_75t_R _28428_ (.A1(_07865_),
    .A2(_09820_),
    .B(_09837_),
    .Y(_03033_));
 NOR2x1_ASAP7_75t_R _28429_ (.A(_00328_),
    .B(_09820_),
    .Y(_09838_));
 AO21x1_ASAP7_75t_R _28430_ (.A1(_07908_),
    .A2(_09820_),
    .B(_09838_),
    .Y(_03034_));
 NOR2x1_ASAP7_75t_R _28431_ (.A(_00691_),
    .B(_09820_),
    .Y(_09839_));
 AO21x1_ASAP7_75t_R _28432_ (.A1(_07950_),
    .A2(_09820_),
    .B(_09839_),
    .Y(_03035_));
 NOR2x1_ASAP7_75t_R _28433_ (.A(_00723_),
    .B(_09820_),
    .Y(_09840_));
 AO21x1_ASAP7_75t_R _28434_ (.A1(_07990_),
    .A2(_09820_),
    .B(_09840_),
    .Y(_03036_));
 NOR2x1_ASAP7_75t_R _28435_ (.A(_00756_),
    .B(_09820_),
    .Y(_09841_));
 AO21x1_ASAP7_75t_R _28436_ (.A1(_08034_),
    .A2(_09820_),
    .B(_09841_),
    .Y(_03037_));
 NOR2x1_ASAP7_75t_R _28437_ (.A(_00789_),
    .B(_09820_),
    .Y(_09842_));
 AO21x1_ASAP7_75t_R _28438_ (.A1(_08073_),
    .A2(_09820_),
    .B(_09842_),
    .Y(_03038_));
 NOR2x1_ASAP7_75t_R _28439_ (.A(_00822_),
    .B(_09820_),
    .Y(_09843_));
 AO21x1_ASAP7_75t_R _28440_ (.A1(_08116_),
    .A2(_09820_),
    .B(_09843_),
    .Y(_03039_));
 TAPCELL_ASAP7_75t_R PHY_527 ();
 NOR2x1_ASAP7_75t_R _28442_ (.A(_00854_),
    .B(_09820_),
    .Y(_09845_));
 AO21x1_ASAP7_75t_R _28443_ (.A1(_08150_),
    .A2(_09820_),
    .B(_09845_),
    .Y(_03040_));
 NOR2x1_ASAP7_75t_R _28444_ (.A(_00887_),
    .B(_09820_),
    .Y(_09846_));
 AO21x1_ASAP7_75t_R _28445_ (.A1(_08187_),
    .A2(_09820_),
    .B(_09846_),
    .Y(_03041_));
 TAPCELL_ASAP7_75t_R PHY_526 ();
 NOR2x1_ASAP7_75t_R _28447_ (.A(_00919_),
    .B(_09820_),
    .Y(_09848_));
 AO21x1_ASAP7_75t_R _28448_ (.A1(_08219_),
    .A2(_09820_),
    .B(_09848_),
    .Y(_03042_));
 NOR2x1_ASAP7_75t_R _28449_ (.A(_00952_),
    .B(_09820_),
    .Y(_09849_));
 AO21x1_ASAP7_75t_R _28450_ (.A1(_08254_),
    .A2(_09820_),
    .B(_09849_),
    .Y(_03043_));
 NOR2x1_ASAP7_75t_R _28451_ (.A(_00984_),
    .B(_09820_),
    .Y(_09850_));
 AO21x1_ASAP7_75t_R _28452_ (.A1(net250),
    .A2(_09820_),
    .B(_09850_),
    .Y(_03044_));
 NOR2x1_ASAP7_75t_R _28453_ (.A(_01018_),
    .B(_09820_),
    .Y(_09851_));
 AO21x1_ASAP7_75t_R _28454_ (.A1(_08319_),
    .A2(_09820_),
    .B(_09851_),
    .Y(_03045_));
 NOR2x1_ASAP7_75t_R _28455_ (.A(_01050_),
    .B(_09820_),
    .Y(_09852_));
 AO21x1_ASAP7_75t_R _28456_ (.A1(_08357_),
    .A2(_09820_),
    .B(_09852_),
    .Y(_03046_));
 NOR2x1_ASAP7_75t_R _28457_ (.A(_01083_),
    .B(_09820_),
    .Y(_09853_));
 AO21x1_ASAP7_75t_R _28458_ (.A1(_08388_),
    .A2(_09820_),
    .B(_09853_),
    .Y(_03047_));
 NOR2x1_ASAP7_75t_R _28459_ (.A(_01115_),
    .B(_09820_),
    .Y(_09854_));
 AO21x1_ASAP7_75t_R _28460_ (.A1(_08419_),
    .A2(_09820_),
    .B(_09854_),
    .Y(_03048_));
 NOR2x1_ASAP7_75t_R _28461_ (.A(_01149_),
    .B(_09820_),
    .Y(_09855_));
 AO21x1_ASAP7_75t_R _28462_ (.A1(_08451_),
    .A2(_09820_),
    .B(_09855_),
    .Y(_03049_));
 NOR2x1_ASAP7_75t_R _28463_ (.A(_01181_),
    .B(_09820_),
    .Y(_09856_));
 AO21x1_ASAP7_75t_R _28464_ (.A1(_08481_),
    .A2(_09820_),
    .B(_09856_),
    .Y(_03050_));
 NOR2x1_ASAP7_75t_R _28465_ (.A(_01215_),
    .B(_09820_),
    .Y(_09857_));
 AO21x1_ASAP7_75t_R _28466_ (.A1(_08512_),
    .A2(_09820_),
    .B(_09857_),
    .Y(_03051_));
 NOR2x1_ASAP7_75t_R _28467_ (.A(_01247_),
    .B(_09820_),
    .Y(_09858_));
 AO21x1_ASAP7_75t_R _28468_ (.A1(_08545_),
    .A2(_09820_),
    .B(_09858_),
    .Y(_03052_));
 NOR2x1_ASAP7_75t_R _28469_ (.A(_01281_),
    .B(_09820_),
    .Y(_09859_));
 AO21x1_ASAP7_75t_R _28470_ (.A1(_08573_),
    .A2(_09820_),
    .B(_09859_),
    .Y(_03053_));
 AND2x6_ASAP7_75t_R _28471_ (.A(_09664_),
    .B(_09779_),
    .Y(_09860_));
 TAPCELL_ASAP7_75t_R PHY_525 ();
 TAPCELL_ASAP7_75t_R PHY_524 ();
 TAPCELL_ASAP7_75t_R PHY_523 ();
 NOR2x1_ASAP7_75t_R _28475_ (.A(_00297_),
    .B(_09860_),
    .Y(_09864_));
 AO21x1_ASAP7_75t_R _28476_ (.A1(_07180_),
    .A2(_09860_),
    .B(_09864_),
    .Y(_03054_));
 NOR2x1_ASAP7_75t_R _28477_ (.A(_00251_),
    .B(_09860_),
    .Y(_09865_));
 AO21x1_ASAP7_75t_R _28478_ (.A1(_07313_),
    .A2(_09860_),
    .B(_09865_),
    .Y(_03055_));
 NOR2x1_ASAP7_75t_R _28479_ (.A(_00359_),
    .B(_09860_),
    .Y(_09866_));
 AO21x1_ASAP7_75t_R _28480_ (.A1(_07398_),
    .A2(_09860_),
    .B(_09866_),
    .Y(_03056_));
 NOR2x1_ASAP7_75t_R _28481_ (.A(_00390_),
    .B(_09860_),
    .Y(_09867_));
 AO21x1_ASAP7_75t_R _28482_ (.A1(_07469_),
    .A2(_09860_),
    .B(_09867_),
    .Y(_03057_));
 NOR2x1_ASAP7_75t_R _28483_ (.A(_00420_),
    .B(_09860_),
    .Y(_09868_));
 AO21x1_ASAP7_75t_R _28484_ (.A1(_07534_),
    .A2(_09860_),
    .B(_09868_),
    .Y(_03058_));
 NOR2x1_ASAP7_75t_R _28485_ (.A(_00450_),
    .B(_09860_),
    .Y(_09869_));
 AO21x1_ASAP7_75t_R _28486_ (.A1(_07581_),
    .A2(_09860_),
    .B(_09869_),
    .Y(_03059_));
 NOR2x1_ASAP7_75t_R _28487_ (.A(_00480_),
    .B(_09860_),
    .Y(_09870_));
 AO21x1_ASAP7_75t_R _28488_ (.A1(net253),
    .A2(_09860_),
    .B(_09870_),
    .Y(_03060_));
 NOR2x1_ASAP7_75t_R _28489_ (.A(_00510_),
    .B(_09860_),
    .Y(_09871_));
 AO21x1_ASAP7_75t_R _28490_ (.A1(_07676_),
    .A2(_09860_),
    .B(_09871_),
    .Y(_03061_));
 TAPCELL_ASAP7_75t_R PHY_522 ();
 NOR2x1_ASAP7_75t_R _28492_ (.A(_00540_),
    .B(_09860_),
    .Y(_09873_));
 AO21x1_ASAP7_75t_R _28493_ (.A1(_07738_),
    .A2(_09860_),
    .B(_09873_),
    .Y(_03062_));
 NOR2x1_ASAP7_75t_R _28494_ (.A(_00570_),
    .B(_09860_),
    .Y(_09874_));
 AO21x1_ASAP7_75t_R _28495_ (.A1(_07780_),
    .A2(_09860_),
    .B(_09874_),
    .Y(_03063_));
 TAPCELL_ASAP7_75t_R PHY_521 ();
 NOR2x1_ASAP7_75t_R _28497_ (.A(_00600_),
    .B(_09860_),
    .Y(_09876_));
 AO21x1_ASAP7_75t_R _28498_ (.A1(_07817_),
    .A2(_09860_),
    .B(_09876_),
    .Y(_03064_));
 NOR2x1_ASAP7_75t_R _28499_ (.A(_00630_),
    .B(_09860_),
    .Y(_09877_));
 AO21x1_ASAP7_75t_R _28500_ (.A1(_07865_),
    .A2(_09860_),
    .B(_09877_),
    .Y(_03065_));
 NOR2x1_ASAP7_75t_R _28501_ (.A(_00329_),
    .B(_09860_),
    .Y(_09878_));
 AO21x1_ASAP7_75t_R _28502_ (.A1(_07908_),
    .A2(_09860_),
    .B(_09878_),
    .Y(_03066_));
 NOR2x1_ASAP7_75t_R _28503_ (.A(_00692_),
    .B(_09860_),
    .Y(_09879_));
 AO21x1_ASAP7_75t_R _28504_ (.A1(_07950_),
    .A2(_09860_),
    .B(_09879_),
    .Y(_03067_));
 NOR2x1_ASAP7_75t_R _28505_ (.A(_00724_),
    .B(_09860_),
    .Y(_09880_));
 AO21x1_ASAP7_75t_R _28506_ (.A1(_07990_),
    .A2(_09860_),
    .B(_09880_),
    .Y(_03068_));
 NOR2x1_ASAP7_75t_R _28507_ (.A(_00757_),
    .B(_09860_),
    .Y(_09881_));
 AO21x1_ASAP7_75t_R _28508_ (.A1(_08034_),
    .A2(_09860_),
    .B(_09881_),
    .Y(_03069_));
 NOR2x1_ASAP7_75t_R _28509_ (.A(_00790_),
    .B(_09860_),
    .Y(_09882_));
 AO21x1_ASAP7_75t_R _28510_ (.A1(_08073_),
    .A2(_09860_),
    .B(_09882_),
    .Y(_03070_));
 NOR2x1_ASAP7_75t_R _28511_ (.A(_00823_),
    .B(_09860_),
    .Y(_09883_));
 AO21x1_ASAP7_75t_R _28512_ (.A1(_08116_),
    .A2(_09860_),
    .B(_09883_),
    .Y(_03071_));
 TAPCELL_ASAP7_75t_R PHY_520 ();
 NOR2x1_ASAP7_75t_R _28514_ (.A(_00855_),
    .B(_09860_),
    .Y(_09885_));
 AO21x1_ASAP7_75t_R _28515_ (.A1(_08150_),
    .A2(_09860_),
    .B(_09885_),
    .Y(_03072_));
 NOR2x1_ASAP7_75t_R _28516_ (.A(_00888_),
    .B(_09860_),
    .Y(_09886_));
 AO21x1_ASAP7_75t_R _28517_ (.A1(_08187_),
    .A2(_09860_),
    .B(_09886_),
    .Y(_03073_));
 TAPCELL_ASAP7_75t_R PHY_519 ();
 NOR2x1_ASAP7_75t_R _28519_ (.A(_00920_),
    .B(_09860_),
    .Y(_09888_));
 AO21x1_ASAP7_75t_R _28520_ (.A1(_08219_),
    .A2(_09860_),
    .B(_09888_),
    .Y(_03074_));
 NOR2x1_ASAP7_75t_R _28521_ (.A(_00953_),
    .B(_09860_),
    .Y(_09889_));
 AO21x1_ASAP7_75t_R _28522_ (.A1(_08254_),
    .A2(_09860_),
    .B(_09889_),
    .Y(_03075_));
 NOR2x1_ASAP7_75t_R _28523_ (.A(_00985_),
    .B(_09860_),
    .Y(_09890_));
 AO21x1_ASAP7_75t_R _28524_ (.A1(net250),
    .A2(_09860_),
    .B(_09890_),
    .Y(_03076_));
 NOR2x1_ASAP7_75t_R _28525_ (.A(_01019_),
    .B(_09860_),
    .Y(_09891_));
 AO21x1_ASAP7_75t_R _28526_ (.A1(_08319_),
    .A2(_09860_),
    .B(_09891_),
    .Y(_03077_));
 NOR2x1_ASAP7_75t_R _28527_ (.A(_01051_),
    .B(_09860_),
    .Y(_09892_));
 AO21x1_ASAP7_75t_R _28528_ (.A1(_08357_),
    .A2(_09860_),
    .B(_09892_),
    .Y(_03078_));
 NOR2x1_ASAP7_75t_R _28529_ (.A(_01084_),
    .B(_09860_),
    .Y(_09893_));
 AO21x1_ASAP7_75t_R _28530_ (.A1(_08388_),
    .A2(_09860_),
    .B(_09893_),
    .Y(_03079_));
 NOR2x1_ASAP7_75t_R _28531_ (.A(_01116_),
    .B(_09860_),
    .Y(_09894_));
 AO21x1_ASAP7_75t_R _28532_ (.A1(_08419_),
    .A2(_09860_),
    .B(_09894_),
    .Y(_03080_));
 NOR2x1_ASAP7_75t_R _28533_ (.A(_01150_),
    .B(_09860_),
    .Y(_09895_));
 AO21x1_ASAP7_75t_R _28534_ (.A1(_08451_),
    .A2(_09860_),
    .B(_09895_),
    .Y(_03081_));
 NOR2x1_ASAP7_75t_R _28535_ (.A(_01182_),
    .B(_09860_),
    .Y(_09896_));
 AO21x1_ASAP7_75t_R _28536_ (.A1(_08481_),
    .A2(_09860_),
    .B(_09896_),
    .Y(_03082_));
 NOR2x1_ASAP7_75t_R _28537_ (.A(_01216_),
    .B(_09860_),
    .Y(_09897_));
 AO21x1_ASAP7_75t_R _28538_ (.A1(_08512_),
    .A2(_09860_),
    .B(_09897_),
    .Y(_03083_));
 NOR2x1_ASAP7_75t_R _28539_ (.A(_01248_),
    .B(_09860_),
    .Y(_09898_));
 AO21x1_ASAP7_75t_R _28540_ (.A1(_08545_),
    .A2(_09860_),
    .B(_09898_),
    .Y(_03084_));
 NOR2x1_ASAP7_75t_R _28541_ (.A(_01282_),
    .B(_09860_),
    .Y(_09899_));
 AO21x1_ASAP7_75t_R _28542_ (.A1(_08573_),
    .A2(_09860_),
    .B(_09899_),
    .Y(_03085_));
 AND2x6_ASAP7_75t_R _28543_ (.A(_09737_),
    .B(_09779_),
    .Y(_09900_));
 TAPCELL_ASAP7_75t_R PHY_518 ();
 TAPCELL_ASAP7_75t_R PHY_517 ();
 TAPCELL_ASAP7_75t_R PHY_516 ();
 NOR2x1_ASAP7_75t_R _28547_ (.A(_00298_),
    .B(_09900_),
    .Y(_09904_));
 AO21x1_ASAP7_75t_R _28548_ (.A1(_07180_),
    .A2(_09900_),
    .B(_09904_),
    .Y(_03086_));
 NOR2x1_ASAP7_75t_R _28549_ (.A(_00252_),
    .B(_09900_),
    .Y(_09905_));
 AO21x1_ASAP7_75t_R _28550_ (.A1(_07313_),
    .A2(_09900_),
    .B(_09905_),
    .Y(_03087_));
 NOR2x1_ASAP7_75t_R _28551_ (.A(_00360_),
    .B(_09900_),
    .Y(_09906_));
 AO21x1_ASAP7_75t_R _28552_ (.A1(_07398_),
    .A2(_09900_),
    .B(_09906_),
    .Y(_03088_));
 NOR2x1_ASAP7_75t_R _28553_ (.A(_00391_),
    .B(_09900_),
    .Y(_09907_));
 AO21x1_ASAP7_75t_R _28554_ (.A1(_07469_),
    .A2(_09900_),
    .B(_09907_),
    .Y(_03089_));
 NOR2x1_ASAP7_75t_R _28555_ (.A(_00421_),
    .B(_09900_),
    .Y(_09908_));
 AO21x1_ASAP7_75t_R _28556_ (.A1(_07534_),
    .A2(_09900_),
    .B(_09908_),
    .Y(_03090_));
 NOR2x1_ASAP7_75t_R _28557_ (.A(_00451_),
    .B(_09900_),
    .Y(_09909_));
 AO21x1_ASAP7_75t_R _28558_ (.A1(_07581_),
    .A2(_09900_),
    .B(_09909_),
    .Y(_03091_));
 NOR2x1_ASAP7_75t_R _28559_ (.A(_00481_),
    .B(_09900_),
    .Y(_09910_));
 AO21x1_ASAP7_75t_R _28560_ (.A1(net253),
    .A2(_09900_),
    .B(_09910_),
    .Y(_03092_));
 NOR2x1_ASAP7_75t_R _28561_ (.A(_00511_),
    .B(_09900_),
    .Y(_09911_));
 AO21x1_ASAP7_75t_R _28562_ (.A1(_07676_),
    .A2(_09900_),
    .B(_09911_),
    .Y(_03093_));
 TAPCELL_ASAP7_75t_R PHY_515 ();
 NOR2x1_ASAP7_75t_R _28564_ (.A(_00541_),
    .B(_09900_),
    .Y(_09913_));
 AO21x1_ASAP7_75t_R _28565_ (.A1(_07738_),
    .A2(_09900_),
    .B(_09913_),
    .Y(_03094_));
 NOR2x1_ASAP7_75t_R _28566_ (.A(_00571_),
    .B(_09900_),
    .Y(_09914_));
 AO21x1_ASAP7_75t_R _28567_ (.A1(_07780_),
    .A2(_09900_),
    .B(_09914_),
    .Y(_03095_));
 TAPCELL_ASAP7_75t_R PHY_514 ();
 NOR2x1_ASAP7_75t_R _28569_ (.A(_00601_),
    .B(_09900_),
    .Y(_09916_));
 AO21x1_ASAP7_75t_R _28570_ (.A1(_07817_),
    .A2(_09900_),
    .B(_09916_),
    .Y(_03096_));
 NOR2x1_ASAP7_75t_R _28571_ (.A(_00631_),
    .B(_09900_),
    .Y(_09917_));
 AO21x1_ASAP7_75t_R _28572_ (.A1(_07865_),
    .A2(_09900_),
    .B(_09917_),
    .Y(_03097_));
 NOR2x1_ASAP7_75t_R _28573_ (.A(_00330_),
    .B(_09900_),
    .Y(_09918_));
 AO21x1_ASAP7_75t_R _28574_ (.A1(_07908_),
    .A2(_09900_),
    .B(_09918_),
    .Y(_03098_));
 NOR2x1_ASAP7_75t_R _28575_ (.A(_00693_),
    .B(_09900_),
    .Y(_09919_));
 AO21x1_ASAP7_75t_R _28576_ (.A1(_07950_),
    .A2(_09900_),
    .B(_09919_),
    .Y(_03099_));
 NOR2x1_ASAP7_75t_R _28577_ (.A(_00725_),
    .B(_09900_),
    .Y(_09920_));
 AO21x1_ASAP7_75t_R _28578_ (.A1(_07990_),
    .A2(_09900_),
    .B(_09920_),
    .Y(_03100_));
 NOR2x1_ASAP7_75t_R _28579_ (.A(_00758_),
    .B(_09900_),
    .Y(_09921_));
 AO21x1_ASAP7_75t_R _28580_ (.A1(_08034_),
    .A2(_09900_),
    .B(_09921_),
    .Y(_03101_));
 NOR2x1_ASAP7_75t_R _28581_ (.A(_00791_),
    .B(_09900_),
    .Y(_09922_));
 AO21x1_ASAP7_75t_R _28582_ (.A1(_08073_),
    .A2(_09900_),
    .B(_09922_),
    .Y(_03102_));
 NOR2x1_ASAP7_75t_R _28583_ (.A(_00824_),
    .B(_09900_),
    .Y(_09923_));
 AO21x1_ASAP7_75t_R _28584_ (.A1(_08116_),
    .A2(_09900_),
    .B(_09923_),
    .Y(_03103_));
 TAPCELL_ASAP7_75t_R PHY_513 ();
 NOR2x1_ASAP7_75t_R _28586_ (.A(_00856_),
    .B(_09900_),
    .Y(_09925_));
 AO21x1_ASAP7_75t_R _28587_ (.A1(_08150_),
    .A2(_09900_),
    .B(_09925_),
    .Y(_03104_));
 NOR2x1_ASAP7_75t_R _28588_ (.A(_00889_),
    .B(_09900_),
    .Y(_09926_));
 AO21x1_ASAP7_75t_R _28589_ (.A1(_08187_),
    .A2(_09900_),
    .B(_09926_),
    .Y(_03105_));
 TAPCELL_ASAP7_75t_R PHY_512 ();
 NOR2x1_ASAP7_75t_R _28591_ (.A(_00921_),
    .B(_09900_),
    .Y(_09928_));
 AO21x1_ASAP7_75t_R _28592_ (.A1(_08219_),
    .A2(_09900_),
    .B(_09928_),
    .Y(_03106_));
 NOR2x1_ASAP7_75t_R _28593_ (.A(_00954_),
    .B(_09900_),
    .Y(_09929_));
 AO21x1_ASAP7_75t_R _28594_ (.A1(_08254_),
    .A2(_09900_),
    .B(_09929_),
    .Y(_03107_));
 NOR2x1_ASAP7_75t_R _28595_ (.A(_00986_),
    .B(_09900_),
    .Y(_09930_));
 AO21x1_ASAP7_75t_R _28596_ (.A1(net250),
    .A2(_09900_),
    .B(_09930_),
    .Y(_03108_));
 NOR2x1_ASAP7_75t_R _28597_ (.A(_01020_),
    .B(_09900_),
    .Y(_09931_));
 AO21x1_ASAP7_75t_R _28598_ (.A1(_08319_),
    .A2(_09900_),
    .B(_09931_),
    .Y(_03109_));
 NOR2x1_ASAP7_75t_R _28599_ (.A(_01052_),
    .B(_09900_),
    .Y(_09932_));
 AO21x1_ASAP7_75t_R _28600_ (.A1(_08357_),
    .A2(_09900_),
    .B(_09932_),
    .Y(_03110_));
 NOR2x1_ASAP7_75t_R _28601_ (.A(_01085_),
    .B(_09900_),
    .Y(_09933_));
 AO21x1_ASAP7_75t_R _28602_ (.A1(_08388_),
    .A2(_09900_),
    .B(_09933_),
    .Y(_03111_));
 NOR2x1_ASAP7_75t_R _28603_ (.A(_01117_),
    .B(_09900_),
    .Y(_09934_));
 AO21x1_ASAP7_75t_R _28604_ (.A1(_08419_),
    .A2(_09900_),
    .B(_09934_),
    .Y(_03112_));
 NOR2x1_ASAP7_75t_R _28605_ (.A(_01151_),
    .B(_09900_),
    .Y(_09935_));
 AO21x1_ASAP7_75t_R _28606_ (.A1(_08451_),
    .A2(_09900_),
    .B(_09935_),
    .Y(_03113_));
 NOR2x1_ASAP7_75t_R _28607_ (.A(_01183_),
    .B(_09900_),
    .Y(_09936_));
 AO21x1_ASAP7_75t_R _28608_ (.A1(_08481_),
    .A2(_09900_),
    .B(_09936_),
    .Y(_03114_));
 NOR2x1_ASAP7_75t_R _28609_ (.A(_01217_),
    .B(_09900_),
    .Y(_09937_));
 AO21x1_ASAP7_75t_R _28610_ (.A1(_08512_),
    .A2(_09900_),
    .B(_09937_),
    .Y(_03115_));
 NOR2x1_ASAP7_75t_R _28611_ (.A(_01249_),
    .B(_09900_),
    .Y(_09938_));
 AO21x1_ASAP7_75t_R _28612_ (.A1(_08545_),
    .A2(_09900_),
    .B(_09938_),
    .Y(_03116_));
 NOR2x1_ASAP7_75t_R _28613_ (.A(_01283_),
    .B(_09900_),
    .Y(_09939_));
 AO21x1_ASAP7_75t_R _28614_ (.A1(_08573_),
    .A2(_09900_),
    .B(_09939_),
    .Y(_03117_));
 AND2x6_ASAP7_75t_R _28615_ (.A(_00187_),
    .B(_14021_),
    .Y(_09940_));
 AND4x2_ASAP7_75t_R _28616_ (.A(_00323_),
    .B(_00184_),
    .C(_09778_),
    .D(_09940_),
    .Y(_09941_));
 TAPCELL_ASAP7_75t_R PHY_511 ();
 TAPCELL_ASAP7_75t_R PHY_510 ();
 TAPCELL_ASAP7_75t_R PHY_509 ();
 NOR2x1_ASAP7_75t_R _28620_ (.A(_00299_),
    .B(net268),
    .Y(_09945_));
 AO21x1_ASAP7_75t_R _28621_ (.A1(_07180_),
    .A2(net268),
    .B(_09945_),
    .Y(_03118_));
 NOR2x1_ASAP7_75t_R _28622_ (.A(_00253_),
    .B(net268),
    .Y(_09946_));
 AO21x1_ASAP7_75t_R _28623_ (.A1(_07313_),
    .A2(net268),
    .B(_09946_),
    .Y(_03119_));
 NOR2x1_ASAP7_75t_R _28624_ (.A(_00361_),
    .B(_09941_),
    .Y(_09947_));
 AO21x1_ASAP7_75t_R _28625_ (.A1(_07398_),
    .A2(_09941_),
    .B(_09947_),
    .Y(_03120_));
 NOR2x1_ASAP7_75t_R _28626_ (.A(_00392_),
    .B(net268),
    .Y(_09948_));
 AO21x1_ASAP7_75t_R _28627_ (.A1(_07469_),
    .A2(net268),
    .B(_09948_),
    .Y(_03121_));
 NOR2x1_ASAP7_75t_R _28628_ (.A(_00422_),
    .B(net268),
    .Y(_09949_));
 AO21x1_ASAP7_75t_R _28629_ (.A1(_07534_),
    .A2(net268),
    .B(_09949_),
    .Y(_03122_));
 NOR2x1_ASAP7_75t_R _28630_ (.A(_00452_),
    .B(_09941_),
    .Y(_09950_));
 AO21x1_ASAP7_75t_R _28631_ (.A1(_07581_),
    .A2(_09941_),
    .B(_09950_),
    .Y(_03123_));
 NOR2x1_ASAP7_75t_R _28632_ (.A(_00482_),
    .B(net268),
    .Y(_09951_));
 AO21x1_ASAP7_75t_R _28633_ (.A1(net253),
    .A2(net268),
    .B(_09951_),
    .Y(_03124_));
 NOR2x1_ASAP7_75t_R _28634_ (.A(_00512_),
    .B(_09941_),
    .Y(_09952_));
 AO21x1_ASAP7_75t_R _28635_ (.A1(_07676_),
    .A2(_09941_),
    .B(_09952_),
    .Y(_03125_));
 TAPCELL_ASAP7_75t_R PHY_508 ();
 NOR2x1_ASAP7_75t_R _28637_ (.A(_00542_),
    .B(net268),
    .Y(_09954_));
 AO21x1_ASAP7_75t_R _28638_ (.A1(net252),
    .A2(net268),
    .B(_09954_),
    .Y(_03126_));
 NOR2x1_ASAP7_75t_R _28639_ (.A(_00572_),
    .B(net268),
    .Y(_09955_));
 AO21x1_ASAP7_75t_R _28640_ (.A1(_07780_),
    .A2(net268),
    .B(_09955_),
    .Y(_03127_));
 TAPCELL_ASAP7_75t_R PHY_507 ();
 NOR2x1_ASAP7_75t_R _28642_ (.A(_00602_),
    .B(_09941_),
    .Y(_09957_));
 AO21x1_ASAP7_75t_R _28643_ (.A1(_07817_),
    .A2(_09941_),
    .B(_09957_),
    .Y(_03128_));
 NOR2x1_ASAP7_75t_R _28644_ (.A(_00632_),
    .B(net268),
    .Y(_09958_));
 AO21x1_ASAP7_75t_R _28645_ (.A1(_07865_),
    .A2(net268),
    .B(_09958_),
    .Y(_03129_));
 NOR2x1_ASAP7_75t_R _28646_ (.A(_00331_),
    .B(net268),
    .Y(_09959_));
 AO21x1_ASAP7_75t_R _28647_ (.A1(_07908_),
    .A2(net268),
    .B(_09959_),
    .Y(_03130_));
 NOR2x1_ASAP7_75t_R _28648_ (.A(_00694_),
    .B(net267),
    .Y(_09960_));
 AO21x1_ASAP7_75t_R _28649_ (.A1(_07950_),
    .A2(net267),
    .B(_09960_),
    .Y(_03131_));
 NOR2x1_ASAP7_75t_R _28650_ (.A(_00726_),
    .B(net268),
    .Y(_09961_));
 AO21x1_ASAP7_75t_R _28651_ (.A1(_07990_),
    .A2(net268),
    .B(_09961_),
    .Y(_03132_));
 NOR2x1_ASAP7_75t_R _28652_ (.A(_00759_),
    .B(_09941_),
    .Y(_09962_));
 AO21x1_ASAP7_75t_R _28653_ (.A1(_08034_),
    .A2(_09941_),
    .B(_09962_),
    .Y(_03133_));
 NOR2x1_ASAP7_75t_R _28654_ (.A(_00792_),
    .B(net267),
    .Y(_09963_));
 AO21x1_ASAP7_75t_R _28655_ (.A1(_08073_),
    .A2(net267),
    .B(_09963_),
    .Y(_03134_));
 NOR2x1_ASAP7_75t_R _28656_ (.A(_00825_),
    .B(_09941_),
    .Y(_09964_));
 AO21x1_ASAP7_75t_R _28657_ (.A1(_08116_),
    .A2(_09941_),
    .B(_09964_),
    .Y(_03135_));
 TAPCELL_ASAP7_75t_R PHY_506 ();
 NOR2x1_ASAP7_75t_R _28659_ (.A(_00857_),
    .B(net267),
    .Y(_09966_));
 AO21x1_ASAP7_75t_R _28660_ (.A1(_08150_),
    .A2(net267),
    .B(_09966_),
    .Y(_03136_));
 NOR2x1_ASAP7_75t_R _28661_ (.A(_00890_),
    .B(net267),
    .Y(_09967_));
 AO21x1_ASAP7_75t_R _28662_ (.A1(_08187_),
    .A2(net267),
    .B(_09967_),
    .Y(_03137_));
 TAPCELL_ASAP7_75t_R PHY_505 ();
 NOR2x1_ASAP7_75t_R _28664_ (.A(_00922_),
    .B(_09941_),
    .Y(_09969_));
 AO21x1_ASAP7_75t_R _28665_ (.A1(_08219_),
    .A2(_09941_),
    .B(_09969_),
    .Y(_03138_));
 NOR2x1_ASAP7_75t_R _28666_ (.A(_00955_),
    .B(net267),
    .Y(_09970_));
 AO21x1_ASAP7_75t_R _28667_ (.A1(_08254_),
    .A2(net267),
    .B(_09970_),
    .Y(_03139_));
 NOR2x1_ASAP7_75t_R _28668_ (.A(_00987_),
    .B(net268),
    .Y(_09971_));
 AO21x1_ASAP7_75t_R _28669_ (.A1(net250),
    .A2(net268),
    .B(_09971_),
    .Y(_03140_));
 NOR2x1_ASAP7_75t_R _28670_ (.A(_01021_),
    .B(net267),
    .Y(_09972_));
 AO21x1_ASAP7_75t_R _28671_ (.A1(_08319_),
    .A2(net267),
    .B(_09972_),
    .Y(_03141_));
 NOR2x1_ASAP7_75t_R _28672_ (.A(_01053_),
    .B(net267),
    .Y(_09973_));
 AO21x1_ASAP7_75t_R _28673_ (.A1(_08357_),
    .A2(net267),
    .B(_09973_),
    .Y(_03142_));
 NOR2x1_ASAP7_75t_R _28674_ (.A(_01086_),
    .B(_09941_),
    .Y(_09974_));
 AO21x1_ASAP7_75t_R _28675_ (.A1(_08388_),
    .A2(_09941_),
    .B(_09974_),
    .Y(_03143_));
 NOR2x1_ASAP7_75t_R _28676_ (.A(_01118_),
    .B(net267),
    .Y(_09975_));
 AO21x1_ASAP7_75t_R _28677_ (.A1(_08419_),
    .A2(net267),
    .B(_09975_),
    .Y(_03144_));
 NOR2x1_ASAP7_75t_R _28678_ (.A(_01152_),
    .B(net267),
    .Y(_09976_));
 AO21x1_ASAP7_75t_R _28679_ (.A1(_08451_),
    .A2(net267),
    .B(_09976_),
    .Y(_03145_));
 NOR2x1_ASAP7_75t_R _28680_ (.A(_01184_),
    .B(_09941_),
    .Y(_09977_));
 AO21x1_ASAP7_75t_R _28681_ (.A1(_08481_),
    .A2(_09941_),
    .B(_09977_),
    .Y(_03146_));
 NOR2x1_ASAP7_75t_R _28682_ (.A(_01218_),
    .B(net267),
    .Y(_09978_));
 AO21x1_ASAP7_75t_R _28683_ (.A1(_08512_),
    .A2(net267),
    .B(_09978_),
    .Y(_03147_));
 NOR2x1_ASAP7_75t_R _28684_ (.A(_01250_),
    .B(_09941_),
    .Y(_09979_));
 AO21x1_ASAP7_75t_R _28685_ (.A1(_08545_),
    .A2(_09941_),
    .B(_09979_),
    .Y(_03148_));
 NOR2x1_ASAP7_75t_R _28686_ (.A(_01284_),
    .B(net268),
    .Y(_09980_));
 AO21x1_ASAP7_75t_R _28687_ (.A1(_08573_),
    .A2(net268),
    .B(_09980_),
    .Y(_03149_));
 AND2x6_ASAP7_75t_R _28688_ (.A(_06923_),
    .B(_09940_),
    .Y(_09981_));
 TAPCELL_ASAP7_75t_R PHY_504 ();
 TAPCELL_ASAP7_75t_R PHY_503 ();
 TAPCELL_ASAP7_75t_R PHY_502 ();
 NOR2x1_ASAP7_75t_R _28692_ (.A(_00300_),
    .B(_09981_),
    .Y(_09985_));
 AO21x1_ASAP7_75t_R _28693_ (.A1(_07180_),
    .A2(_09981_),
    .B(_09985_),
    .Y(_03150_));
 NOR2x1_ASAP7_75t_R _28694_ (.A(_00254_),
    .B(_09981_),
    .Y(_09986_));
 AO21x1_ASAP7_75t_R _28695_ (.A1(_07313_),
    .A2(_09981_),
    .B(_09986_),
    .Y(_03151_));
 NOR2x1_ASAP7_75t_R _28696_ (.A(_00362_),
    .B(_09981_),
    .Y(_09987_));
 AO21x1_ASAP7_75t_R _28697_ (.A1(_07398_),
    .A2(_09981_),
    .B(_09987_),
    .Y(_03152_));
 NOR2x1_ASAP7_75t_R _28698_ (.A(_00393_),
    .B(_09981_),
    .Y(_09988_));
 AO21x1_ASAP7_75t_R _28699_ (.A1(_07469_),
    .A2(_09981_),
    .B(_09988_),
    .Y(_03153_));
 NOR2x1_ASAP7_75t_R _28700_ (.A(_00423_),
    .B(_09981_),
    .Y(_09989_));
 AO21x1_ASAP7_75t_R _28701_ (.A1(_07534_),
    .A2(_09981_),
    .B(_09989_),
    .Y(_03154_));
 NOR2x1_ASAP7_75t_R _28702_ (.A(_00453_),
    .B(_09981_),
    .Y(_09990_));
 AO21x1_ASAP7_75t_R _28703_ (.A1(_07581_),
    .A2(_09981_),
    .B(_09990_),
    .Y(_03155_));
 NOR2x1_ASAP7_75t_R _28704_ (.A(_00483_),
    .B(_09981_),
    .Y(_09991_));
 AO21x1_ASAP7_75t_R _28705_ (.A1(net253),
    .A2(_09981_),
    .B(_09991_),
    .Y(_03156_));
 NOR2x1_ASAP7_75t_R _28706_ (.A(_00513_),
    .B(_09981_),
    .Y(_09992_));
 AO21x1_ASAP7_75t_R _28707_ (.A1(_07676_),
    .A2(_09981_),
    .B(_09992_),
    .Y(_03157_));
 TAPCELL_ASAP7_75t_R PHY_501 ();
 NOR2x1_ASAP7_75t_R _28709_ (.A(_00543_),
    .B(_09981_),
    .Y(_09994_));
 AO21x1_ASAP7_75t_R _28710_ (.A1(net252),
    .A2(_09981_),
    .B(_09994_),
    .Y(_03158_));
 NOR2x1_ASAP7_75t_R _28711_ (.A(_00573_),
    .B(_09981_),
    .Y(_09995_));
 AO21x1_ASAP7_75t_R _28712_ (.A1(_07780_),
    .A2(_09981_),
    .B(_09995_),
    .Y(_03159_));
 TAPCELL_ASAP7_75t_R PHY_500 ();
 NOR2x1_ASAP7_75t_R _28714_ (.A(_00603_),
    .B(_09981_),
    .Y(_09997_));
 AO21x1_ASAP7_75t_R _28715_ (.A1(_07817_),
    .A2(_09981_),
    .B(_09997_),
    .Y(_03160_));
 NOR2x1_ASAP7_75t_R _28716_ (.A(_00633_),
    .B(_09981_),
    .Y(_09998_));
 AO21x1_ASAP7_75t_R _28717_ (.A1(_07865_),
    .A2(_09981_),
    .B(_09998_),
    .Y(_03161_));
 NOR2x1_ASAP7_75t_R _28718_ (.A(_00332_),
    .B(_09981_),
    .Y(_09999_));
 AO21x1_ASAP7_75t_R _28719_ (.A1(_07908_),
    .A2(_09981_),
    .B(_09999_),
    .Y(_03162_));
 NOR2x1_ASAP7_75t_R _28720_ (.A(_00695_),
    .B(_09981_),
    .Y(_10000_));
 AO21x1_ASAP7_75t_R _28721_ (.A1(_07950_),
    .A2(_09981_),
    .B(_10000_),
    .Y(_03163_));
 NOR2x1_ASAP7_75t_R _28722_ (.A(_00727_),
    .B(_09981_),
    .Y(_10001_));
 AO21x1_ASAP7_75t_R _28723_ (.A1(_07990_),
    .A2(_09981_),
    .B(_10001_),
    .Y(_03164_));
 NOR2x1_ASAP7_75t_R _28724_ (.A(_00760_),
    .B(_09981_),
    .Y(_10002_));
 AO21x1_ASAP7_75t_R _28725_ (.A1(_08034_),
    .A2(_09981_),
    .B(_10002_),
    .Y(_03165_));
 NOR2x1_ASAP7_75t_R _28726_ (.A(_00793_),
    .B(_09981_),
    .Y(_10003_));
 AO21x1_ASAP7_75t_R _28727_ (.A1(_08073_),
    .A2(_09981_),
    .B(_10003_),
    .Y(_03166_));
 NOR2x1_ASAP7_75t_R _28728_ (.A(_00826_),
    .B(_09981_),
    .Y(_10004_));
 AO21x1_ASAP7_75t_R _28729_ (.A1(_08116_),
    .A2(_09981_),
    .B(_10004_),
    .Y(_03167_));
 TAPCELL_ASAP7_75t_R PHY_499 ();
 NOR2x1_ASAP7_75t_R _28731_ (.A(_00858_),
    .B(_09981_),
    .Y(_10006_));
 AO21x1_ASAP7_75t_R _28732_ (.A1(_08150_),
    .A2(_09981_),
    .B(_10006_),
    .Y(_03168_));
 NOR2x1_ASAP7_75t_R _28733_ (.A(_00891_),
    .B(_09981_),
    .Y(_10007_));
 AO21x1_ASAP7_75t_R _28734_ (.A1(_08187_),
    .A2(_09981_),
    .B(_10007_),
    .Y(_03169_));
 TAPCELL_ASAP7_75t_R PHY_498 ();
 NOR2x1_ASAP7_75t_R _28736_ (.A(_00923_),
    .B(_09981_),
    .Y(_10009_));
 AO21x1_ASAP7_75t_R _28737_ (.A1(_08219_),
    .A2(_09981_),
    .B(_10009_),
    .Y(_03170_));
 NOR2x1_ASAP7_75t_R _28738_ (.A(_00956_),
    .B(_09981_),
    .Y(_10010_));
 AO21x1_ASAP7_75t_R _28739_ (.A1(_08254_),
    .A2(_09981_),
    .B(_10010_),
    .Y(_03171_));
 NOR2x1_ASAP7_75t_R _28740_ (.A(_00988_),
    .B(_09981_),
    .Y(_10011_));
 AO21x1_ASAP7_75t_R _28741_ (.A1(net250),
    .A2(_09981_),
    .B(_10011_),
    .Y(_03172_));
 NOR2x1_ASAP7_75t_R _28742_ (.A(_01022_),
    .B(_09981_),
    .Y(_10012_));
 AO21x1_ASAP7_75t_R _28743_ (.A1(_08319_),
    .A2(_09981_),
    .B(_10012_),
    .Y(_03173_));
 NOR2x1_ASAP7_75t_R _28744_ (.A(_01054_),
    .B(_09981_),
    .Y(_10013_));
 AO21x1_ASAP7_75t_R _28745_ (.A1(_08357_),
    .A2(_09981_),
    .B(_10013_),
    .Y(_03174_));
 NOR2x1_ASAP7_75t_R _28746_ (.A(_01087_),
    .B(_09981_),
    .Y(_10014_));
 AO21x1_ASAP7_75t_R _28747_ (.A1(_08388_),
    .A2(_09981_),
    .B(_10014_),
    .Y(_03175_));
 NOR2x1_ASAP7_75t_R _28748_ (.A(_01119_),
    .B(_09981_),
    .Y(_10015_));
 AO21x1_ASAP7_75t_R _28749_ (.A1(_08419_),
    .A2(_09981_),
    .B(_10015_),
    .Y(_03176_));
 NOR2x1_ASAP7_75t_R _28750_ (.A(_01153_),
    .B(_09981_),
    .Y(_10016_));
 AO21x1_ASAP7_75t_R _28751_ (.A1(_08451_),
    .A2(_09981_),
    .B(_10016_),
    .Y(_03177_));
 NOR2x1_ASAP7_75t_R _28752_ (.A(_01185_),
    .B(_09981_),
    .Y(_10017_));
 AO21x1_ASAP7_75t_R _28753_ (.A1(_08481_),
    .A2(_09981_),
    .B(_10017_),
    .Y(_03178_));
 NOR2x1_ASAP7_75t_R _28754_ (.A(_01219_),
    .B(_09981_),
    .Y(_10018_));
 AO21x1_ASAP7_75t_R _28755_ (.A1(_08512_),
    .A2(_09981_),
    .B(_10018_),
    .Y(_03179_));
 NOR2x1_ASAP7_75t_R _28756_ (.A(_01251_),
    .B(_09981_),
    .Y(_10019_));
 AO21x1_ASAP7_75t_R _28757_ (.A1(_08545_),
    .A2(_09981_),
    .B(_10019_),
    .Y(_03180_));
 NOR2x1_ASAP7_75t_R _28758_ (.A(_01285_),
    .B(_09981_),
    .Y(_10020_));
 AO21x1_ASAP7_75t_R _28759_ (.A1(_08573_),
    .A2(_09981_),
    .B(_10020_),
    .Y(_03181_));
 AND2x6_ASAP7_75t_R _28760_ (.A(_09664_),
    .B(_09940_),
    .Y(_10021_));
 TAPCELL_ASAP7_75t_R PHY_497 ();
 TAPCELL_ASAP7_75t_R PHY_496 ();
 TAPCELL_ASAP7_75t_R PHY_495 ();
 NOR2x1_ASAP7_75t_R _28764_ (.A(_00301_),
    .B(_10021_),
    .Y(_10025_));
 AO21x1_ASAP7_75t_R _28765_ (.A1(_07180_),
    .A2(_10021_),
    .B(_10025_),
    .Y(_03182_));
 NOR2x1_ASAP7_75t_R _28766_ (.A(_00255_),
    .B(_10021_),
    .Y(_10026_));
 AO21x1_ASAP7_75t_R _28767_ (.A1(_07313_),
    .A2(_10021_),
    .B(_10026_),
    .Y(_03183_));
 NOR2x1_ASAP7_75t_R _28768_ (.A(_00363_),
    .B(_10021_),
    .Y(_10027_));
 AO21x1_ASAP7_75t_R _28769_ (.A1(_07398_),
    .A2(_10021_),
    .B(_10027_),
    .Y(_03184_));
 NOR2x1_ASAP7_75t_R _28770_ (.A(_00394_),
    .B(_10021_),
    .Y(_10028_));
 AO21x1_ASAP7_75t_R _28771_ (.A1(_07469_),
    .A2(_10021_),
    .B(_10028_),
    .Y(_03185_));
 NOR2x1_ASAP7_75t_R _28772_ (.A(_00424_),
    .B(_10021_),
    .Y(_10029_));
 AO21x1_ASAP7_75t_R _28773_ (.A1(_07534_),
    .A2(_10021_),
    .B(_10029_),
    .Y(_03186_));
 NOR2x1_ASAP7_75t_R _28774_ (.A(_00454_),
    .B(_10021_),
    .Y(_10030_));
 AO21x1_ASAP7_75t_R _28775_ (.A1(_07581_),
    .A2(_10021_),
    .B(_10030_),
    .Y(_03187_));
 NOR2x1_ASAP7_75t_R _28776_ (.A(_00484_),
    .B(_10021_),
    .Y(_10031_));
 AO21x1_ASAP7_75t_R _28777_ (.A1(net253),
    .A2(_10021_),
    .B(_10031_),
    .Y(_03188_));
 NOR2x1_ASAP7_75t_R _28778_ (.A(_00514_),
    .B(_10021_),
    .Y(_10032_));
 AO21x1_ASAP7_75t_R _28779_ (.A1(_07676_),
    .A2(_10021_),
    .B(_10032_),
    .Y(_03189_));
 TAPCELL_ASAP7_75t_R PHY_494 ();
 NOR2x1_ASAP7_75t_R _28781_ (.A(_00544_),
    .B(_10021_),
    .Y(_10034_));
 AO21x1_ASAP7_75t_R _28782_ (.A1(net252),
    .A2(_10021_),
    .B(_10034_),
    .Y(_03190_));
 NOR2x1_ASAP7_75t_R _28783_ (.A(_00574_),
    .B(_10021_),
    .Y(_10035_));
 AO21x1_ASAP7_75t_R _28784_ (.A1(_07780_),
    .A2(_10021_),
    .B(_10035_),
    .Y(_03191_));
 TAPCELL_ASAP7_75t_R PHY_493 ();
 NOR2x1_ASAP7_75t_R _28786_ (.A(_00604_),
    .B(_10021_),
    .Y(_10037_));
 AO21x1_ASAP7_75t_R _28787_ (.A1(_07817_),
    .A2(_10021_),
    .B(_10037_),
    .Y(_03192_));
 NOR2x1_ASAP7_75t_R _28788_ (.A(_00634_),
    .B(_10021_),
    .Y(_10038_));
 AO21x1_ASAP7_75t_R _28789_ (.A1(_07865_),
    .A2(_10021_),
    .B(_10038_),
    .Y(_03193_));
 NOR2x1_ASAP7_75t_R _28790_ (.A(_00333_),
    .B(_10021_),
    .Y(_10039_));
 AO21x1_ASAP7_75t_R _28791_ (.A1(_07908_),
    .A2(_10021_),
    .B(_10039_),
    .Y(_03194_));
 NOR2x1_ASAP7_75t_R _28792_ (.A(_00696_),
    .B(_10021_),
    .Y(_10040_));
 AO21x1_ASAP7_75t_R _28793_ (.A1(_07950_),
    .A2(_10021_),
    .B(_10040_),
    .Y(_03195_));
 NOR2x1_ASAP7_75t_R _28794_ (.A(_00728_),
    .B(_10021_),
    .Y(_10041_));
 AO21x1_ASAP7_75t_R _28795_ (.A1(_07990_),
    .A2(_10021_),
    .B(_10041_),
    .Y(_03196_));
 NOR2x1_ASAP7_75t_R _28796_ (.A(_00761_),
    .B(_10021_),
    .Y(_10042_));
 AO21x1_ASAP7_75t_R _28797_ (.A1(_08034_),
    .A2(_10021_),
    .B(_10042_),
    .Y(_03197_));
 NOR2x1_ASAP7_75t_R _28798_ (.A(_00794_),
    .B(_10021_),
    .Y(_10043_));
 AO21x1_ASAP7_75t_R _28799_ (.A1(_08073_),
    .A2(_10021_),
    .B(_10043_),
    .Y(_03198_));
 NOR2x1_ASAP7_75t_R _28800_ (.A(_00827_),
    .B(_10021_),
    .Y(_10044_));
 AO21x1_ASAP7_75t_R _28801_ (.A1(_08116_),
    .A2(_10021_),
    .B(_10044_),
    .Y(_03199_));
 TAPCELL_ASAP7_75t_R PHY_492 ();
 NOR2x1_ASAP7_75t_R _28803_ (.A(_00859_),
    .B(_10021_),
    .Y(_10046_));
 AO21x1_ASAP7_75t_R _28804_ (.A1(_08150_),
    .A2(_10021_),
    .B(_10046_),
    .Y(_03200_));
 NOR2x1_ASAP7_75t_R _28805_ (.A(_00892_),
    .B(_10021_),
    .Y(_10047_));
 AO21x1_ASAP7_75t_R _28806_ (.A1(_08187_),
    .A2(_10021_),
    .B(_10047_),
    .Y(_03201_));
 TAPCELL_ASAP7_75t_R PHY_491 ();
 NOR2x1_ASAP7_75t_R _28808_ (.A(_00924_),
    .B(_10021_),
    .Y(_10049_));
 AO21x1_ASAP7_75t_R _28809_ (.A1(_08219_),
    .A2(_10021_),
    .B(_10049_),
    .Y(_03202_));
 NOR2x1_ASAP7_75t_R _28810_ (.A(_00957_),
    .B(_10021_),
    .Y(_10050_));
 AO21x1_ASAP7_75t_R _28811_ (.A1(_08254_),
    .A2(_10021_),
    .B(_10050_),
    .Y(_03203_));
 NOR2x1_ASAP7_75t_R _28812_ (.A(_00989_),
    .B(_10021_),
    .Y(_10051_));
 AO21x1_ASAP7_75t_R _28813_ (.A1(net250),
    .A2(_10021_),
    .B(_10051_),
    .Y(_03204_));
 NOR2x1_ASAP7_75t_R _28814_ (.A(_01023_),
    .B(_10021_),
    .Y(_10052_));
 AO21x1_ASAP7_75t_R _28815_ (.A1(_08319_),
    .A2(_10021_),
    .B(_10052_),
    .Y(_03205_));
 NOR2x1_ASAP7_75t_R _28816_ (.A(_01055_),
    .B(_10021_),
    .Y(_10053_));
 AO21x1_ASAP7_75t_R _28817_ (.A1(_08357_),
    .A2(_10021_),
    .B(_10053_),
    .Y(_03206_));
 NOR2x1_ASAP7_75t_R _28818_ (.A(_01088_),
    .B(_10021_),
    .Y(_10054_));
 AO21x1_ASAP7_75t_R _28819_ (.A1(_08388_),
    .A2(_10021_),
    .B(_10054_),
    .Y(_03207_));
 NOR2x1_ASAP7_75t_R _28820_ (.A(_01120_),
    .B(_10021_),
    .Y(_10055_));
 AO21x1_ASAP7_75t_R _28821_ (.A1(_08419_),
    .A2(_10021_),
    .B(_10055_),
    .Y(_03208_));
 NOR2x1_ASAP7_75t_R _28822_ (.A(_01154_),
    .B(_10021_),
    .Y(_10056_));
 AO21x1_ASAP7_75t_R _28823_ (.A1(_08451_),
    .A2(_10021_),
    .B(_10056_),
    .Y(_03209_));
 NOR2x1_ASAP7_75t_R _28824_ (.A(_01186_),
    .B(_10021_),
    .Y(_10057_));
 AO21x1_ASAP7_75t_R _28825_ (.A1(_08481_),
    .A2(_10021_),
    .B(_10057_),
    .Y(_03210_));
 NOR2x1_ASAP7_75t_R _28826_ (.A(_01220_),
    .B(_10021_),
    .Y(_10058_));
 AO21x1_ASAP7_75t_R _28827_ (.A1(_08512_),
    .A2(_10021_),
    .B(_10058_),
    .Y(_03211_));
 NOR2x1_ASAP7_75t_R _28828_ (.A(_01252_),
    .B(_10021_),
    .Y(_10059_));
 AO21x1_ASAP7_75t_R _28829_ (.A1(_08545_),
    .A2(_10021_),
    .B(_10059_),
    .Y(_03212_));
 NOR2x1_ASAP7_75t_R _28830_ (.A(_01286_),
    .B(_10021_),
    .Y(_10060_));
 AO21x1_ASAP7_75t_R _28831_ (.A1(_08573_),
    .A2(_10021_),
    .B(_10060_),
    .Y(_03213_));
 AND2x6_ASAP7_75t_R _28832_ (.A(_09737_),
    .B(_09940_),
    .Y(_10061_));
 TAPCELL_ASAP7_75t_R PHY_490 ();
 TAPCELL_ASAP7_75t_R PHY_489 ();
 TAPCELL_ASAP7_75t_R PHY_488 ();
 NOR2x1_ASAP7_75t_R _28836_ (.A(_00302_),
    .B(_10061_),
    .Y(_10065_));
 AO21x1_ASAP7_75t_R _28837_ (.A1(_07180_),
    .A2(_10061_),
    .B(_10065_),
    .Y(_03214_));
 NOR2x1_ASAP7_75t_R _28838_ (.A(_00256_),
    .B(_10061_),
    .Y(_10066_));
 AO21x1_ASAP7_75t_R _28839_ (.A1(_07313_),
    .A2(_10061_),
    .B(_10066_),
    .Y(_03215_));
 NOR2x1_ASAP7_75t_R _28840_ (.A(_00364_),
    .B(_10061_),
    .Y(_10067_));
 AO21x1_ASAP7_75t_R _28841_ (.A1(_07398_),
    .A2(_10061_),
    .B(_10067_),
    .Y(_03216_));
 NOR2x1_ASAP7_75t_R _28842_ (.A(_00395_),
    .B(_10061_),
    .Y(_10068_));
 AO21x1_ASAP7_75t_R _28843_ (.A1(_07469_),
    .A2(_10061_),
    .B(_10068_),
    .Y(_03217_));
 NOR2x1_ASAP7_75t_R _28844_ (.A(_00425_),
    .B(_10061_),
    .Y(_10069_));
 AO21x1_ASAP7_75t_R _28845_ (.A1(_07534_),
    .A2(_10061_),
    .B(_10069_),
    .Y(_03218_));
 NOR2x1_ASAP7_75t_R _28846_ (.A(_00455_),
    .B(_10061_),
    .Y(_10070_));
 AO21x1_ASAP7_75t_R _28847_ (.A1(_07581_),
    .A2(_10061_),
    .B(_10070_),
    .Y(_03219_));
 NOR2x1_ASAP7_75t_R _28848_ (.A(_00485_),
    .B(_10061_),
    .Y(_10071_));
 AO21x1_ASAP7_75t_R _28849_ (.A1(net253),
    .A2(_10061_),
    .B(_10071_),
    .Y(_03220_));
 NOR2x1_ASAP7_75t_R _28850_ (.A(_00515_),
    .B(_10061_),
    .Y(_10072_));
 AO21x1_ASAP7_75t_R _28851_ (.A1(_07676_),
    .A2(_10061_),
    .B(_10072_),
    .Y(_03221_));
 TAPCELL_ASAP7_75t_R PHY_487 ();
 NOR2x1_ASAP7_75t_R _28853_ (.A(_00545_),
    .B(_10061_),
    .Y(_10074_));
 AO21x1_ASAP7_75t_R _28854_ (.A1(net252),
    .A2(_10061_),
    .B(_10074_),
    .Y(_03222_));
 NOR2x1_ASAP7_75t_R _28855_ (.A(_00575_),
    .B(_10061_),
    .Y(_10075_));
 AO21x1_ASAP7_75t_R _28856_ (.A1(_07780_),
    .A2(_10061_),
    .B(_10075_),
    .Y(_03223_));
 TAPCELL_ASAP7_75t_R PHY_486 ();
 NOR2x1_ASAP7_75t_R _28858_ (.A(_00605_),
    .B(_10061_),
    .Y(_10077_));
 AO21x1_ASAP7_75t_R _28859_ (.A1(_07817_),
    .A2(_10061_),
    .B(_10077_),
    .Y(_03224_));
 NOR2x1_ASAP7_75t_R _28860_ (.A(_00635_),
    .B(_10061_),
    .Y(_10078_));
 AO21x1_ASAP7_75t_R _28861_ (.A1(_07865_),
    .A2(_10061_),
    .B(_10078_),
    .Y(_03225_));
 NOR2x1_ASAP7_75t_R _28862_ (.A(_00334_),
    .B(_10061_),
    .Y(_10079_));
 AO21x1_ASAP7_75t_R _28863_ (.A1(_07908_),
    .A2(_10061_),
    .B(_10079_),
    .Y(_03226_));
 NOR2x1_ASAP7_75t_R _28864_ (.A(_00697_),
    .B(_10061_),
    .Y(_10080_));
 AO21x1_ASAP7_75t_R _28865_ (.A1(_07950_),
    .A2(_10061_),
    .B(_10080_),
    .Y(_03227_));
 NOR2x1_ASAP7_75t_R _28866_ (.A(_00729_),
    .B(_10061_),
    .Y(_10081_));
 AO21x1_ASAP7_75t_R _28867_ (.A1(_07990_),
    .A2(_10061_),
    .B(_10081_),
    .Y(_03228_));
 NOR2x1_ASAP7_75t_R _28868_ (.A(_00762_),
    .B(_10061_),
    .Y(_10082_));
 AO21x1_ASAP7_75t_R _28869_ (.A1(_08034_),
    .A2(_10061_),
    .B(_10082_),
    .Y(_03229_));
 NOR2x1_ASAP7_75t_R _28870_ (.A(_00795_),
    .B(_10061_),
    .Y(_10083_));
 AO21x1_ASAP7_75t_R _28871_ (.A1(_08073_),
    .A2(_10061_),
    .B(_10083_),
    .Y(_03230_));
 NOR2x1_ASAP7_75t_R _28872_ (.A(_00828_),
    .B(_10061_),
    .Y(_10084_));
 AO21x1_ASAP7_75t_R _28873_ (.A1(_08116_),
    .A2(_10061_),
    .B(_10084_),
    .Y(_03231_));
 TAPCELL_ASAP7_75t_R PHY_485 ();
 NOR2x1_ASAP7_75t_R _28875_ (.A(_00860_),
    .B(_10061_),
    .Y(_10086_));
 AO21x1_ASAP7_75t_R _28876_ (.A1(_08150_),
    .A2(_10061_),
    .B(_10086_),
    .Y(_03232_));
 NOR2x1_ASAP7_75t_R _28877_ (.A(_00893_),
    .B(_10061_),
    .Y(_10087_));
 AO21x1_ASAP7_75t_R _28878_ (.A1(_08187_),
    .A2(_10061_),
    .B(_10087_),
    .Y(_03233_));
 TAPCELL_ASAP7_75t_R PHY_484 ();
 NOR2x1_ASAP7_75t_R _28880_ (.A(_00925_),
    .B(_10061_),
    .Y(_10089_));
 AO21x1_ASAP7_75t_R _28881_ (.A1(_08219_),
    .A2(_10061_),
    .B(_10089_),
    .Y(_03234_));
 NOR2x1_ASAP7_75t_R _28882_ (.A(_00958_),
    .B(_10061_),
    .Y(_10090_));
 AO21x1_ASAP7_75t_R _28883_ (.A1(_08254_),
    .A2(_10061_),
    .B(_10090_),
    .Y(_03235_));
 NOR2x1_ASAP7_75t_R _28884_ (.A(_00990_),
    .B(_10061_),
    .Y(_10091_));
 AO21x1_ASAP7_75t_R _28885_ (.A1(net250),
    .A2(_10061_),
    .B(_10091_),
    .Y(_03236_));
 NOR2x1_ASAP7_75t_R _28886_ (.A(_01024_),
    .B(_10061_),
    .Y(_10092_));
 AO21x1_ASAP7_75t_R _28887_ (.A1(_08319_),
    .A2(_10061_),
    .B(_10092_),
    .Y(_03237_));
 NOR2x1_ASAP7_75t_R _28888_ (.A(_01056_),
    .B(_10061_),
    .Y(_10093_));
 AO21x1_ASAP7_75t_R _28889_ (.A1(_08357_),
    .A2(_10061_),
    .B(_10093_),
    .Y(_03238_));
 NOR2x1_ASAP7_75t_R _28890_ (.A(_01089_),
    .B(_10061_),
    .Y(_10094_));
 AO21x1_ASAP7_75t_R _28891_ (.A1(_08388_),
    .A2(_10061_),
    .B(_10094_),
    .Y(_03239_));
 NOR2x1_ASAP7_75t_R _28892_ (.A(_01121_),
    .B(_10061_),
    .Y(_10095_));
 AO21x1_ASAP7_75t_R _28893_ (.A1(_08419_),
    .A2(_10061_),
    .B(_10095_),
    .Y(_03240_));
 NOR2x1_ASAP7_75t_R _28894_ (.A(_01155_),
    .B(_10061_),
    .Y(_10096_));
 AO21x1_ASAP7_75t_R _28895_ (.A1(_08451_),
    .A2(_10061_),
    .B(_10096_),
    .Y(_03241_));
 NOR2x1_ASAP7_75t_R _28896_ (.A(_01187_),
    .B(_10061_),
    .Y(_10097_));
 AO21x1_ASAP7_75t_R _28897_ (.A1(_08481_),
    .A2(_10061_),
    .B(_10097_),
    .Y(_03242_));
 NOR2x1_ASAP7_75t_R _28898_ (.A(_01221_),
    .B(_10061_),
    .Y(_10098_));
 AO21x1_ASAP7_75t_R _28899_ (.A1(_08512_),
    .A2(_10061_),
    .B(_10098_),
    .Y(_03243_));
 NOR2x1_ASAP7_75t_R _28900_ (.A(_01253_),
    .B(_10061_),
    .Y(_10099_));
 AO21x1_ASAP7_75t_R _28901_ (.A1(_08545_),
    .A2(_10061_),
    .B(_10099_),
    .Y(_03244_));
 NOR2x1_ASAP7_75t_R _28902_ (.A(_01287_),
    .B(_10061_),
    .Y(_10100_));
 AO21x1_ASAP7_75t_R _28903_ (.A1(_08573_),
    .A2(_10061_),
    .B(_10100_),
    .Y(_03245_));
 TAPCELL_ASAP7_75t_R PHY_483 ();
 NOR2x2_ASAP7_75t_R _28905_ (.A(_00187_),
    .B(_00191_),
    .Y(_10102_));
 AND4x2_ASAP7_75t_R _28906_ (.A(_00323_),
    .B(_00184_),
    .C(_09778_),
    .D(_10102_),
    .Y(_10103_));
 TAPCELL_ASAP7_75t_R PHY_482 ();
 TAPCELL_ASAP7_75t_R PHY_481 ();
 TAPCELL_ASAP7_75t_R PHY_480 ();
 NOR2x1_ASAP7_75t_R _28910_ (.A(_00303_),
    .B(net265),
    .Y(_10107_));
 AO21x1_ASAP7_75t_R _28911_ (.A1(_07180_),
    .A2(net265),
    .B(_10107_),
    .Y(_03246_));
 TAPCELL_ASAP7_75t_R PHY_479 ();
 NOR2x1_ASAP7_75t_R _28913_ (.A(_00257_),
    .B(net265),
    .Y(_10109_));
 AO21x1_ASAP7_75t_R _28914_ (.A1(_07313_),
    .A2(net265),
    .B(_10109_),
    .Y(_03247_));
 TAPCELL_ASAP7_75t_R PHY_478 ();
 NOR2x1_ASAP7_75t_R _28916_ (.A(_00365_),
    .B(net265),
    .Y(_10111_));
 AO21x1_ASAP7_75t_R _28917_ (.A1(_07398_),
    .A2(net265),
    .B(_10111_),
    .Y(_03248_));
 TAPCELL_ASAP7_75t_R PHY_477 ();
 NOR2x1_ASAP7_75t_R _28919_ (.A(_00396_),
    .B(net265),
    .Y(_10113_));
 AO21x1_ASAP7_75t_R _28920_ (.A1(_07469_),
    .A2(net265),
    .B(_10113_),
    .Y(_03249_));
 TAPCELL_ASAP7_75t_R PHY_476 ();
 NOR2x1_ASAP7_75t_R _28922_ (.A(_00426_),
    .B(_10103_),
    .Y(_10115_));
 AO21x1_ASAP7_75t_R _28923_ (.A1(_07534_),
    .A2(_10103_),
    .B(_10115_),
    .Y(_03250_));
 TAPCELL_ASAP7_75t_R PHY_475 ();
 NOR2x1_ASAP7_75t_R _28925_ (.A(_00456_),
    .B(net264),
    .Y(_10117_));
 AO21x1_ASAP7_75t_R _28926_ (.A1(_07581_),
    .A2(net264),
    .B(_10117_),
    .Y(_03251_));
 TAPCELL_ASAP7_75t_R PHY_474 ();
 NOR2x1_ASAP7_75t_R _28928_ (.A(_00486_),
    .B(_10103_),
    .Y(_10119_));
 AO21x1_ASAP7_75t_R _28929_ (.A1(net253),
    .A2(_10103_),
    .B(_10119_),
    .Y(_03252_));
 TAPCELL_ASAP7_75t_R PHY_473 ();
 NOR2x1_ASAP7_75t_R _28931_ (.A(_00516_),
    .B(net265),
    .Y(_10121_));
 AO21x1_ASAP7_75t_R _28932_ (.A1(_07676_),
    .A2(net265),
    .B(_10121_),
    .Y(_03253_));
 TAPCELL_ASAP7_75t_R PHY_472 ();
 TAPCELL_ASAP7_75t_R PHY_471 ();
 NOR2x1_ASAP7_75t_R _28935_ (.A(_00546_),
    .B(net265),
    .Y(_10124_));
 AO21x1_ASAP7_75t_R _28936_ (.A1(net252),
    .A2(net265),
    .B(_10124_),
    .Y(_03254_));
 TAPCELL_ASAP7_75t_R PHY_470 ();
 NOR2x1_ASAP7_75t_R _28938_ (.A(_00576_),
    .B(_10103_),
    .Y(_10126_));
 AO21x1_ASAP7_75t_R _28939_ (.A1(_07780_),
    .A2(_10103_),
    .B(_10126_),
    .Y(_03255_));
 TAPCELL_ASAP7_75t_R PHY_469 ();
 TAPCELL_ASAP7_75t_R PHY_468 ();
 NOR2x1_ASAP7_75t_R _28942_ (.A(_00606_),
    .B(net264),
    .Y(_10129_));
 AO21x1_ASAP7_75t_R _28943_ (.A1(_07817_),
    .A2(net264),
    .B(_10129_),
    .Y(_03256_));
 TAPCELL_ASAP7_75t_R PHY_467 ();
 NOR2x1_ASAP7_75t_R _28945_ (.A(_00636_),
    .B(net265),
    .Y(_10131_));
 AO21x1_ASAP7_75t_R _28946_ (.A1(_07865_),
    .A2(net265),
    .B(_10131_),
    .Y(_03257_));
 TAPCELL_ASAP7_75t_R PHY_466 ();
 NOR2x1_ASAP7_75t_R _28948_ (.A(_00335_),
    .B(net265),
    .Y(_10133_));
 AO21x1_ASAP7_75t_R _28949_ (.A1(_07908_),
    .A2(net265),
    .B(_10133_),
    .Y(_03258_));
 TAPCELL_ASAP7_75t_R PHY_465 ();
 NOR2x1_ASAP7_75t_R _28951_ (.A(_00698_),
    .B(net264),
    .Y(_10135_));
 AO21x1_ASAP7_75t_R _28952_ (.A1(_07950_),
    .A2(net264),
    .B(_10135_),
    .Y(_03259_));
 TAPCELL_ASAP7_75t_R PHY_464 ();
 NOR2x1_ASAP7_75t_R _28954_ (.A(_00730_),
    .B(_10103_),
    .Y(_10137_));
 AO21x1_ASAP7_75t_R _28955_ (.A1(_07990_),
    .A2(_10103_),
    .B(_10137_),
    .Y(_03260_));
 TAPCELL_ASAP7_75t_R PHY_463 ();
 NOR2x1_ASAP7_75t_R _28957_ (.A(_00763_),
    .B(net264),
    .Y(_10139_));
 AO21x1_ASAP7_75t_R _28958_ (.A1(_08034_),
    .A2(net264),
    .B(_10139_),
    .Y(_03261_));
 TAPCELL_ASAP7_75t_R PHY_462 ();
 NOR2x1_ASAP7_75t_R _28960_ (.A(_00796_),
    .B(net264),
    .Y(_10141_));
 AO21x1_ASAP7_75t_R _28961_ (.A1(_08073_),
    .A2(net264),
    .B(_10141_),
    .Y(_03262_));
 TAPCELL_ASAP7_75t_R PHY_461 ();
 NOR2x1_ASAP7_75t_R _28963_ (.A(_00829_),
    .B(net264),
    .Y(_10143_));
 AO21x1_ASAP7_75t_R _28964_ (.A1(_08116_),
    .A2(net264),
    .B(_10143_),
    .Y(_03263_));
 TAPCELL_ASAP7_75t_R PHY_460 ();
 TAPCELL_ASAP7_75t_R PHY_459 ();
 NOR2x1_ASAP7_75t_R _28967_ (.A(_00861_),
    .B(net266),
    .Y(_10146_));
 AO21x1_ASAP7_75t_R _28968_ (.A1(net251),
    .A2(net266),
    .B(_10146_),
    .Y(_03264_));
 TAPCELL_ASAP7_75t_R PHY_458 ();
 NOR2x1_ASAP7_75t_R _28970_ (.A(_00894_),
    .B(net266),
    .Y(_10148_));
 AO21x1_ASAP7_75t_R _28971_ (.A1(_08187_),
    .A2(net266),
    .B(_10148_),
    .Y(_03265_));
 TAPCELL_ASAP7_75t_R PHY_457 ();
 TAPCELL_ASAP7_75t_R PHY_456 ();
 NOR2x1_ASAP7_75t_R _28974_ (.A(_00926_),
    .B(net264),
    .Y(_10151_));
 AO21x1_ASAP7_75t_R _28975_ (.A1(_08219_),
    .A2(net264),
    .B(_10151_),
    .Y(_03266_));
 TAPCELL_ASAP7_75t_R PHY_455 ();
 NOR2x1_ASAP7_75t_R _28977_ (.A(_00959_),
    .B(net266),
    .Y(_10153_));
 AO21x1_ASAP7_75t_R _28978_ (.A1(_08254_),
    .A2(net266),
    .B(_10153_),
    .Y(_03267_));
 TAPCELL_ASAP7_75t_R PHY_454 ();
 NOR2x1_ASAP7_75t_R _28980_ (.A(_00991_),
    .B(_10103_),
    .Y(_10155_));
 AO21x1_ASAP7_75t_R _28981_ (.A1(net250),
    .A2(_10103_),
    .B(_10155_),
    .Y(_03268_));
 TAPCELL_ASAP7_75t_R PHY_453 ();
 NOR2x1_ASAP7_75t_R _28983_ (.A(_01025_),
    .B(net266),
    .Y(_10157_));
 AO21x1_ASAP7_75t_R _28984_ (.A1(_08319_),
    .A2(net266),
    .B(_10157_),
    .Y(_03269_));
 TAPCELL_ASAP7_75t_R PHY_452 ();
 NOR2x1_ASAP7_75t_R _28986_ (.A(_01057_),
    .B(net264),
    .Y(_10159_));
 AO21x1_ASAP7_75t_R _28987_ (.A1(_08357_),
    .A2(net264),
    .B(_10159_),
    .Y(_03270_));
 TAPCELL_ASAP7_75t_R PHY_451 ();
 NOR2x1_ASAP7_75t_R _28989_ (.A(_01090_),
    .B(net264),
    .Y(_10161_));
 AO21x1_ASAP7_75t_R _28990_ (.A1(_08388_),
    .A2(net264),
    .B(_10161_),
    .Y(_03271_));
 TAPCELL_ASAP7_75t_R PHY_450 ();
 NOR2x1_ASAP7_75t_R _28992_ (.A(_01122_),
    .B(net264),
    .Y(_10163_));
 AO21x1_ASAP7_75t_R _28993_ (.A1(_08419_),
    .A2(net264),
    .B(_10163_),
    .Y(_03272_));
 TAPCELL_ASAP7_75t_R PHY_449 ();
 NOR2x1_ASAP7_75t_R _28995_ (.A(_01156_),
    .B(net266),
    .Y(_10165_));
 AO21x1_ASAP7_75t_R _28996_ (.A1(_08451_),
    .A2(net266),
    .B(_10165_),
    .Y(_03273_));
 TAPCELL_ASAP7_75t_R PHY_448 ();
 NOR2x1_ASAP7_75t_R _28998_ (.A(_01188_),
    .B(_10103_),
    .Y(_10167_));
 AO21x1_ASAP7_75t_R _28999_ (.A1(_08481_),
    .A2(_10103_),
    .B(_10167_),
    .Y(_03274_));
 TAPCELL_ASAP7_75t_R PHY_447 ();
 NOR2x1_ASAP7_75t_R _29001_ (.A(_01222_),
    .B(net266),
    .Y(_10169_));
 AO21x1_ASAP7_75t_R _29002_ (.A1(_08512_),
    .A2(net266),
    .B(_10169_),
    .Y(_03275_));
 TAPCELL_ASAP7_75t_R PHY_446 ();
 NOR2x1_ASAP7_75t_R _29004_ (.A(_01254_),
    .B(net264),
    .Y(_10171_));
 AO21x1_ASAP7_75t_R _29005_ (.A1(_08545_),
    .A2(net264),
    .B(_10171_),
    .Y(_03276_));
 TAPCELL_ASAP7_75t_R PHY_445 ();
 NOR2x1_ASAP7_75t_R _29007_ (.A(_01288_),
    .B(net265),
    .Y(_10173_));
 AO21x1_ASAP7_75t_R _29008_ (.A1(_08573_),
    .A2(net265),
    .B(_10173_),
    .Y(_03277_));
 AND2x6_ASAP7_75t_R _29009_ (.A(_06923_),
    .B(_10102_),
    .Y(_10174_));
 TAPCELL_ASAP7_75t_R PHY_444 ();
 TAPCELL_ASAP7_75t_R PHY_443 ();
 TAPCELL_ASAP7_75t_R PHY_442 ();
 NOR2x1_ASAP7_75t_R _29013_ (.A(_00304_),
    .B(_10174_),
    .Y(_10178_));
 AO21x1_ASAP7_75t_R _29014_ (.A1(_07180_),
    .A2(_10174_),
    .B(_10178_),
    .Y(_03278_));
 NOR2x1_ASAP7_75t_R _29015_ (.A(_00258_),
    .B(_10174_),
    .Y(_10179_));
 AO21x1_ASAP7_75t_R _29016_ (.A1(_07313_),
    .A2(_10174_),
    .B(_10179_),
    .Y(_03279_));
 NOR2x1_ASAP7_75t_R _29017_ (.A(_00366_),
    .B(_10174_),
    .Y(_10180_));
 AO21x1_ASAP7_75t_R _29018_ (.A1(_07398_),
    .A2(_10174_),
    .B(_10180_),
    .Y(_03280_));
 NOR2x1_ASAP7_75t_R _29019_ (.A(_00397_),
    .B(_10174_),
    .Y(_10181_));
 AO21x1_ASAP7_75t_R _29020_ (.A1(_07469_),
    .A2(_10174_),
    .B(_10181_),
    .Y(_03281_));
 NOR2x1_ASAP7_75t_R _29021_ (.A(_00427_),
    .B(_10174_),
    .Y(_10182_));
 AO21x1_ASAP7_75t_R _29022_ (.A1(_07534_),
    .A2(_10174_),
    .B(_10182_),
    .Y(_03282_));
 NOR2x1_ASAP7_75t_R _29023_ (.A(_00457_),
    .B(_10174_),
    .Y(_10183_));
 AO21x1_ASAP7_75t_R _29024_ (.A1(_07581_),
    .A2(_10174_),
    .B(_10183_),
    .Y(_03283_));
 NOR2x1_ASAP7_75t_R _29025_ (.A(_00487_),
    .B(_10174_),
    .Y(_10184_));
 AO21x1_ASAP7_75t_R _29026_ (.A1(net253),
    .A2(_10174_),
    .B(_10184_),
    .Y(_03284_));
 NOR2x1_ASAP7_75t_R _29027_ (.A(_00517_),
    .B(_10174_),
    .Y(_10185_));
 AO21x1_ASAP7_75t_R _29028_ (.A1(_07676_),
    .A2(_10174_),
    .B(_10185_),
    .Y(_03285_));
 TAPCELL_ASAP7_75t_R PHY_441 ();
 NOR2x1_ASAP7_75t_R _29030_ (.A(_00547_),
    .B(_10174_),
    .Y(_10187_));
 AO21x1_ASAP7_75t_R _29031_ (.A1(net252),
    .A2(_10174_),
    .B(_10187_),
    .Y(_03286_));
 NOR2x1_ASAP7_75t_R _29032_ (.A(_00577_),
    .B(_10174_),
    .Y(_10188_));
 AO21x1_ASAP7_75t_R _29033_ (.A1(_07780_),
    .A2(_10174_),
    .B(_10188_),
    .Y(_03287_));
 TAPCELL_ASAP7_75t_R PHY_440 ();
 NOR2x1_ASAP7_75t_R _29035_ (.A(_00607_),
    .B(_10174_),
    .Y(_10190_));
 AO21x1_ASAP7_75t_R _29036_ (.A1(_07817_),
    .A2(_10174_),
    .B(_10190_),
    .Y(_03288_));
 NOR2x1_ASAP7_75t_R _29037_ (.A(_00637_),
    .B(_10174_),
    .Y(_10191_));
 AO21x1_ASAP7_75t_R _29038_ (.A1(_07865_),
    .A2(_10174_),
    .B(_10191_),
    .Y(_03289_));
 NOR2x1_ASAP7_75t_R _29039_ (.A(_00336_),
    .B(_10174_),
    .Y(_10192_));
 AO21x1_ASAP7_75t_R _29040_ (.A1(_07908_),
    .A2(_10174_),
    .B(_10192_),
    .Y(_03290_));
 NOR2x1_ASAP7_75t_R _29041_ (.A(_00699_),
    .B(_10174_),
    .Y(_10193_));
 AO21x1_ASAP7_75t_R _29042_ (.A1(_07950_),
    .A2(_10174_),
    .B(_10193_),
    .Y(_03291_));
 NOR2x1_ASAP7_75t_R _29043_ (.A(_00731_),
    .B(_10174_),
    .Y(_10194_));
 AO21x1_ASAP7_75t_R _29044_ (.A1(_07990_),
    .A2(_10174_),
    .B(_10194_),
    .Y(_03292_));
 NOR2x1_ASAP7_75t_R _29045_ (.A(_00764_),
    .B(_10174_),
    .Y(_10195_));
 AO21x1_ASAP7_75t_R _29046_ (.A1(_08034_),
    .A2(_10174_),
    .B(_10195_),
    .Y(_03293_));
 NOR2x1_ASAP7_75t_R _29047_ (.A(_00797_),
    .B(_10174_),
    .Y(_10196_));
 AO21x1_ASAP7_75t_R _29048_ (.A1(_08073_),
    .A2(_10174_),
    .B(_10196_),
    .Y(_03294_));
 NOR2x1_ASAP7_75t_R _29049_ (.A(_00830_),
    .B(_10174_),
    .Y(_10197_));
 AO21x1_ASAP7_75t_R _29050_ (.A1(_08116_),
    .A2(_10174_),
    .B(_10197_),
    .Y(_03295_));
 TAPCELL_ASAP7_75t_R PHY_439 ();
 NOR2x1_ASAP7_75t_R _29052_ (.A(_00862_),
    .B(_10174_),
    .Y(_10199_));
 AO21x1_ASAP7_75t_R _29053_ (.A1(_08150_),
    .A2(_10174_),
    .B(_10199_),
    .Y(_03296_));
 NOR2x1_ASAP7_75t_R _29054_ (.A(_00895_),
    .B(_10174_),
    .Y(_10200_));
 AO21x1_ASAP7_75t_R _29055_ (.A1(_08187_),
    .A2(_10174_),
    .B(_10200_),
    .Y(_03297_));
 TAPCELL_ASAP7_75t_R PHY_438 ();
 NOR2x1_ASAP7_75t_R _29057_ (.A(_00927_),
    .B(_10174_),
    .Y(_10202_));
 AO21x1_ASAP7_75t_R _29058_ (.A1(_08219_),
    .A2(_10174_),
    .B(_10202_),
    .Y(_03298_));
 NOR2x1_ASAP7_75t_R _29059_ (.A(_00960_),
    .B(_10174_),
    .Y(_10203_));
 AO21x1_ASAP7_75t_R _29060_ (.A1(_08254_),
    .A2(_10174_),
    .B(_10203_),
    .Y(_03299_));
 NOR2x1_ASAP7_75t_R _29061_ (.A(_00992_),
    .B(_10174_),
    .Y(_10204_));
 AO21x1_ASAP7_75t_R _29062_ (.A1(net250),
    .A2(_10174_),
    .B(_10204_),
    .Y(_03300_));
 NOR2x1_ASAP7_75t_R _29063_ (.A(_01026_),
    .B(_10174_),
    .Y(_10205_));
 AO21x1_ASAP7_75t_R _29064_ (.A1(_08319_),
    .A2(_10174_),
    .B(_10205_),
    .Y(_03301_));
 NOR2x1_ASAP7_75t_R _29065_ (.A(_01058_),
    .B(_10174_),
    .Y(_10206_));
 AO21x1_ASAP7_75t_R _29066_ (.A1(_08357_),
    .A2(_10174_),
    .B(_10206_),
    .Y(_03302_));
 NOR2x1_ASAP7_75t_R _29067_ (.A(_01091_),
    .B(_10174_),
    .Y(_10207_));
 AO21x1_ASAP7_75t_R _29068_ (.A1(_08388_),
    .A2(_10174_),
    .B(_10207_),
    .Y(_03303_));
 NOR2x1_ASAP7_75t_R _29069_ (.A(_01123_),
    .B(_10174_),
    .Y(_10208_));
 AO21x1_ASAP7_75t_R _29070_ (.A1(_08419_),
    .A2(_10174_),
    .B(_10208_),
    .Y(_03304_));
 NOR2x1_ASAP7_75t_R _29071_ (.A(_01157_),
    .B(_10174_),
    .Y(_10209_));
 AO21x1_ASAP7_75t_R _29072_ (.A1(_08451_),
    .A2(_10174_),
    .B(_10209_),
    .Y(_03305_));
 NOR2x1_ASAP7_75t_R _29073_ (.A(_01189_),
    .B(_10174_),
    .Y(_10210_));
 AO21x1_ASAP7_75t_R _29074_ (.A1(_08481_),
    .A2(_10174_),
    .B(_10210_),
    .Y(_03306_));
 NOR2x1_ASAP7_75t_R _29075_ (.A(_01223_),
    .B(_10174_),
    .Y(_10211_));
 AO21x1_ASAP7_75t_R _29076_ (.A1(_08512_),
    .A2(_10174_),
    .B(_10211_),
    .Y(_03307_));
 NOR2x1_ASAP7_75t_R _29077_ (.A(_01255_),
    .B(_10174_),
    .Y(_10212_));
 AO21x1_ASAP7_75t_R _29078_ (.A1(_08545_),
    .A2(_10174_),
    .B(_10212_),
    .Y(_03308_));
 NOR2x1_ASAP7_75t_R _29079_ (.A(_01289_),
    .B(_10174_),
    .Y(_10213_));
 AO21x1_ASAP7_75t_R _29080_ (.A1(_08573_),
    .A2(_10174_),
    .B(_10213_),
    .Y(_03309_));
 AND2x6_ASAP7_75t_R _29081_ (.A(_09664_),
    .B(_10102_),
    .Y(_10214_));
 TAPCELL_ASAP7_75t_R PHY_437 ();
 TAPCELL_ASAP7_75t_R PHY_436 ();
 TAPCELL_ASAP7_75t_R PHY_435 ();
 NOR2x1_ASAP7_75t_R _29085_ (.A(_00305_),
    .B(_10214_),
    .Y(_10218_));
 AO21x1_ASAP7_75t_R _29086_ (.A1(_07180_),
    .A2(_10214_),
    .B(_10218_),
    .Y(_03310_));
 NOR2x1_ASAP7_75t_R _29087_ (.A(_00259_),
    .B(_10214_),
    .Y(_10219_));
 AO21x1_ASAP7_75t_R _29088_ (.A1(_07313_),
    .A2(_10214_),
    .B(_10219_),
    .Y(_03311_));
 NOR2x1_ASAP7_75t_R _29089_ (.A(_00367_),
    .B(_10214_),
    .Y(_10220_));
 AO21x1_ASAP7_75t_R _29090_ (.A1(_07398_),
    .A2(_10214_),
    .B(_10220_),
    .Y(_03312_));
 NOR2x1_ASAP7_75t_R _29091_ (.A(_00398_),
    .B(_10214_),
    .Y(_10221_));
 AO21x1_ASAP7_75t_R _29092_ (.A1(_07469_),
    .A2(_10214_),
    .B(_10221_),
    .Y(_03313_));
 NOR2x1_ASAP7_75t_R _29093_ (.A(_00428_),
    .B(_10214_),
    .Y(_10222_));
 AO21x1_ASAP7_75t_R _29094_ (.A1(_07534_),
    .A2(_10214_),
    .B(_10222_),
    .Y(_03314_));
 NOR2x1_ASAP7_75t_R _29095_ (.A(_00458_),
    .B(_10214_),
    .Y(_10223_));
 AO21x1_ASAP7_75t_R _29096_ (.A1(_07581_),
    .A2(_10214_),
    .B(_10223_),
    .Y(_03315_));
 NOR2x1_ASAP7_75t_R _29097_ (.A(_00488_),
    .B(_10214_),
    .Y(_10224_));
 AO21x1_ASAP7_75t_R _29098_ (.A1(net253),
    .A2(_10214_),
    .B(_10224_),
    .Y(_03316_));
 NOR2x1_ASAP7_75t_R _29099_ (.A(_00518_),
    .B(_10214_),
    .Y(_10225_));
 AO21x1_ASAP7_75t_R _29100_ (.A1(_07676_),
    .A2(_10214_),
    .B(_10225_),
    .Y(_03317_));
 TAPCELL_ASAP7_75t_R PHY_434 ();
 NOR2x1_ASAP7_75t_R _29102_ (.A(_00548_),
    .B(_10214_),
    .Y(_10227_));
 AO21x1_ASAP7_75t_R _29103_ (.A1(net252),
    .A2(_10214_),
    .B(_10227_),
    .Y(_03318_));
 NOR2x1_ASAP7_75t_R _29104_ (.A(_00578_),
    .B(_10214_),
    .Y(_10228_));
 AO21x1_ASAP7_75t_R _29105_ (.A1(_07780_),
    .A2(_10214_),
    .B(_10228_),
    .Y(_03319_));
 TAPCELL_ASAP7_75t_R PHY_433 ();
 NOR2x1_ASAP7_75t_R _29107_ (.A(_00608_),
    .B(_10214_),
    .Y(_10230_));
 AO21x1_ASAP7_75t_R _29108_ (.A1(_07817_),
    .A2(_10214_),
    .B(_10230_),
    .Y(_03320_));
 NOR2x1_ASAP7_75t_R _29109_ (.A(_00638_),
    .B(_10214_),
    .Y(_10231_));
 AO21x1_ASAP7_75t_R _29110_ (.A1(_07865_),
    .A2(_10214_),
    .B(_10231_),
    .Y(_03321_));
 NOR2x1_ASAP7_75t_R _29111_ (.A(_00337_),
    .B(_10214_),
    .Y(_10232_));
 AO21x1_ASAP7_75t_R _29112_ (.A1(_07908_),
    .A2(_10214_),
    .B(_10232_),
    .Y(_03322_));
 NOR2x1_ASAP7_75t_R _29113_ (.A(_00700_),
    .B(_10214_),
    .Y(_10233_));
 AO21x1_ASAP7_75t_R _29114_ (.A1(_07950_),
    .A2(_10214_),
    .B(_10233_),
    .Y(_03323_));
 NOR2x1_ASAP7_75t_R _29115_ (.A(_00732_),
    .B(_10214_),
    .Y(_10234_));
 AO21x1_ASAP7_75t_R _29116_ (.A1(_07990_),
    .A2(_10214_),
    .B(_10234_),
    .Y(_03324_));
 NOR2x1_ASAP7_75t_R _29117_ (.A(_00765_),
    .B(_10214_),
    .Y(_10235_));
 AO21x1_ASAP7_75t_R _29118_ (.A1(_08034_),
    .A2(_10214_),
    .B(_10235_),
    .Y(_03325_));
 NOR2x1_ASAP7_75t_R _29119_ (.A(_00798_),
    .B(_10214_),
    .Y(_10236_));
 AO21x1_ASAP7_75t_R _29120_ (.A1(_08073_),
    .A2(_10214_),
    .B(_10236_),
    .Y(_03326_));
 NOR2x1_ASAP7_75t_R _29121_ (.A(_00831_),
    .B(_10214_),
    .Y(_10237_));
 AO21x1_ASAP7_75t_R _29122_ (.A1(_08116_),
    .A2(_10214_),
    .B(_10237_),
    .Y(_03327_));
 TAPCELL_ASAP7_75t_R PHY_432 ();
 NOR2x1_ASAP7_75t_R _29124_ (.A(_00863_),
    .B(_10214_),
    .Y(_10239_));
 AO21x1_ASAP7_75t_R _29125_ (.A1(net251),
    .A2(_10214_),
    .B(_10239_),
    .Y(_03328_));
 NOR2x1_ASAP7_75t_R _29126_ (.A(_00896_),
    .B(_10214_),
    .Y(_10240_));
 AO21x1_ASAP7_75t_R _29127_ (.A1(_08187_),
    .A2(_10214_),
    .B(_10240_),
    .Y(_03329_));
 TAPCELL_ASAP7_75t_R PHY_431 ();
 NOR2x1_ASAP7_75t_R _29129_ (.A(_00928_),
    .B(_10214_),
    .Y(_10242_));
 AO21x1_ASAP7_75t_R _29130_ (.A1(_08219_),
    .A2(_10214_),
    .B(_10242_),
    .Y(_03330_));
 NOR2x1_ASAP7_75t_R _29131_ (.A(_00961_),
    .B(_10214_),
    .Y(_10243_));
 AO21x1_ASAP7_75t_R _29132_ (.A1(_08254_),
    .A2(_10214_),
    .B(_10243_),
    .Y(_03331_));
 NOR2x1_ASAP7_75t_R _29133_ (.A(_00993_),
    .B(_10214_),
    .Y(_10244_));
 AO21x1_ASAP7_75t_R _29134_ (.A1(net250),
    .A2(_10214_),
    .B(_10244_),
    .Y(_03332_));
 NOR2x1_ASAP7_75t_R _29135_ (.A(_01027_),
    .B(_10214_),
    .Y(_10245_));
 AO21x1_ASAP7_75t_R _29136_ (.A1(_08319_),
    .A2(_10214_),
    .B(_10245_),
    .Y(_03333_));
 NOR2x1_ASAP7_75t_R _29137_ (.A(_01059_),
    .B(_10214_),
    .Y(_10246_));
 AO21x1_ASAP7_75t_R _29138_ (.A1(_08357_),
    .A2(_10214_),
    .B(_10246_),
    .Y(_03334_));
 NOR2x1_ASAP7_75t_R _29139_ (.A(_01092_),
    .B(_10214_),
    .Y(_10247_));
 AO21x1_ASAP7_75t_R _29140_ (.A1(_08388_),
    .A2(_10214_),
    .B(_10247_),
    .Y(_03335_));
 NOR2x1_ASAP7_75t_R _29141_ (.A(_01124_),
    .B(_10214_),
    .Y(_10248_));
 AO21x1_ASAP7_75t_R _29142_ (.A1(_08419_),
    .A2(_10214_),
    .B(_10248_),
    .Y(_03336_));
 NOR2x1_ASAP7_75t_R _29143_ (.A(_01158_),
    .B(_10214_),
    .Y(_10249_));
 AO21x1_ASAP7_75t_R _29144_ (.A1(_08451_),
    .A2(_10214_),
    .B(_10249_),
    .Y(_03337_));
 NOR2x1_ASAP7_75t_R _29145_ (.A(_01190_),
    .B(_10214_),
    .Y(_10250_));
 AO21x1_ASAP7_75t_R _29146_ (.A1(_08481_),
    .A2(_10214_),
    .B(_10250_),
    .Y(_03338_));
 NOR2x1_ASAP7_75t_R _29147_ (.A(_01224_),
    .B(_10214_),
    .Y(_10251_));
 AO21x1_ASAP7_75t_R _29148_ (.A1(_08512_),
    .A2(_10214_),
    .B(_10251_),
    .Y(_03339_));
 NOR2x1_ASAP7_75t_R _29149_ (.A(_01256_),
    .B(_10214_),
    .Y(_10252_));
 AO21x1_ASAP7_75t_R _29150_ (.A1(_08545_),
    .A2(_10214_),
    .B(_10252_),
    .Y(_03340_));
 NOR2x1_ASAP7_75t_R _29151_ (.A(_01290_),
    .B(_10214_),
    .Y(_10253_));
 AO21x1_ASAP7_75t_R _29152_ (.A1(_08573_),
    .A2(_10214_),
    .B(_10253_),
    .Y(_03341_));
 AND2x6_ASAP7_75t_R _29153_ (.A(_09737_),
    .B(_10102_),
    .Y(_10254_));
 TAPCELL_ASAP7_75t_R PHY_430 ();
 TAPCELL_ASAP7_75t_R PHY_429 ();
 TAPCELL_ASAP7_75t_R PHY_428 ();
 NOR2x1_ASAP7_75t_R _29157_ (.A(_00306_),
    .B(_10254_),
    .Y(_10258_));
 AO21x1_ASAP7_75t_R _29158_ (.A1(_07180_),
    .A2(_10254_),
    .B(_10258_),
    .Y(_03342_));
 NOR2x1_ASAP7_75t_R _29159_ (.A(_00260_),
    .B(_10254_),
    .Y(_10259_));
 AO21x1_ASAP7_75t_R _29160_ (.A1(_07313_),
    .A2(_10254_),
    .B(_10259_),
    .Y(_03343_));
 NOR2x1_ASAP7_75t_R _29161_ (.A(_00368_),
    .B(_10254_),
    .Y(_10260_));
 AO21x1_ASAP7_75t_R _29162_ (.A1(_07398_),
    .A2(_10254_),
    .B(_10260_),
    .Y(_03344_));
 NOR2x1_ASAP7_75t_R _29163_ (.A(_00399_),
    .B(_10254_),
    .Y(_10261_));
 AO21x1_ASAP7_75t_R _29164_ (.A1(_07469_),
    .A2(_10254_),
    .B(_10261_),
    .Y(_03345_));
 NOR2x1_ASAP7_75t_R _29165_ (.A(_00429_),
    .B(_10254_),
    .Y(_10262_));
 AO21x1_ASAP7_75t_R _29166_ (.A1(_07534_),
    .A2(_10254_),
    .B(_10262_),
    .Y(_03346_));
 NOR2x1_ASAP7_75t_R _29167_ (.A(_00459_),
    .B(_10254_),
    .Y(_10263_));
 AO21x1_ASAP7_75t_R _29168_ (.A1(_07581_),
    .A2(_10254_),
    .B(_10263_),
    .Y(_03347_));
 NOR2x1_ASAP7_75t_R _29169_ (.A(_00489_),
    .B(_10254_),
    .Y(_10264_));
 AO21x1_ASAP7_75t_R _29170_ (.A1(net253),
    .A2(_10254_),
    .B(_10264_),
    .Y(_03348_));
 NOR2x1_ASAP7_75t_R _29171_ (.A(_00519_),
    .B(_10254_),
    .Y(_10265_));
 AO21x1_ASAP7_75t_R _29172_ (.A1(_07676_),
    .A2(_10254_),
    .B(_10265_),
    .Y(_03349_));
 TAPCELL_ASAP7_75t_R PHY_427 ();
 NOR2x1_ASAP7_75t_R _29174_ (.A(_00549_),
    .B(_10254_),
    .Y(_10267_));
 AO21x1_ASAP7_75t_R _29175_ (.A1(net252),
    .A2(_10254_),
    .B(_10267_),
    .Y(_03350_));
 NOR2x1_ASAP7_75t_R _29176_ (.A(_00579_),
    .B(_10254_),
    .Y(_10268_));
 AO21x1_ASAP7_75t_R _29177_ (.A1(_07780_),
    .A2(_10254_),
    .B(_10268_),
    .Y(_03351_));
 TAPCELL_ASAP7_75t_R PHY_426 ();
 NOR2x1_ASAP7_75t_R _29179_ (.A(_00609_),
    .B(_10254_),
    .Y(_10270_));
 AO21x1_ASAP7_75t_R _29180_ (.A1(_07817_),
    .A2(_10254_),
    .B(_10270_),
    .Y(_03352_));
 NOR2x1_ASAP7_75t_R _29181_ (.A(_00639_),
    .B(_10254_),
    .Y(_10271_));
 AO21x1_ASAP7_75t_R _29182_ (.A1(_07865_),
    .A2(_10254_),
    .B(_10271_),
    .Y(_03353_));
 NOR2x1_ASAP7_75t_R _29183_ (.A(_00338_),
    .B(_10254_),
    .Y(_10272_));
 AO21x1_ASAP7_75t_R _29184_ (.A1(_07908_),
    .A2(_10254_),
    .B(_10272_),
    .Y(_03354_));
 NOR2x1_ASAP7_75t_R _29185_ (.A(_00701_),
    .B(_10254_),
    .Y(_10273_));
 AO21x1_ASAP7_75t_R _29186_ (.A1(_07950_),
    .A2(_10254_),
    .B(_10273_),
    .Y(_03355_));
 NOR2x1_ASAP7_75t_R _29187_ (.A(_00733_),
    .B(_10254_),
    .Y(_10274_));
 AO21x1_ASAP7_75t_R _29188_ (.A1(_07990_),
    .A2(_10254_),
    .B(_10274_),
    .Y(_03356_));
 NOR2x1_ASAP7_75t_R _29189_ (.A(_00766_),
    .B(_10254_),
    .Y(_10275_));
 AO21x1_ASAP7_75t_R _29190_ (.A1(_08034_),
    .A2(_10254_),
    .B(_10275_),
    .Y(_03357_));
 NOR2x1_ASAP7_75t_R _29191_ (.A(_00799_),
    .B(_10254_),
    .Y(_10276_));
 AO21x1_ASAP7_75t_R _29192_ (.A1(_08073_),
    .A2(_10254_),
    .B(_10276_),
    .Y(_03358_));
 NOR2x1_ASAP7_75t_R _29193_ (.A(_00832_),
    .B(_10254_),
    .Y(_10277_));
 AO21x1_ASAP7_75t_R _29194_ (.A1(_08116_),
    .A2(_10254_),
    .B(_10277_),
    .Y(_03359_));
 TAPCELL_ASAP7_75t_R PHY_425 ();
 NOR2x1_ASAP7_75t_R _29196_ (.A(_00864_),
    .B(_10254_),
    .Y(_10279_));
 AO21x1_ASAP7_75t_R _29197_ (.A1(_08150_),
    .A2(_10254_),
    .B(_10279_),
    .Y(_03360_));
 NOR2x1_ASAP7_75t_R _29198_ (.A(_00897_),
    .B(_10254_),
    .Y(_10280_));
 AO21x1_ASAP7_75t_R _29199_ (.A1(_08187_),
    .A2(_10254_),
    .B(_10280_),
    .Y(_03361_));
 TAPCELL_ASAP7_75t_R PHY_424 ();
 NOR2x1_ASAP7_75t_R _29201_ (.A(_00929_),
    .B(_10254_),
    .Y(_10282_));
 AO21x1_ASAP7_75t_R _29202_ (.A1(_08219_),
    .A2(_10254_),
    .B(_10282_),
    .Y(_03362_));
 NOR2x1_ASAP7_75t_R _29203_ (.A(_00962_),
    .B(_10254_),
    .Y(_10283_));
 AO21x1_ASAP7_75t_R _29204_ (.A1(_08254_),
    .A2(_10254_),
    .B(_10283_),
    .Y(_03363_));
 NOR2x1_ASAP7_75t_R _29205_ (.A(_00994_),
    .B(_10254_),
    .Y(_10284_));
 AO21x1_ASAP7_75t_R _29206_ (.A1(net250),
    .A2(_10254_),
    .B(_10284_),
    .Y(_03364_));
 NOR2x1_ASAP7_75t_R _29207_ (.A(_01028_),
    .B(_10254_),
    .Y(_10285_));
 AO21x1_ASAP7_75t_R _29208_ (.A1(_08319_),
    .A2(_10254_),
    .B(_10285_),
    .Y(_03365_));
 NOR2x1_ASAP7_75t_R _29209_ (.A(_01060_),
    .B(_10254_),
    .Y(_10286_));
 AO21x1_ASAP7_75t_R _29210_ (.A1(_08357_),
    .A2(_10254_),
    .B(_10286_),
    .Y(_03366_));
 NOR2x1_ASAP7_75t_R _29211_ (.A(_01093_),
    .B(_10254_),
    .Y(_10287_));
 AO21x1_ASAP7_75t_R _29212_ (.A1(_08388_),
    .A2(_10254_),
    .B(_10287_),
    .Y(_03367_));
 NOR2x1_ASAP7_75t_R _29213_ (.A(_01125_),
    .B(_10254_),
    .Y(_10288_));
 AO21x1_ASAP7_75t_R _29214_ (.A1(_08419_),
    .A2(_10254_),
    .B(_10288_),
    .Y(_03368_));
 NOR2x1_ASAP7_75t_R _29215_ (.A(_01159_),
    .B(_10254_),
    .Y(_10289_));
 AO21x1_ASAP7_75t_R _29216_ (.A1(_08451_),
    .A2(_10254_),
    .B(_10289_),
    .Y(_03369_));
 NOR2x1_ASAP7_75t_R _29217_ (.A(_01191_),
    .B(_10254_),
    .Y(_10290_));
 AO21x1_ASAP7_75t_R _29218_ (.A1(_08481_),
    .A2(_10254_),
    .B(_10290_),
    .Y(_03370_));
 NOR2x1_ASAP7_75t_R _29219_ (.A(_01225_),
    .B(_10254_),
    .Y(_10291_));
 AO21x1_ASAP7_75t_R _29220_ (.A1(_08512_),
    .A2(_10254_),
    .B(_10291_),
    .Y(_03371_));
 NOR2x1_ASAP7_75t_R _29221_ (.A(_01257_),
    .B(_10254_),
    .Y(_10292_));
 AO21x1_ASAP7_75t_R _29222_ (.A1(_08545_),
    .A2(_10254_),
    .B(_10292_),
    .Y(_03372_));
 NOR2x1_ASAP7_75t_R _29223_ (.A(_01291_),
    .B(_10254_),
    .Y(_10293_));
 AO21x1_ASAP7_75t_R _29224_ (.A1(_08573_),
    .A2(_10254_),
    .B(_10293_),
    .Y(_03373_));
 AND3x4_ASAP7_75t_R _29225_ (.A(_14027_),
    .B(_14606_),
    .C(_06922_),
    .Y(_10294_));
 TAPCELL_ASAP7_75t_R PHY_423 ();
 TAPCELL_ASAP7_75t_R PHY_422 ();
 TAPCELL_ASAP7_75t_R PHY_421 ();
 NOR2x1_ASAP7_75t_R _29229_ (.A(_00307_),
    .B(_10294_),
    .Y(_10298_));
 AO21x1_ASAP7_75t_R _29230_ (.A1(_07180_),
    .A2(_10294_),
    .B(_10298_),
    .Y(_03374_));
 NOR2x1_ASAP7_75t_R _29231_ (.A(_00261_),
    .B(_10294_),
    .Y(_10299_));
 AO21x1_ASAP7_75t_R _29232_ (.A1(_07313_),
    .A2(_10294_),
    .B(_10299_),
    .Y(_03375_));
 NOR2x1_ASAP7_75t_R _29233_ (.A(_00369_),
    .B(_10294_),
    .Y(_10300_));
 AO21x1_ASAP7_75t_R _29234_ (.A1(_07398_),
    .A2(_10294_),
    .B(_10300_),
    .Y(_03376_));
 NOR2x1_ASAP7_75t_R _29235_ (.A(_00400_),
    .B(_10294_),
    .Y(_10301_));
 AO21x1_ASAP7_75t_R _29236_ (.A1(_07469_),
    .A2(_10294_),
    .B(_10301_),
    .Y(_03377_));
 NOR2x1_ASAP7_75t_R _29237_ (.A(_00430_),
    .B(_10294_),
    .Y(_10302_));
 AO21x1_ASAP7_75t_R _29238_ (.A1(_07534_),
    .A2(_10294_),
    .B(_10302_),
    .Y(_03378_));
 NOR2x1_ASAP7_75t_R _29239_ (.A(_00460_),
    .B(_10294_),
    .Y(_10303_));
 AO21x1_ASAP7_75t_R _29240_ (.A1(_07581_),
    .A2(_10294_),
    .B(_10303_),
    .Y(_03379_));
 NOR2x1_ASAP7_75t_R _29241_ (.A(_00490_),
    .B(_10294_),
    .Y(_10304_));
 AO21x1_ASAP7_75t_R _29242_ (.A1(_07620_),
    .A2(_10294_),
    .B(_10304_),
    .Y(_03380_));
 NOR2x1_ASAP7_75t_R _29243_ (.A(_00520_),
    .B(_10294_),
    .Y(_10305_));
 AO21x1_ASAP7_75t_R _29244_ (.A1(_07676_),
    .A2(_10294_),
    .B(_10305_),
    .Y(_03381_));
 TAPCELL_ASAP7_75t_R PHY_420 ();
 NOR2x1_ASAP7_75t_R _29246_ (.A(_00550_),
    .B(_10294_),
    .Y(_10307_));
 AO21x1_ASAP7_75t_R _29247_ (.A1(_07738_),
    .A2(_10294_),
    .B(_10307_),
    .Y(_03382_));
 NOR2x1_ASAP7_75t_R _29248_ (.A(_00580_),
    .B(_10294_),
    .Y(_10308_));
 AO21x1_ASAP7_75t_R _29249_ (.A1(_07780_),
    .A2(_10294_),
    .B(_10308_),
    .Y(_03383_));
 TAPCELL_ASAP7_75t_R PHY_419 ();
 NOR2x1_ASAP7_75t_R _29251_ (.A(_00610_),
    .B(_10294_),
    .Y(_10310_));
 AO21x1_ASAP7_75t_R _29252_ (.A1(_07817_),
    .A2(_10294_),
    .B(_10310_),
    .Y(_03384_));
 NOR2x1_ASAP7_75t_R _29253_ (.A(_00640_),
    .B(_10294_),
    .Y(_10311_));
 AO21x1_ASAP7_75t_R _29254_ (.A1(_07865_),
    .A2(_10294_),
    .B(_10311_),
    .Y(_03385_));
 NOR2x1_ASAP7_75t_R _29255_ (.A(_00339_),
    .B(_10294_),
    .Y(_10312_));
 AO21x1_ASAP7_75t_R _29256_ (.A1(_07908_),
    .A2(_10294_),
    .B(_10312_),
    .Y(_03386_));
 NOR2x1_ASAP7_75t_R _29257_ (.A(_00702_),
    .B(_10294_),
    .Y(_10313_));
 AO21x1_ASAP7_75t_R _29258_ (.A1(_07950_),
    .A2(_10294_),
    .B(_10313_),
    .Y(_03387_));
 NOR2x1_ASAP7_75t_R _29259_ (.A(_00734_),
    .B(_10294_),
    .Y(_10314_));
 AO21x1_ASAP7_75t_R _29260_ (.A1(_07990_),
    .A2(_10294_),
    .B(_10314_),
    .Y(_03388_));
 NOR2x1_ASAP7_75t_R _29261_ (.A(_00767_),
    .B(_10294_),
    .Y(_10315_));
 AO21x1_ASAP7_75t_R _29262_ (.A1(_08034_),
    .A2(_10294_),
    .B(_10315_),
    .Y(_03389_));
 NOR2x1_ASAP7_75t_R _29263_ (.A(_00800_),
    .B(_10294_),
    .Y(_10316_));
 AO21x1_ASAP7_75t_R _29264_ (.A1(_08073_),
    .A2(_10294_),
    .B(_10316_),
    .Y(_03390_));
 NOR2x1_ASAP7_75t_R _29265_ (.A(_00833_),
    .B(_10294_),
    .Y(_10317_));
 AO21x1_ASAP7_75t_R _29266_ (.A1(_08116_),
    .A2(_10294_),
    .B(_10317_),
    .Y(_03391_));
 TAPCELL_ASAP7_75t_R PHY_418 ();
 NOR2x1_ASAP7_75t_R _29268_ (.A(_00865_),
    .B(_10294_),
    .Y(_10319_));
 AO21x1_ASAP7_75t_R _29269_ (.A1(net251),
    .A2(_10294_),
    .B(_10319_),
    .Y(_03392_));
 NOR2x1_ASAP7_75t_R _29270_ (.A(_00898_),
    .B(_10294_),
    .Y(_10320_));
 AO21x1_ASAP7_75t_R _29271_ (.A1(_08187_),
    .A2(_10294_),
    .B(_10320_),
    .Y(_03393_));
 TAPCELL_ASAP7_75t_R PHY_417 ();
 NOR2x1_ASAP7_75t_R _29273_ (.A(_00930_),
    .B(_10294_),
    .Y(_10322_));
 AO21x1_ASAP7_75t_R _29274_ (.A1(_08219_),
    .A2(_10294_),
    .B(_10322_),
    .Y(_03394_));
 NOR2x1_ASAP7_75t_R _29275_ (.A(_00963_),
    .B(_10294_),
    .Y(_10323_));
 AO21x1_ASAP7_75t_R _29276_ (.A1(_08254_),
    .A2(_10294_),
    .B(_10323_),
    .Y(_03395_));
 NOR2x1_ASAP7_75t_R _29277_ (.A(_00995_),
    .B(_10294_),
    .Y(_10324_));
 AO21x1_ASAP7_75t_R _29278_ (.A1(net250),
    .A2(_10294_),
    .B(_10324_),
    .Y(_03396_));
 NOR2x1_ASAP7_75t_R _29279_ (.A(_01029_),
    .B(_10294_),
    .Y(_10325_));
 AO21x1_ASAP7_75t_R _29280_ (.A1(_08319_),
    .A2(_10294_),
    .B(_10325_),
    .Y(_03397_));
 NOR2x1_ASAP7_75t_R _29281_ (.A(_01061_),
    .B(_10294_),
    .Y(_10326_));
 AO21x1_ASAP7_75t_R _29282_ (.A1(_08357_),
    .A2(_10294_),
    .B(_10326_),
    .Y(_03398_));
 NOR2x1_ASAP7_75t_R _29283_ (.A(_01094_),
    .B(_10294_),
    .Y(_10327_));
 AO21x1_ASAP7_75t_R _29284_ (.A1(_08388_),
    .A2(_10294_),
    .B(_10327_),
    .Y(_03399_));
 NOR2x1_ASAP7_75t_R _29285_ (.A(_01126_),
    .B(_10294_),
    .Y(_10328_));
 AO21x1_ASAP7_75t_R _29286_ (.A1(_08419_),
    .A2(_10294_),
    .B(_10328_),
    .Y(_03400_));
 NOR2x1_ASAP7_75t_R _29287_ (.A(_01160_),
    .B(_10294_),
    .Y(_10329_));
 AO21x1_ASAP7_75t_R _29288_ (.A1(_08451_),
    .A2(_10294_),
    .B(_10329_),
    .Y(_03401_));
 NOR2x1_ASAP7_75t_R _29289_ (.A(_01192_),
    .B(_10294_),
    .Y(_10330_));
 AO21x1_ASAP7_75t_R _29290_ (.A1(_08481_),
    .A2(_10294_),
    .B(_10330_),
    .Y(_03402_));
 NOR2x1_ASAP7_75t_R _29291_ (.A(_01226_),
    .B(_10294_),
    .Y(_10331_));
 AO21x1_ASAP7_75t_R _29292_ (.A1(_08512_),
    .A2(_10294_),
    .B(_10331_),
    .Y(_03403_));
 NOR2x1_ASAP7_75t_R _29293_ (.A(_01258_),
    .B(_10294_),
    .Y(_10332_));
 AO21x1_ASAP7_75t_R _29294_ (.A1(_08545_),
    .A2(_10294_),
    .B(_10332_),
    .Y(_03404_));
 NOR2x1_ASAP7_75t_R _29295_ (.A(_01292_),
    .B(_10294_),
    .Y(_10333_));
 AO21x1_ASAP7_75t_R _29296_ (.A1(_08573_),
    .A2(_10294_),
    .B(_10333_),
    .Y(_03405_));
 AND2x6_ASAP7_75t_R _29297_ (.A(_14027_),
    .B(_06922_),
    .Y(_10334_));
 TAPCELL_ASAP7_75t_R PHY_416 ();
 AND3x4_ASAP7_75t_R _29299_ (.A(_06881_),
    .B(_06882_),
    .C(_10334_),
    .Y(_10336_));
 TAPCELL_ASAP7_75t_R PHY_415 ();
 TAPCELL_ASAP7_75t_R PHY_414 ();
 TAPCELL_ASAP7_75t_R PHY_413 ();
 NOR2x1_ASAP7_75t_R _29303_ (.A(_00308_),
    .B(_10336_),
    .Y(_10340_));
 AO21x1_ASAP7_75t_R _29304_ (.A1(_07180_),
    .A2(_10336_),
    .B(_10340_),
    .Y(_03406_));
 NOR2x1_ASAP7_75t_R _29305_ (.A(_00262_),
    .B(_10336_),
    .Y(_10341_));
 AO21x1_ASAP7_75t_R _29306_ (.A1(_07313_),
    .A2(_10336_),
    .B(_10341_),
    .Y(_03407_));
 NOR2x1_ASAP7_75t_R _29307_ (.A(_00370_),
    .B(_10336_),
    .Y(_10342_));
 AO21x1_ASAP7_75t_R _29308_ (.A1(_07398_),
    .A2(_10336_),
    .B(_10342_),
    .Y(_03408_));
 NOR2x1_ASAP7_75t_R _29309_ (.A(_00401_),
    .B(_10336_),
    .Y(_10343_));
 AO21x1_ASAP7_75t_R _29310_ (.A1(_07469_),
    .A2(_10336_),
    .B(_10343_),
    .Y(_03409_));
 NOR2x1_ASAP7_75t_R _29311_ (.A(_00431_),
    .B(_10336_),
    .Y(_10344_));
 AO21x1_ASAP7_75t_R _29312_ (.A1(_07534_),
    .A2(_10336_),
    .B(_10344_),
    .Y(_03410_));
 NOR2x1_ASAP7_75t_R _29313_ (.A(_00461_),
    .B(_10336_),
    .Y(_10345_));
 AO21x1_ASAP7_75t_R _29314_ (.A1(_07581_),
    .A2(_10336_),
    .B(_10345_),
    .Y(_03411_));
 NOR2x1_ASAP7_75t_R _29315_ (.A(_00491_),
    .B(_10336_),
    .Y(_10346_));
 AO21x1_ASAP7_75t_R _29316_ (.A1(_07620_),
    .A2(_10336_),
    .B(_10346_),
    .Y(_03412_));
 NOR2x1_ASAP7_75t_R _29317_ (.A(_00521_),
    .B(_10336_),
    .Y(_10347_));
 AO21x1_ASAP7_75t_R _29318_ (.A1(_07676_),
    .A2(_10336_),
    .B(_10347_),
    .Y(_03413_));
 TAPCELL_ASAP7_75t_R PHY_412 ();
 NOR2x1_ASAP7_75t_R _29320_ (.A(_00551_),
    .B(_10336_),
    .Y(_10349_));
 AO21x1_ASAP7_75t_R _29321_ (.A1(net252),
    .A2(_10336_),
    .B(_10349_),
    .Y(_03414_));
 NOR2x1_ASAP7_75t_R _29322_ (.A(_00581_),
    .B(_10336_),
    .Y(_10350_));
 AO21x1_ASAP7_75t_R _29323_ (.A1(_07780_),
    .A2(_10336_),
    .B(_10350_),
    .Y(_03415_));
 TAPCELL_ASAP7_75t_R PHY_411 ();
 NOR2x1_ASAP7_75t_R _29325_ (.A(_00611_),
    .B(_10336_),
    .Y(_10352_));
 AO21x1_ASAP7_75t_R _29326_ (.A1(_07817_),
    .A2(_10336_),
    .B(_10352_),
    .Y(_03416_));
 NOR2x1_ASAP7_75t_R _29327_ (.A(_00641_),
    .B(_10336_),
    .Y(_10353_));
 AO21x1_ASAP7_75t_R _29328_ (.A1(_07865_),
    .A2(_10336_),
    .B(_10353_),
    .Y(_03417_));
 NOR2x1_ASAP7_75t_R _29329_ (.A(_00340_),
    .B(_10336_),
    .Y(_10354_));
 AO21x1_ASAP7_75t_R _29330_ (.A1(_07908_),
    .A2(_10336_),
    .B(_10354_),
    .Y(_03418_));
 NOR2x1_ASAP7_75t_R _29331_ (.A(_00703_),
    .B(_10336_),
    .Y(_10355_));
 AO21x1_ASAP7_75t_R _29332_ (.A1(_07950_),
    .A2(_10336_),
    .B(_10355_),
    .Y(_03419_));
 NOR2x1_ASAP7_75t_R _29333_ (.A(_00735_),
    .B(_10336_),
    .Y(_10356_));
 AO21x1_ASAP7_75t_R _29334_ (.A1(_07990_),
    .A2(_10336_),
    .B(_10356_),
    .Y(_03420_));
 NOR2x1_ASAP7_75t_R _29335_ (.A(_00768_),
    .B(_10336_),
    .Y(_10357_));
 AO21x1_ASAP7_75t_R _29336_ (.A1(_08034_),
    .A2(_10336_),
    .B(_10357_),
    .Y(_03421_));
 NOR2x1_ASAP7_75t_R _29337_ (.A(_00801_),
    .B(_10336_),
    .Y(_10358_));
 AO21x1_ASAP7_75t_R _29338_ (.A1(_08073_),
    .A2(_10336_),
    .B(_10358_),
    .Y(_03422_));
 NOR2x1_ASAP7_75t_R _29339_ (.A(_00834_),
    .B(_10336_),
    .Y(_10359_));
 AO21x1_ASAP7_75t_R _29340_ (.A1(_08116_),
    .A2(_10336_),
    .B(_10359_),
    .Y(_03423_));
 TAPCELL_ASAP7_75t_R PHY_410 ();
 NOR2x1_ASAP7_75t_R _29342_ (.A(_00866_),
    .B(_10336_),
    .Y(_10361_));
 AO21x1_ASAP7_75t_R _29343_ (.A1(net251),
    .A2(_10336_),
    .B(_10361_),
    .Y(_03424_));
 NOR2x1_ASAP7_75t_R _29344_ (.A(_00899_),
    .B(_10336_),
    .Y(_10362_));
 AO21x1_ASAP7_75t_R _29345_ (.A1(_08187_),
    .A2(_10336_),
    .B(_10362_),
    .Y(_03425_));
 TAPCELL_ASAP7_75t_R PHY_409 ();
 NOR2x1_ASAP7_75t_R _29347_ (.A(_00931_),
    .B(_10336_),
    .Y(_10364_));
 AO21x1_ASAP7_75t_R _29348_ (.A1(_08219_),
    .A2(_10336_),
    .B(_10364_),
    .Y(_03426_));
 NOR2x1_ASAP7_75t_R _29349_ (.A(_00964_),
    .B(_10336_),
    .Y(_10365_));
 AO21x1_ASAP7_75t_R _29350_ (.A1(_08254_),
    .A2(_10336_),
    .B(_10365_),
    .Y(_03427_));
 NOR2x1_ASAP7_75t_R _29351_ (.A(_00996_),
    .B(_10336_),
    .Y(_10366_));
 AO21x1_ASAP7_75t_R _29352_ (.A1(net250),
    .A2(_10336_),
    .B(_10366_),
    .Y(_03428_));
 NOR2x1_ASAP7_75t_R _29353_ (.A(_01030_),
    .B(_10336_),
    .Y(_10367_));
 AO21x1_ASAP7_75t_R _29354_ (.A1(_08319_),
    .A2(_10336_),
    .B(_10367_),
    .Y(_03429_));
 NOR2x1_ASAP7_75t_R _29355_ (.A(_01062_),
    .B(_10336_),
    .Y(_10368_));
 AO21x1_ASAP7_75t_R _29356_ (.A1(_08357_),
    .A2(_10336_),
    .B(_10368_),
    .Y(_03430_));
 NOR2x1_ASAP7_75t_R _29357_ (.A(_01095_),
    .B(_10336_),
    .Y(_10369_));
 AO21x1_ASAP7_75t_R _29358_ (.A1(_08388_),
    .A2(_10336_),
    .B(_10369_),
    .Y(_03431_));
 NOR2x1_ASAP7_75t_R _29359_ (.A(_01127_),
    .B(_10336_),
    .Y(_10370_));
 AO21x1_ASAP7_75t_R _29360_ (.A1(_08419_),
    .A2(_10336_),
    .B(_10370_),
    .Y(_03432_));
 NOR2x1_ASAP7_75t_R _29361_ (.A(_01161_),
    .B(_10336_),
    .Y(_10371_));
 AO21x1_ASAP7_75t_R _29362_ (.A1(_08451_),
    .A2(_10336_),
    .B(_10371_),
    .Y(_03433_));
 NOR2x1_ASAP7_75t_R _29363_ (.A(_01193_),
    .B(_10336_),
    .Y(_10372_));
 AO21x1_ASAP7_75t_R _29364_ (.A1(_08481_),
    .A2(_10336_),
    .B(_10372_),
    .Y(_03434_));
 NOR2x1_ASAP7_75t_R _29365_ (.A(_01227_),
    .B(_10336_),
    .Y(_10373_));
 AO21x1_ASAP7_75t_R _29366_ (.A1(_08512_),
    .A2(_10336_),
    .B(_10373_),
    .Y(_03435_));
 NOR2x1_ASAP7_75t_R _29367_ (.A(_01259_),
    .B(_10336_),
    .Y(_10374_));
 AO21x1_ASAP7_75t_R _29368_ (.A1(_08545_),
    .A2(_10336_),
    .B(_10374_),
    .Y(_03436_));
 NOR2x1_ASAP7_75t_R _29369_ (.A(_01293_),
    .B(_10336_),
    .Y(_10375_));
 AO21x1_ASAP7_75t_R _29370_ (.A1(_08573_),
    .A2(_10336_),
    .B(_10375_),
    .Y(_03437_));
 AND3x4_ASAP7_75t_R _29371_ (.A(_06881_),
    .B(_09663_),
    .C(_10334_),
    .Y(_10376_));
 TAPCELL_ASAP7_75t_R PHY_408 ();
 TAPCELL_ASAP7_75t_R PHY_407 ();
 TAPCELL_ASAP7_75t_R PHY_406 ();
 NOR2x1_ASAP7_75t_R _29375_ (.A(_00309_),
    .B(_10376_),
    .Y(_10380_));
 AO21x1_ASAP7_75t_R _29376_ (.A1(_07180_),
    .A2(_10376_),
    .B(_10380_),
    .Y(_03438_));
 NOR2x1_ASAP7_75t_R _29377_ (.A(_00263_),
    .B(_10376_),
    .Y(_10381_));
 AO21x1_ASAP7_75t_R _29378_ (.A1(_07313_),
    .A2(_10376_),
    .B(_10381_),
    .Y(_03439_));
 NOR2x1_ASAP7_75t_R _29379_ (.A(_00371_),
    .B(_10376_),
    .Y(_10382_));
 AO21x1_ASAP7_75t_R _29380_ (.A1(_07398_),
    .A2(_10376_),
    .B(_10382_),
    .Y(_03440_));
 NOR2x1_ASAP7_75t_R _29381_ (.A(_00402_),
    .B(_10376_),
    .Y(_10383_));
 AO21x1_ASAP7_75t_R _29382_ (.A1(_07469_),
    .A2(_10376_),
    .B(_10383_),
    .Y(_03441_));
 NOR2x1_ASAP7_75t_R _29383_ (.A(_00432_),
    .B(_10376_),
    .Y(_10384_));
 AO21x1_ASAP7_75t_R _29384_ (.A1(_07534_),
    .A2(_10376_),
    .B(_10384_),
    .Y(_03442_));
 NOR2x1_ASAP7_75t_R _29385_ (.A(_00462_),
    .B(_10376_),
    .Y(_10385_));
 AO21x1_ASAP7_75t_R _29386_ (.A1(_07581_),
    .A2(_10376_),
    .B(_10385_),
    .Y(_03443_));
 NOR2x1_ASAP7_75t_R _29387_ (.A(_00492_),
    .B(_10376_),
    .Y(_10386_));
 AO21x1_ASAP7_75t_R _29388_ (.A1(_07620_),
    .A2(_10376_),
    .B(_10386_),
    .Y(_03444_));
 NOR2x1_ASAP7_75t_R _29389_ (.A(_00522_),
    .B(_10376_),
    .Y(_10387_));
 AO21x1_ASAP7_75t_R _29390_ (.A1(_07676_),
    .A2(_10376_),
    .B(_10387_),
    .Y(_03445_));
 TAPCELL_ASAP7_75t_R PHY_405 ();
 NOR2x1_ASAP7_75t_R _29392_ (.A(_00552_),
    .B(_10376_),
    .Y(_10389_));
 AO21x1_ASAP7_75t_R _29393_ (.A1(_07738_),
    .A2(_10376_),
    .B(_10389_),
    .Y(_03446_));
 NOR2x1_ASAP7_75t_R _29394_ (.A(_00582_),
    .B(_10376_),
    .Y(_10390_));
 AO21x1_ASAP7_75t_R _29395_ (.A1(_07780_),
    .A2(_10376_),
    .B(_10390_),
    .Y(_03447_));
 TAPCELL_ASAP7_75t_R PHY_404 ();
 NOR2x1_ASAP7_75t_R _29397_ (.A(_00612_),
    .B(_10376_),
    .Y(_10392_));
 AO21x1_ASAP7_75t_R _29398_ (.A1(_07817_),
    .A2(_10376_),
    .B(_10392_),
    .Y(_03448_));
 NOR2x1_ASAP7_75t_R _29399_ (.A(_00642_),
    .B(_10376_),
    .Y(_10393_));
 AO21x1_ASAP7_75t_R _29400_ (.A1(_07865_),
    .A2(_10376_),
    .B(_10393_),
    .Y(_03449_));
 NOR2x1_ASAP7_75t_R _29401_ (.A(_00341_),
    .B(_10376_),
    .Y(_10394_));
 AO21x1_ASAP7_75t_R _29402_ (.A1(_07908_),
    .A2(_10376_),
    .B(_10394_),
    .Y(_03450_));
 NOR2x1_ASAP7_75t_R _29403_ (.A(_00704_),
    .B(_10376_),
    .Y(_10395_));
 AO21x1_ASAP7_75t_R _29404_ (.A1(_07950_),
    .A2(_10376_),
    .B(_10395_),
    .Y(_03451_));
 NOR2x1_ASAP7_75t_R _29405_ (.A(_00736_),
    .B(_10376_),
    .Y(_10396_));
 AO21x1_ASAP7_75t_R _29406_ (.A1(_07990_),
    .A2(_10376_),
    .B(_10396_),
    .Y(_03452_));
 NOR2x1_ASAP7_75t_R _29407_ (.A(_00769_),
    .B(_10376_),
    .Y(_10397_));
 AO21x1_ASAP7_75t_R _29408_ (.A1(_08034_),
    .A2(_10376_),
    .B(_10397_),
    .Y(_03453_));
 NOR2x1_ASAP7_75t_R _29409_ (.A(_00802_),
    .B(_10376_),
    .Y(_10398_));
 AO21x1_ASAP7_75t_R _29410_ (.A1(_08073_),
    .A2(_10376_),
    .B(_10398_),
    .Y(_03454_));
 NOR2x1_ASAP7_75t_R _29411_ (.A(_00835_),
    .B(_10376_),
    .Y(_10399_));
 AO21x1_ASAP7_75t_R _29412_ (.A1(_08116_),
    .A2(_10376_),
    .B(_10399_),
    .Y(_03455_));
 TAPCELL_ASAP7_75t_R PHY_403 ();
 NOR2x1_ASAP7_75t_R _29414_ (.A(_00867_),
    .B(_10376_),
    .Y(_10401_));
 AO21x1_ASAP7_75t_R _29415_ (.A1(net251),
    .A2(_10376_),
    .B(_10401_),
    .Y(_03456_));
 NOR2x1_ASAP7_75t_R _29416_ (.A(_00900_),
    .B(_10376_),
    .Y(_10402_));
 AO21x1_ASAP7_75t_R _29417_ (.A1(_08187_),
    .A2(_10376_),
    .B(_10402_),
    .Y(_03457_));
 TAPCELL_ASAP7_75t_R PHY_402 ();
 NOR2x1_ASAP7_75t_R _29419_ (.A(_00932_),
    .B(_10376_),
    .Y(_10404_));
 AO21x1_ASAP7_75t_R _29420_ (.A1(_08219_),
    .A2(_10376_),
    .B(_10404_),
    .Y(_03458_));
 NOR2x1_ASAP7_75t_R _29421_ (.A(_00965_),
    .B(_10376_),
    .Y(_10405_));
 AO21x1_ASAP7_75t_R _29422_ (.A1(_08254_),
    .A2(_10376_),
    .B(_10405_),
    .Y(_03459_));
 NOR2x1_ASAP7_75t_R _29423_ (.A(_00997_),
    .B(_10376_),
    .Y(_10406_));
 AO21x1_ASAP7_75t_R _29424_ (.A1(net250),
    .A2(_10376_),
    .B(_10406_),
    .Y(_03460_));
 NOR2x1_ASAP7_75t_R _29425_ (.A(_01031_),
    .B(_10376_),
    .Y(_10407_));
 AO21x1_ASAP7_75t_R _29426_ (.A1(_08319_),
    .A2(_10376_),
    .B(_10407_),
    .Y(_03461_));
 NOR2x1_ASAP7_75t_R _29427_ (.A(_01063_),
    .B(_10376_),
    .Y(_10408_));
 AO21x1_ASAP7_75t_R _29428_ (.A1(_08357_),
    .A2(_10376_),
    .B(_10408_),
    .Y(_03462_));
 NOR2x1_ASAP7_75t_R _29429_ (.A(_01096_),
    .B(_10376_),
    .Y(_10409_));
 AO21x1_ASAP7_75t_R _29430_ (.A1(_08388_),
    .A2(_10376_),
    .B(_10409_),
    .Y(_03463_));
 NOR2x1_ASAP7_75t_R _29431_ (.A(_01128_),
    .B(_10376_),
    .Y(_10410_));
 AO21x1_ASAP7_75t_R _29432_ (.A1(_08419_),
    .A2(_10376_),
    .B(_10410_),
    .Y(_03464_));
 NOR2x1_ASAP7_75t_R _29433_ (.A(_01162_),
    .B(_10376_),
    .Y(_10411_));
 AO21x1_ASAP7_75t_R _29434_ (.A1(_08451_),
    .A2(_10376_),
    .B(_10411_),
    .Y(_03465_));
 NOR2x1_ASAP7_75t_R _29435_ (.A(_01194_),
    .B(_10376_),
    .Y(_10412_));
 AO21x1_ASAP7_75t_R _29436_ (.A1(_08481_),
    .A2(_10376_),
    .B(_10412_),
    .Y(_03466_));
 NOR2x1_ASAP7_75t_R _29437_ (.A(_01228_),
    .B(_10376_),
    .Y(_10413_));
 AO21x1_ASAP7_75t_R _29438_ (.A1(_08512_),
    .A2(_10376_),
    .B(_10413_),
    .Y(_03467_));
 NOR2x1_ASAP7_75t_R _29439_ (.A(_01260_),
    .B(_10376_),
    .Y(_10414_));
 AO21x1_ASAP7_75t_R _29440_ (.A1(_08545_),
    .A2(_10376_),
    .B(_10414_),
    .Y(_03468_));
 NOR2x1_ASAP7_75t_R _29441_ (.A(_01294_),
    .B(_10376_),
    .Y(_10415_));
 AO21x1_ASAP7_75t_R _29442_ (.A1(_08573_),
    .A2(_10376_),
    .B(_10415_),
    .Y(_03469_));
 AND3x4_ASAP7_75t_R _29443_ (.A(_06881_),
    .B(_09736_),
    .C(_10334_),
    .Y(_10416_));
 TAPCELL_ASAP7_75t_R PHY_401 ();
 TAPCELL_ASAP7_75t_R PHY_400 ();
 TAPCELL_ASAP7_75t_R PHY_399 ();
 NOR2x1_ASAP7_75t_R _29447_ (.A(_00310_),
    .B(_10416_),
    .Y(_10420_));
 AO21x1_ASAP7_75t_R _29448_ (.A1(_07180_),
    .A2(_10416_),
    .B(_10420_),
    .Y(_03470_));
 NOR2x1_ASAP7_75t_R _29449_ (.A(_00264_),
    .B(_10416_),
    .Y(_10421_));
 AO21x1_ASAP7_75t_R _29450_ (.A1(_07313_),
    .A2(_10416_),
    .B(_10421_),
    .Y(_03471_));
 NOR2x1_ASAP7_75t_R _29451_ (.A(_00372_),
    .B(_10416_),
    .Y(_10422_));
 AO21x1_ASAP7_75t_R _29452_ (.A1(_07398_),
    .A2(_10416_),
    .B(_10422_),
    .Y(_03472_));
 NOR2x1_ASAP7_75t_R _29453_ (.A(_00403_),
    .B(_10416_),
    .Y(_10423_));
 AO21x1_ASAP7_75t_R _29454_ (.A1(_07469_),
    .A2(_10416_),
    .B(_10423_),
    .Y(_03473_));
 NOR2x1_ASAP7_75t_R _29455_ (.A(_00433_),
    .B(_10416_),
    .Y(_10424_));
 AO21x1_ASAP7_75t_R _29456_ (.A1(_07534_),
    .A2(_10416_),
    .B(_10424_),
    .Y(_03474_));
 NOR2x1_ASAP7_75t_R _29457_ (.A(_00463_),
    .B(_10416_),
    .Y(_10425_));
 AO21x1_ASAP7_75t_R _29458_ (.A1(_07581_),
    .A2(_10416_),
    .B(_10425_),
    .Y(_03475_));
 NOR2x1_ASAP7_75t_R _29459_ (.A(_00493_),
    .B(_10416_),
    .Y(_10426_));
 AO21x1_ASAP7_75t_R _29460_ (.A1(net253),
    .A2(_10416_),
    .B(_10426_),
    .Y(_03476_));
 NOR2x1_ASAP7_75t_R _29461_ (.A(_00523_),
    .B(_10416_),
    .Y(_10427_));
 AO21x1_ASAP7_75t_R _29462_ (.A1(_07676_),
    .A2(_10416_),
    .B(_10427_),
    .Y(_03477_));
 TAPCELL_ASAP7_75t_R PHY_398 ();
 NOR2x1_ASAP7_75t_R _29464_ (.A(_00553_),
    .B(_10416_),
    .Y(_10429_));
 AO21x1_ASAP7_75t_R _29465_ (.A1(net252),
    .A2(_10416_),
    .B(_10429_),
    .Y(_03478_));
 NOR2x1_ASAP7_75t_R _29466_ (.A(_00583_),
    .B(_10416_),
    .Y(_10430_));
 AO21x1_ASAP7_75t_R _29467_ (.A1(_07780_),
    .A2(_10416_),
    .B(_10430_),
    .Y(_03479_));
 TAPCELL_ASAP7_75t_R PHY_397 ();
 NOR2x1_ASAP7_75t_R _29469_ (.A(_00613_),
    .B(_10416_),
    .Y(_10432_));
 AO21x1_ASAP7_75t_R _29470_ (.A1(_07817_),
    .A2(_10416_),
    .B(_10432_),
    .Y(_03480_));
 NOR2x1_ASAP7_75t_R _29471_ (.A(_00643_),
    .B(_10416_),
    .Y(_10433_));
 AO21x1_ASAP7_75t_R _29472_ (.A1(_07865_),
    .A2(_10416_),
    .B(_10433_),
    .Y(_03481_));
 NOR2x1_ASAP7_75t_R _29473_ (.A(_00342_),
    .B(_10416_),
    .Y(_10434_));
 AO21x1_ASAP7_75t_R _29474_ (.A1(_07908_),
    .A2(_10416_),
    .B(_10434_),
    .Y(_03482_));
 NOR2x1_ASAP7_75t_R _29475_ (.A(_00705_),
    .B(_10416_),
    .Y(_10435_));
 AO21x1_ASAP7_75t_R _29476_ (.A1(_07950_),
    .A2(_10416_),
    .B(_10435_),
    .Y(_03483_));
 NOR2x1_ASAP7_75t_R _29477_ (.A(_00737_),
    .B(_10416_),
    .Y(_10436_));
 AO21x1_ASAP7_75t_R _29478_ (.A1(_07990_),
    .A2(_10416_),
    .B(_10436_),
    .Y(_03484_));
 NOR2x1_ASAP7_75t_R _29479_ (.A(_00770_),
    .B(_10416_),
    .Y(_10437_));
 AO21x1_ASAP7_75t_R _29480_ (.A1(_08034_),
    .A2(_10416_),
    .B(_10437_),
    .Y(_03485_));
 NOR2x1_ASAP7_75t_R _29481_ (.A(_00803_),
    .B(_10416_),
    .Y(_10438_));
 AO21x1_ASAP7_75t_R _29482_ (.A1(_08073_),
    .A2(_10416_),
    .B(_10438_),
    .Y(_03486_));
 NOR2x1_ASAP7_75t_R _29483_ (.A(_00836_),
    .B(_10416_),
    .Y(_10439_));
 AO21x1_ASAP7_75t_R _29484_ (.A1(_08116_),
    .A2(_10416_),
    .B(_10439_),
    .Y(_03487_));
 TAPCELL_ASAP7_75t_R PHY_396 ();
 NOR2x1_ASAP7_75t_R _29486_ (.A(_00868_),
    .B(_10416_),
    .Y(_10441_));
 AO21x1_ASAP7_75t_R _29487_ (.A1(net251),
    .A2(_10416_),
    .B(_10441_),
    .Y(_03488_));
 NOR2x1_ASAP7_75t_R _29488_ (.A(_00901_),
    .B(_10416_),
    .Y(_10442_));
 AO21x1_ASAP7_75t_R _29489_ (.A1(_08187_),
    .A2(_10416_),
    .B(_10442_),
    .Y(_03489_));
 TAPCELL_ASAP7_75t_R PHY_395 ();
 NOR2x1_ASAP7_75t_R _29491_ (.A(_00933_),
    .B(_10416_),
    .Y(_10444_));
 AO21x1_ASAP7_75t_R _29492_ (.A1(_08219_),
    .A2(_10416_),
    .B(_10444_),
    .Y(_03490_));
 NOR2x1_ASAP7_75t_R _29493_ (.A(_00966_),
    .B(_10416_),
    .Y(_10445_));
 AO21x1_ASAP7_75t_R _29494_ (.A1(_08254_),
    .A2(_10416_),
    .B(_10445_),
    .Y(_03491_));
 NOR2x1_ASAP7_75t_R _29495_ (.A(_00998_),
    .B(_10416_),
    .Y(_10446_));
 AO21x1_ASAP7_75t_R _29496_ (.A1(net250),
    .A2(_10416_),
    .B(_10446_),
    .Y(_03492_));
 NOR2x1_ASAP7_75t_R _29497_ (.A(_01032_),
    .B(_10416_),
    .Y(_10447_));
 AO21x1_ASAP7_75t_R _29498_ (.A1(_08319_),
    .A2(_10416_),
    .B(_10447_),
    .Y(_03493_));
 NOR2x1_ASAP7_75t_R _29499_ (.A(_01064_),
    .B(_10416_),
    .Y(_10448_));
 AO21x1_ASAP7_75t_R _29500_ (.A1(_08357_),
    .A2(_10416_),
    .B(_10448_),
    .Y(_03494_));
 NOR2x1_ASAP7_75t_R _29501_ (.A(_01097_),
    .B(_10416_),
    .Y(_10449_));
 AO21x1_ASAP7_75t_R _29502_ (.A1(_08388_),
    .A2(_10416_),
    .B(_10449_),
    .Y(_03495_));
 NOR2x1_ASAP7_75t_R _29503_ (.A(_01129_),
    .B(_10416_),
    .Y(_10450_));
 AO21x1_ASAP7_75t_R _29504_ (.A1(_08419_),
    .A2(_10416_),
    .B(_10450_),
    .Y(_03496_));
 NOR2x1_ASAP7_75t_R _29505_ (.A(_01163_),
    .B(_10416_),
    .Y(_10451_));
 AO21x1_ASAP7_75t_R _29506_ (.A1(_08451_),
    .A2(_10416_),
    .B(_10451_),
    .Y(_03497_));
 NOR2x1_ASAP7_75t_R _29507_ (.A(_01195_),
    .B(_10416_),
    .Y(_10452_));
 AO21x1_ASAP7_75t_R _29508_ (.A1(_08481_),
    .A2(_10416_),
    .B(_10452_),
    .Y(_03498_));
 NOR2x1_ASAP7_75t_R _29509_ (.A(_01229_),
    .B(_10416_),
    .Y(_10453_));
 AO21x1_ASAP7_75t_R _29510_ (.A1(_08512_),
    .A2(_10416_),
    .B(_10453_),
    .Y(_03499_));
 NOR2x1_ASAP7_75t_R _29511_ (.A(_01261_),
    .B(_10416_),
    .Y(_10454_));
 AO21x1_ASAP7_75t_R _29512_ (.A1(_08545_),
    .A2(_10416_),
    .B(_10454_),
    .Y(_03500_));
 NOR2x1_ASAP7_75t_R _29513_ (.A(_01295_),
    .B(_10416_),
    .Y(_10455_));
 AO21x1_ASAP7_75t_R _29514_ (.A1(_08573_),
    .A2(_10416_),
    .B(_10455_),
    .Y(_03501_));
 AND4x2_ASAP7_75t_R _29515_ (.A(_00323_),
    .B(_00184_),
    .C(_09779_),
    .D(_10334_),
    .Y(_10456_));
 TAPCELL_ASAP7_75t_R PHY_394 ();
 TAPCELL_ASAP7_75t_R PHY_393 ();
 TAPCELL_ASAP7_75t_R PHY_392 ();
 NOR2x1_ASAP7_75t_R _29519_ (.A(_00311_),
    .B(_10456_),
    .Y(_10460_));
 AO21x1_ASAP7_75t_R _29520_ (.A1(_07180_),
    .A2(_10456_),
    .B(_10460_),
    .Y(_03502_));
 NOR2x1_ASAP7_75t_R _29521_ (.A(_00265_),
    .B(_10456_),
    .Y(_10461_));
 AO21x1_ASAP7_75t_R _29522_ (.A1(_07313_),
    .A2(_10456_),
    .B(_10461_),
    .Y(_03503_));
 NOR2x1_ASAP7_75t_R _29523_ (.A(_00373_),
    .B(_10456_),
    .Y(_10462_));
 AO21x1_ASAP7_75t_R _29524_ (.A1(_07398_),
    .A2(net263),
    .B(_10462_),
    .Y(_03504_));
 NOR2x1_ASAP7_75t_R _29525_ (.A(_00404_),
    .B(net263),
    .Y(_10463_));
 AO21x1_ASAP7_75t_R _29526_ (.A1(_07469_),
    .A2(net263),
    .B(_10463_),
    .Y(_03505_));
 NOR2x1_ASAP7_75t_R _29527_ (.A(_00434_),
    .B(_10456_),
    .Y(_10464_));
 AO21x1_ASAP7_75t_R _29528_ (.A1(_07534_),
    .A2(_10456_),
    .B(_10464_),
    .Y(_03506_));
 NOR2x1_ASAP7_75t_R _29529_ (.A(_00464_),
    .B(net263),
    .Y(_10465_));
 AO21x1_ASAP7_75t_R _29530_ (.A1(_07581_),
    .A2(net263),
    .B(_10465_),
    .Y(_03507_));
 NOR2x1_ASAP7_75t_R _29531_ (.A(_00494_),
    .B(_10456_),
    .Y(_10466_));
 AO21x1_ASAP7_75t_R _29532_ (.A1(net253),
    .A2(_10456_),
    .B(_10466_),
    .Y(_03508_));
 NOR2x1_ASAP7_75t_R _29533_ (.A(_00524_),
    .B(net263),
    .Y(_10467_));
 AO21x1_ASAP7_75t_R _29534_ (.A1(_07676_),
    .A2(net263),
    .B(_10467_),
    .Y(_03509_));
 TAPCELL_ASAP7_75t_R PHY_391 ();
 NOR2x1_ASAP7_75t_R _29536_ (.A(_00554_),
    .B(_10456_),
    .Y(_10469_));
 AO21x1_ASAP7_75t_R _29537_ (.A1(_07738_),
    .A2(_10456_),
    .B(_10469_),
    .Y(_03510_));
 NOR2x1_ASAP7_75t_R _29538_ (.A(_00584_),
    .B(_10456_),
    .Y(_10470_));
 AO21x1_ASAP7_75t_R _29539_ (.A1(_07780_),
    .A2(_10456_),
    .B(_10470_),
    .Y(_03511_));
 TAPCELL_ASAP7_75t_R PHY_390 ();
 NOR2x1_ASAP7_75t_R _29541_ (.A(_00614_),
    .B(net263),
    .Y(_10472_));
 AO21x1_ASAP7_75t_R _29542_ (.A1(_07817_),
    .A2(net263),
    .B(_10472_),
    .Y(_03512_));
 NOR2x1_ASAP7_75t_R _29543_ (.A(_00644_),
    .B(_10456_),
    .Y(_10473_));
 AO21x1_ASAP7_75t_R _29544_ (.A1(_07865_),
    .A2(_10456_),
    .B(_10473_),
    .Y(_03513_));
 NOR2x1_ASAP7_75t_R _29545_ (.A(_00343_),
    .B(_10456_),
    .Y(_10474_));
 AO21x1_ASAP7_75t_R _29546_ (.A1(_07908_),
    .A2(_10456_),
    .B(_10474_),
    .Y(_03514_));
 NOR2x1_ASAP7_75t_R _29547_ (.A(_00706_),
    .B(net262),
    .Y(_10475_));
 AO21x1_ASAP7_75t_R _29548_ (.A1(_07950_),
    .A2(net262),
    .B(_10475_),
    .Y(_03515_));
 NOR2x1_ASAP7_75t_R _29549_ (.A(_00738_),
    .B(_10456_),
    .Y(_10476_));
 AO21x1_ASAP7_75t_R _29550_ (.A1(_07990_),
    .A2(_10456_),
    .B(_10476_),
    .Y(_03516_));
 NOR2x1_ASAP7_75t_R _29551_ (.A(_00771_),
    .B(net262),
    .Y(_10477_));
 AO21x1_ASAP7_75t_R _29552_ (.A1(_08034_),
    .A2(net262),
    .B(_10477_),
    .Y(_03517_));
 NOR2x1_ASAP7_75t_R _29553_ (.A(_00804_),
    .B(net262),
    .Y(_10478_));
 AO21x1_ASAP7_75t_R _29554_ (.A1(_08073_),
    .A2(net262),
    .B(_10478_),
    .Y(_03518_));
 NOR2x1_ASAP7_75t_R _29555_ (.A(_00837_),
    .B(net263),
    .Y(_10479_));
 AO21x1_ASAP7_75t_R _29556_ (.A1(_08116_),
    .A2(net263),
    .B(_10479_),
    .Y(_03519_));
 TAPCELL_ASAP7_75t_R PHY_389 ();
 NOR2x1_ASAP7_75t_R _29558_ (.A(_00869_),
    .B(net262),
    .Y(_10481_));
 AO21x1_ASAP7_75t_R _29559_ (.A1(net251),
    .A2(net262),
    .B(_10481_),
    .Y(_03520_));
 NOR2x1_ASAP7_75t_R _29560_ (.A(_00902_),
    .B(net262),
    .Y(_10482_));
 AO21x1_ASAP7_75t_R _29561_ (.A1(_08187_),
    .A2(net262),
    .B(_10482_),
    .Y(_03521_));
 TAPCELL_ASAP7_75t_R PHY_388 ();
 NOR2x1_ASAP7_75t_R _29563_ (.A(_00934_),
    .B(net263),
    .Y(_10484_));
 AO21x1_ASAP7_75t_R _29564_ (.A1(_08219_),
    .A2(net263),
    .B(_10484_),
    .Y(_03522_));
 NOR2x1_ASAP7_75t_R _29565_ (.A(_00967_),
    .B(net262),
    .Y(_10485_));
 AO21x1_ASAP7_75t_R _29566_ (.A1(_08254_),
    .A2(net262),
    .B(_10485_),
    .Y(_03523_));
 NOR2x1_ASAP7_75t_R _29567_ (.A(_00999_),
    .B(_10456_),
    .Y(_10486_));
 AO21x1_ASAP7_75t_R _29568_ (.A1(net250),
    .A2(_10456_),
    .B(_10486_),
    .Y(_03524_));
 NOR2x1_ASAP7_75t_R _29569_ (.A(_01033_),
    .B(net263),
    .Y(_10487_));
 AO21x1_ASAP7_75t_R _29570_ (.A1(_08319_),
    .A2(net263),
    .B(_10487_),
    .Y(_03525_));
 NOR2x1_ASAP7_75t_R _29571_ (.A(_01065_),
    .B(net262),
    .Y(_10488_));
 AO21x1_ASAP7_75t_R _29572_ (.A1(_08357_),
    .A2(net262),
    .B(_10488_),
    .Y(_03526_));
 NOR2x1_ASAP7_75t_R _29573_ (.A(_01098_),
    .B(net262),
    .Y(_10489_));
 AO21x1_ASAP7_75t_R _29574_ (.A1(_08388_),
    .A2(net262),
    .B(_10489_),
    .Y(_03527_));
 NOR2x1_ASAP7_75t_R _29575_ (.A(_01130_),
    .B(net262),
    .Y(_10490_));
 AO21x1_ASAP7_75t_R _29576_ (.A1(_08419_),
    .A2(net262),
    .B(_10490_),
    .Y(_03528_));
 NOR2x1_ASAP7_75t_R _29577_ (.A(_01164_),
    .B(net262),
    .Y(_10491_));
 AO21x1_ASAP7_75t_R _29578_ (.A1(_08451_),
    .A2(net262),
    .B(_10491_),
    .Y(_03529_));
 NOR2x1_ASAP7_75t_R _29579_ (.A(_01196_),
    .B(_10456_),
    .Y(_10492_));
 AO21x1_ASAP7_75t_R _29580_ (.A1(_08481_),
    .A2(_10456_),
    .B(_10492_),
    .Y(_03530_));
 NOR2x1_ASAP7_75t_R _29581_ (.A(_01230_),
    .B(net263),
    .Y(_10493_));
 AO21x1_ASAP7_75t_R _29582_ (.A1(_08512_),
    .A2(net263),
    .B(_10493_),
    .Y(_03531_));
 NOR2x1_ASAP7_75t_R _29583_ (.A(_01262_),
    .B(net262),
    .Y(_10494_));
 AO21x1_ASAP7_75t_R _29584_ (.A1(_08545_),
    .A2(net262),
    .B(_10494_),
    .Y(_03532_));
 NOR2x1_ASAP7_75t_R _29585_ (.A(_01296_),
    .B(_10456_),
    .Y(_10495_));
 AO21x1_ASAP7_75t_R _29586_ (.A1(_08573_),
    .A2(_10456_),
    .B(_10495_),
    .Y(_03533_));
 AND3x4_ASAP7_75t_R _29587_ (.A(_06882_),
    .B(_09779_),
    .C(_10334_),
    .Y(_10496_));
 TAPCELL_ASAP7_75t_R PHY_387 ();
 TAPCELL_ASAP7_75t_R PHY_386 ();
 TAPCELL_ASAP7_75t_R PHY_385 ();
 NOR2x1_ASAP7_75t_R _29591_ (.A(_00312_),
    .B(_10496_),
    .Y(_10500_));
 AO21x1_ASAP7_75t_R _29592_ (.A1(_07180_),
    .A2(_10496_),
    .B(_10500_),
    .Y(_03534_));
 NOR2x1_ASAP7_75t_R _29593_ (.A(_00266_),
    .B(_10496_),
    .Y(_10501_));
 AO21x1_ASAP7_75t_R _29594_ (.A1(_07313_),
    .A2(_10496_),
    .B(_10501_),
    .Y(_03535_));
 NOR2x1_ASAP7_75t_R _29595_ (.A(_00374_),
    .B(_10496_),
    .Y(_10502_));
 AO21x1_ASAP7_75t_R _29596_ (.A1(_07398_),
    .A2(_10496_),
    .B(_10502_),
    .Y(_03536_));
 NOR2x1_ASAP7_75t_R _29597_ (.A(_00405_),
    .B(_10496_),
    .Y(_10503_));
 AO21x1_ASAP7_75t_R _29598_ (.A1(_07469_),
    .A2(_10496_),
    .B(_10503_),
    .Y(_03537_));
 NOR2x1_ASAP7_75t_R _29599_ (.A(_00435_),
    .B(_10496_),
    .Y(_10504_));
 AO21x1_ASAP7_75t_R _29600_ (.A1(_07534_),
    .A2(_10496_),
    .B(_10504_),
    .Y(_03538_));
 NOR2x1_ASAP7_75t_R _29601_ (.A(_00465_),
    .B(_10496_),
    .Y(_10505_));
 AO21x1_ASAP7_75t_R _29602_ (.A1(_07581_),
    .A2(_10496_),
    .B(_10505_),
    .Y(_03539_));
 NOR2x1_ASAP7_75t_R _29603_ (.A(_00495_),
    .B(_10496_),
    .Y(_10506_));
 AO21x1_ASAP7_75t_R _29604_ (.A1(net253),
    .A2(_10496_),
    .B(_10506_),
    .Y(_03540_));
 NOR2x1_ASAP7_75t_R _29605_ (.A(_00525_),
    .B(_10496_),
    .Y(_10507_));
 AO21x1_ASAP7_75t_R _29606_ (.A1(_07676_),
    .A2(_10496_),
    .B(_10507_),
    .Y(_03541_));
 TAPCELL_ASAP7_75t_R PHY_384 ();
 NOR2x1_ASAP7_75t_R _29608_ (.A(_00555_),
    .B(_10496_),
    .Y(_10509_));
 AO21x1_ASAP7_75t_R _29609_ (.A1(net252),
    .A2(_10496_),
    .B(_10509_),
    .Y(_03542_));
 NOR2x1_ASAP7_75t_R _29610_ (.A(_00585_),
    .B(_10496_),
    .Y(_10510_));
 AO21x1_ASAP7_75t_R _29611_ (.A1(_07780_),
    .A2(_10496_),
    .B(_10510_),
    .Y(_03543_));
 TAPCELL_ASAP7_75t_R PHY_383 ();
 NOR2x1_ASAP7_75t_R _29613_ (.A(_00615_),
    .B(_10496_),
    .Y(_10512_));
 AO21x1_ASAP7_75t_R _29614_ (.A1(_07817_),
    .A2(_10496_),
    .B(_10512_),
    .Y(_03544_));
 NOR2x1_ASAP7_75t_R _29615_ (.A(_00645_),
    .B(_10496_),
    .Y(_10513_));
 AO21x1_ASAP7_75t_R _29616_ (.A1(_07865_),
    .A2(_10496_),
    .B(_10513_),
    .Y(_03545_));
 NOR2x1_ASAP7_75t_R _29617_ (.A(_00344_),
    .B(_10496_),
    .Y(_10514_));
 AO21x1_ASAP7_75t_R _29618_ (.A1(_07908_),
    .A2(_10496_),
    .B(_10514_),
    .Y(_03546_));
 NOR2x1_ASAP7_75t_R _29619_ (.A(_00707_),
    .B(_10496_),
    .Y(_10515_));
 AO21x1_ASAP7_75t_R _29620_ (.A1(_07950_),
    .A2(_10496_),
    .B(_10515_),
    .Y(_03547_));
 NOR2x1_ASAP7_75t_R _29621_ (.A(_00739_),
    .B(_10496_),
    .Y(_10516_));
 AO21x1_ASAP7_75t_R _29622_ (.A1(_07990_),
    .A2(_10496_),
    .B(_10516_),
    .Y(_03548_));
 NOR2x1_ASAP7_75t_R _29623_ (.A(_00772_),
    .B(_10496_),
    .Y(_10517_));
 AO21x1_ASAP7_75t_R _29624_ (.A1(_08034_),
    .A2(_10496_),
    .B(_10517_),
    .Y(_03549_));
 NOR2x1_ASAP7_75t_R _29625_ (.A(_00805_),
    .B(_10496_),
    .Y(_10518_));
 AO21x1_ASAP7_75t_R _29626_ (.A1(_08073_),
    .A2(_10496_),
    .B(_10518_),
    .Y(_03550_));
 NOR2x1_ASAP7_75t_R _29627_ (.A(_00838_),
    .B(_10496_),
    .Y(_10519_));
 AO21x1_ASAP7_75t_R _29628_ (.A1(_08116_),
    .A2(_10496_),
    .B(_10519_),
    .Y(_03551_));
 TAPCELL_ASAP7_75t_R PHY_382 ();
 NOR2x1_ASAP7_75t_R _29630_ (.A(_00870_),
    .B(_10496_),
    .Y(_10521_));
 AO21x1_ASAP7_75t_R _29631_ (.A1(net251),
    .A2(_10496_),
    .B(_10521_),
    .Y(_03552_));
 NOR2x1_ASAP7_75t_R _29632_ (.A(_00903_),
    .B(_10496_),
    .Y(_10522_));
 AO21x1_ASAP7_75t_R _29633_ (.A1(_08187_),
    .A2(_10496_),
    .B(_10522_),
    .Y(_03553_));
 TAPCELL_ASAP7_75t_R PHY_381 ();
 NOR2x1_ASAP7_75t_R _29635_ (.A(_00935_),
    .B(_10496_),
    .Y(_10524_));
 AO21x1_ASAP7_75t_R _29636_ (.A1(_08219_),
    .A2(_10496_),
    .B(_10524_),
    .Y(_03554_));
 NOR2x1_ASAP7_75t_R _29637_ (.A(_00968_),
    .B(_10496_),
    .Y(_10525_));
 AO21x1_ASAP7_75t_R _29638_ (.A1(_08254_),
    .A2(_10496_),
    .B(_10525_),
    .Y(_03555_));
 NOR2x1_ASAP7_75t_R _29639_ (.A(_01000_),
    .B(_10496_),
    .Y(_10526_));
 AO21x1_ASAP7_75t_R _29640_ (.A1(net250),
    .A2(_10496_),
    .B(_10526_),
    .Y(_03556_));
 NOR2x1_ASAP7_75t_R _29641_ (.A(_01034_),
    .B(_10496_),
    .Y(_10527_));
 AO21x1_ASAP7_75t_R _29642_ (.A1(_08319_),
    .A2(_10496_),
    .B(_10527_),
    .Y(_03557_));
 NOR2x1_ASAP7_75t_R _29643_ (.A(_01066_),
    .B(_10496_),
    .Y(_10528_));
 AO21x1_ASAP7_75t_R _29644_ (.A1(_08357_),
    .A2(_10496_),
    .B(_10528_),
    .Y(_03558_));
 NOR2x1_ASAP7_75t_R _29645_ (.A(_01099_),
    .B(_10496_),
    .Y(_10529_));
 AO21x1_ASAP7_75t_R _29646_ (.A1(_08388_),
    .A2(_10496_),
    .B(_10529_),
    .Y(_03559_));
 NOR2x1_ASAP7_75t_R _29647_ (.A(_01131_),
    .B(_10496_),
    .Y(_10530_));
 AO21x1_ASAP7_75t_R _29648_ (.A1(_08419_),
    .A2(_10496_),
    .B(_10530_),
    .Y(_03560_));
 NOR2x1_ASAP7_75t_R _29649_ (.A(_01165_),
    .B(_10496_),
    .Y(_10531_));
 AO21x1_ASAP7_75t_R _29650_ (.A1(_08451_),
    .A2(_10496_),
    .B(_10531_),
    .Y(_03561_));
 NOR2x1_ASAP7_75t_R _29651_ (.A(_01197_),
    .B(_10496_),
    .Y(_10532_));
 AO21x1_ASAP7_75t_R _29652_ (.A1(_08481_),
    .A2(_10496_),
    .B(_10532_),
    .Y(_03562_));
 NOR2x1_ASAP7_75t_R _29653_ (.A(_01231_),
    .B(_10496_),
    .Y(_10533_));
 AO21x1_ASAP7_75t_R _29654_ (.A1(_08512_),
    .A2(_10496_),
    .B(_10533_),
    .Y(_03563_));
 NOR2x1_ASAP7_75t_R _29655_ (.A(_01263_),
    .B(_10496_),
    .Y(_10534_));
 AO21x1_ASAP7_75t_R _29656_ (.A1(_08545_),
    .A2(_10496_),
    .B(_10534_),
    .Y(_03564_));
 NOR2x1_ASAP7_75t_R _29657_ (.A(_01297_),
    .B(_10496_),
    .Y(_10535_));
 AO21x1_ASAP7_75t_R _29658_ (.A1(_08573_),
    .A2(_10496_),
    .B(_10535_),
    .Y(_03565_));
 TAPCELL_ASAP7_75t_R PHY_380 ();
 AND3x4_ASAP7_75t_R _29660_ (.A(_09663_),
    .B(_09779_),
    .C(_10334_),
    .Y(_10537_));
 TAPCELL_ASAP7_75t_R PHY_379 ();
 TAPCELL_ASAP7_75t_R PHY_378 ();
 TAPCELL_ASAP7_75t_R PHY_377 ();
 NOR2x1_ASAP7_75t_R _29664_ (.A(_00313_),
    .B(_10537_),
    .Y(_10541_));
 AO21x1_ASAP7_75t_R _29665_ (.A1(_07180_),
    .A2(_10537_),
    .B(_10541_),
    .Y(_03566_));
 TAPCELL_ASAP7_75t_R PHY_376 ();
 NOR2x1_ASAP7_75t_R _29667_ (.A(_00267_),
    .B(_10537_),
    .Y(_10543_));
 AO21x1_ASAP7_75t_R _29668_ (.A1(_07313_),
    .A2(_10537_),
    .B(_10543_),
    .Y(_03567_));
 TAPCELL_ASAP7_75t_R PHY_375 ();
 NOR2x1_ASAP7_75t_R _29670_ (.A(_00375_),
    .B(_10537_),
    .Y(_10545_));
 AO21x1_ASAP7_75t_R _29671_ (.A1(_07398_),
    .A2(_10537_),
    .B(_10545_),
    .Y(_03568_));
 TAPCELL_ASAP7_75t_R PHY_374 ();
 NOR2x1_ASAP7_75t_R _29673_ (.A(_00406_),
    .B(_10537_),
    .Y(_10547_));
 AO21x1_ASAP7_75t_R _29674_ (.A1(_07469_),
    .A2(_10537_),
    .B(_10547_),
    .Y(_03569_));
 TAPCELL_ASAP7_75t_R PHY_373 ();
 NOR2x1_ASAP7_75t_R _29676_ (.A(_00436_),
    .B(_10537_),
    .Y(_10549_));
 AO21x1_ASAP7_75t_R _29677_ (.A1(_07534_),
    .A2(_10537_),
    .B(_10549_),
    .Y(_03570_));
 TAPCELL_ASAP7_75t_R PHY_372 ();
 NOR2x1_ASAP7_75t_R _29679_ (.A(_00466_),
    .B(_10537_),
    .Y(_10551_));
 AO21x1_ASAP7_75t_R _29680_ (.A1(_07581_),
    .A2(_10537_),
    .B(_10551_),
    .Y(_03571_));
 TAPCELL_ASAP7_75t_R PHY_371 ();
 NOR2x1_ASAP7_75t_R _29682_ (.A(_00496_),
    .B(_10537_),
    .Y(_10553_));
 AO21x1_ASAP7_75t_R _29683_ (.A1(net253),
    .A2(_10537_),
    .B(_10553_),
    .Y(_03572_));
 TAPCELL_ASAP7_75t_R PHY_370 ();
 NOR2x1_ASAP7_75t_R _29685_ (.A(_00526_),
    .B(_10537_),
    .Y(_10555_));
 AO21x1_ASAP7_75t_R _29686_ (.A1(_07676_),
    .A2(_10537_),
    .B(_10555_),
    .Y(_03573_));
 TAPCELL_ASAP7_75t_R PHY_369 ();
 TAPCELL_ASAP7_75t_R PHY_368 ();
 NOR2x1_ASAP7_75t_R _29689_ (.A(_00556_),
    .B(_10537_),
    .Y(_10558_));
 AO21x1_ASAP7_75t_R _29690_ (.A1(_07738_),
    .A2(_10537_),
    .B(_10558_),
    .Y(_03574_));
 TAPCELL_ASAP7_75t_R PHY_367 ();
 NOR2x1_ASAP7_75t_R _29692_ (.A(_00586_),
    .B(_10537_),
    .Y(_10560_));
 AO21x1_ASAP7_75t_R _29693_ (.A1(_07780_),
    .A2(_10537_),
    .B(_10560_),
    .Y(_03575_));
 TAPCELL_ASAP7_75t_R PHY_366 ();
 TAPCELL_ASAP7_75t_R PHY_365 ();
 NOR2x1_ASAP7_75t_R _29696_ (.A(_00616_),
    .B(_10537_),
    .Y(_10563_));
 AO21x1_ASAP7_75t_R _29697_ (.A1(_07817_),
    .A2(_10537_),
    .B(_10563_),
    .Y(_03576_));
 TAPCELL_ASAP7_75t_R PHY_364 ();
 NOR2x1_ASAP7_75t_R _29699_ (.A(_00646_),
    .B(_10537_),
    .Y(_10565_));
 AO21x1_ASAP7_75t_R _29700_ (.A1(_07865_),
    .A2(_10537_),
    .B(_10565_),
    .Y(_03577_));
 TAPCELL_ASAP7_75t_R PHY_363 ();
 NOR2x1_ASAP7_75t_R _29702_ (.A(_00345_),
    .B(_10537_),
    .Y(_10567_));
 AO21x1_ASAP7_75t_R _29703_ (.A1(_07908_),
    .A2(_10537_),
    .B(_10567_),
    .Y(_03578_));
 TAPCELL_ASAP7_75t_R PHY_362 ();
 NOR2x1_ASAP7_75t_R _29705_ (.A(_00708_),
    .B(_10537_),
    .Y(_10569_));
 AO21x1_ASAP7_75t_R _29706_ (.A1(_07950_),
    .A2(_10537_),
    .B(_10569_),
    .Y(_03579_));
 TAPCELL_ASAP7_75t_R PHY_361 ();
 NOR2x1_ASAP7_75t_R _29708_ (.A(_00740_),
    .B(_10537_),
    .Y(_10571_));
 AO21x1_ASAP7_75t_R _29709_ (.A1(_07990_),
    .A2(_10537_),
    .B(_10571_),
    .Y(_03580_));
 TAPCELL_ASAP7_75t_R PHY_360 ();
 NOR2x1_ASAP7_75t_R _29711_ (.A(_00773_),
    .B(_10537_),
    .Y(_10573_));
 AO21x1_ASAP7_75t_R _29712_ (.A1(_08034_),
    .A2(_10537_),
    .B(_10573_),
    .Y(_03581_));
 TAPCELL_ASAP7_75t_R PHY_359 ();
 NOR2x1_ASAP7_75t_R _29714_ (.A(_00806_),
    .B(_10537_),
    .Y(_10575_));
 AO21x1_ASAP7_75t_R _29715_ (.A1(_08073_),
    .A2(_10537_),
    .B(_10575_),
    .Y(_03582_));
 TAPCELL_ASAP7_75t_R PHY_358 ();
 NOR2x1_ASAP7_75t_R _29717_ (.A(_00839_),
    .B(_10537_),
    .Y(_10577_));
 AO21x1_ASAP7_75t_R _29718_ (.A1(_08116_),
    .A2(_10537_),
    .B(_10577_),
    .Y(_03583_));
 TAPCELL_ASAP7_75t_R PHY_357 ();
 TAPCELL_ASAP7_75t_R PHY_356 ();
 NOR2x1_ASAP7_75t_R _29721_ (.A(_00871_),
    .B(_10537_),
    .Y(_10580_));
 AO21x1_ASAP7_75t_R _29722_ (.A1(net251),
    .A2(_10537_),
    .B(_10580_),
    .Y(_03584_));
 TAPCELL_ASAP7_75t_R PHY_355 ();
 NOR2x1_ASAP7_75t_R _29724_ (.A(_00904_),
    .B(_10537_),
    .Y(_10582_));
 AO21x1_ASAP7_75t_R _29725_ (.A1(_08187_),
    .A2(_10537_),
    .B(_10582_),
    .Y(_03585_));
 TAPCELL_ASAP7_75t_R PHY_354 ();
 TAPCELL_ASAP7_75t_R PHY_353 ();
 NOR2x1_ASAP7_75t_R _29728_ (.A(_00936_),
    .B(_10537_),
    .Y(_10585_));
 AO21x1_ASAP7_75t_R _29729_ (.A1(_08219_),
    .A2(_10537_),
    .B(_10585_),
    .Y(_03586_));
 TAPCELL_ASAP7_75t_R PHY_352 ();
 NOR2x1_ASAP7_75t_R _29731_ (.A(_00969_),
    .B(_10537_),
    .Y(_10587_));
 AO21x1_ASAP7_75t_R _29732_ (.A1(_08254_),
    .A2(_10537_),
    .B(_10587_),
    .Y(_03587_));
 TAPCELL_ASAP7_75t_R PHY_351 ();
 NOR2x1_ASAP7_75t_R _29734_ (.A(_01001_),
    .B(_10537_),
    .Y(_10589_));
 AO21x1_ASAP7_75t_R _29735_ (.A1(net250),
    .A2(_10537_),
    .B(_10589_),
    .Y(_03588_));
 TAPCELL_ASAP7_75t_R PHY_350 ();
 NOR2x1_ASAP7_75t_R _29737_ (.A(_01035_),
    .B(_10537_),
    .Y(_10591_));
 AO21x1_ASAP7_75t_R _29738_ (.A1(_08319_),
    .A2(_10537_),
    .B(_10591_),
    .Y(_03589_));
 TAPCELL_ASAP7_75t_R PHY_349 ();
 NOR2x1_ASAP7_75t_R _29740_ (.A(_01067_),
    .B(_10537_),
    .Y(_10593_));
 AO21x1_ASAP7_75t_R _29741_ (.A1(_08357_),
    .A2(_10537_),
    .B(_10593_),
    .Y(_03590_));
 TAPCELL_ASAP7_75t_R PHY_348 ();
 NOR2x1_ASAP7_75t_R _29743_ (.A(_01100_),
    .B(_10537_),
    .Y(_10595_));
 AO21x1_ASAP7_75t_R _29744_ (.A1(_08388_),
    .A2(_10537_),
    .B(_10595_),
    .Y(_03591_));
 TAPCELL_ASAP7_75t_R PHY_347 ();
 NOR2x1_ASAP7_75t_R _29746_ (.A(_01132_),
    .B(_10537_),
    .Y(_10597_));
 AO21x1_ASAP7_75t_R _29747_ (.A1(_08419_),
    .A2(_10537_),
    .B(_10597_),
    .Y(_03592_));
 TAPCELL_ASAP7_75t_R PHY_346 ();
 NOR2x1_ASAP7_75t_R _29749_ (.A(_01166_),
    .B(_10537_),
    .Y(_10599_));
 AO21x1_ASAP7_75t_R _29750_ (.A1(_08451_),
    .A2(_10537_),
    .B(_10599_),
    .Y(_03593_));
 TAPCELL_ASAP7_75t_R PHY_345 ();
 NOR2x1_ASAP7_75t_R _29752_ (.A(_01198_),
    .B(_10537_),
    .Y(_10601_));
 AO21x1_ASAP7_75t_R _29753_ (.A1(_08481_),
    .A2(_10537_),
    .B(_10601_),
    .Y(_03594_));
 TAPCELL_ASAP7_75t_R PHY_344 ();
 NOR2x1_ASAP7_75t_R _29755_ (.A(_01232_),
    .B(_10537_),
    .Y(_10603_));
 AO21x1_ASAP7_75t_R _29756_ (.A1(_08512_),
    .A2(_10537_),
    .B(_10603_),
    .Y(_03595_));
 TAPCELL_ASAP7_75t_R PHY_343 ();
 NOR2x1_ASAP7_75t_R _29758_ (.A(_01264_),
    .B(_10537_),
    .Y(_10605_));
 AO21x1_ASAP7_75t_R _29759_ (.A1(_08545_),
    .A2(_10537_),
    .B(_10605_),
    .Y(_03596_));
 TAPCELL_ASAP7_75t_R PHY_342 ();
 NOR2x1_ASAP7_75t_R _29761_ (.A(_01298_),
    .B(_10537_),
    .Y(_10607_));
 AO21x1_ASAP7_75t_R _29762_ (.A1(_08573_),
    .A2(_10537_),
    .B(_10607_),
    .Y(_03597_));
 AND3x4_ASAP7_75t_R _29763_ (.A(_09736_),
    .B(_09779_),
    .C(_10334_),
    .Y(_10608_));
 TAPCELL_ASAP7_75t_R PHY_341 ();
 TAPCELL_ASAP7_75t_R PHY_340 ();
 TAPCELL_ASAP7_75t_R PHY_339 ();
 NOR2x1_ASAP7_75t_R _29767_ (.A(_00314_),
    .B(_10608_),
    .Y(_10612_));
 AO21x1_ASAP7_75t_R _29768_ (.A1(_07180_),
    .A2(_10608_),
    .B(_10612_),
    .Y(_03598_));
 NOR2x1_ASAP7_75t_R _29769_ (.A(_00268_),
    .B(_10608_),
    .Y(_10613_));
 AO21x1_ASAP7_75t_R _29770_ (.A1(_07313_),
    .A2(_10608_),
    .B(_10613_),
    .Y(_03599_));
 NOR2x1_ASAP7_75t_R _29771_ (.A(_00376_),
    .B(_10608_),
    .Y(_10614_));
 AO21x1_ASAP7_75t_R _29772_ (.A1(_07398_),
    .A2(_10608_),
    .B(_10614_),
    .Y(_03600_));
 NOR2x1_ASAP7_75t_R _29773_ (.A(_00407_),
    .B(_10608_),
    .Y(_10615_));
 AO21x1_ASAP7_75t_R _29774_ (.A1(_07469_),
    .A2(_10608_),
    .B(_10615_),
    .Y(_03601_));
 NOR2x1_ASAP7_75t_R _29775_ (.A(_00437_),
    .B(_10608_),
    .Y(_10616_));
 AO21x1_ASAP7_75t_R _29776_ (.A1(_07534_),
    .A2(_10608_),
    .B(_10616_),
    .Y(_03602_));
 NOR2x1_ASAP7_75t_R _29777_ (.A(_00467_),
    .B(_10608_),
    .Y(_10617_));
 AO21x1_ASAP7_75t_R _29778_ (.A1(_07581_),
    .A2(_10608_),
    .B(_10617_),
    .Y(_03603_));
 NOR2x1_ASAP7_75t_R _29779_ (.A(_00497_),
    .B(_10608_),
    .Y(_10618_));
 AO21x1_ASAP7_75t_R _29780_ (.A1(net253),
    .A2(_10608_),
    .B(_10618_),
    .Y(_03604_));
 NOR2x1_ASAP7_75t_R _29781_ (.A(_00527_),
    .B(_10608_),
    .Y(_10619_));
 AO21x1_ASAP7_75t_R _29782_ (.A1(_07676_),
    .A2(_10608_),
    .B(_10619_),
    .Y(_03605_));
 TAPCELL_ASAP7_75t_R PHY_338 ();
 NOR2x1_ASAP7_75t_R _29784_ (.A(_00557_),
    .B(_10608_),
    .Y(_10621_));
 AO21x1_ASAP7_75t_R _29785_ (.A1(net252),
    .A2(_10608_),
    .B(_10621_),
    .Y(_03606_));
 NOR2x1_ASAP7_75t_R _29786_ (.A(_00587_),
    .B(_10608_),
    .Y(_10622_));
 AO21x1_ASAP7_75t_R _29787_ (.A1(_07780_),
    .A2(_10608_),
    .B(_10622_),
    .Y(_03607_));
 TAPCELL_ASAP7_75t_R PHY_337 ();
 NOR2x1_ASAP7_75t_R _29789_ (.A(_00617_),
    .B(_10608_),
    .Y(_10624_));
 AO21x1_ASAP7_75t_R _29790_ (.A1(_07817_),
    .A2(_10608_),
    .B(_10624_),
    .Y(_03608_));
 NOR2x1_ASAP7_75t_R _29791_ (.A(_00647_),
    .B(_10608_),
    .Y(_10625_));
 AO21x1_ASAP7_75t_R _29792_ (.A1(_07865_),
    .A2(_10608_),
    .B(_10625_),
    .Y(_03609_));
 NOR2x1_ASAP7_75t_R _29793_ (.A(_00346_),
    .B(_10608_),
    .Y(_10626_));
 AO21x1_ASAP7_75t_R _29794_ (.A1(_07908_),
    .A2(_10608_),
    .B(_10626_),
    .Y(_03610_));
 NOR2x1_ASAP7_75t_R _29795_ (.A(_00709_),
    .B(_10608_),
    .Y(_10627_));
 AO21x1_ASAP7_75t_R _29796_ (.A1(_07950_),
    .A2(_10608_),
    .B(_10627_),
    .Y(_03611_));
 NOR2x1_ASAP7_75t_R _29797_ (.A(_00741_),
    .B(_10608_),
    .Y(_10628_));
 AO21x1_ASAP7_75t_R _29798_ (.A1(_07990_),
    .A2(_10608_),
    .B(_10628_),
    .Y(_03612_));
 NOR2x1_ASAP7_75t_R _29799_ (.A(_00774_),
    .B(_10608_),
    .Y(_10629_));
 AO21x1_ASAP7_75t_R _29800_ (.A1(_08034_),
    .A2(_10608_),
    .B(_10629_),
    .Y(_03613_));
 NOR2x1_ASAP7_75t_R _29801_ (.A(_00807_),
    .B(_10608_),
    .Y(_10630_));
 AO21x1_ASAP7_75t_R _29802_ (.A1(_08073_),
    .A2(_10608_),
    .B(_10630_),
    .Y(_03614_));
 NOR2x1_ASAP7_75t_R _29803_ (.A(_00840_),
    .B(_10608_),
    .Y(_10631_));
 AO21x1_ASAP7_75t_R _29804_ (.A1(_08116_),
    .A2(_10608_),
    .B(_10631_),
    .Y(_03615_));
 TAPCELL_ASAP7_75t_R PHY_336 ();
 NOR2x1_ASAP7_75t_R _29806_ (.A(_00872_),
    .B(_10608_),
    .Y(_10633_));
 AO21x1_ASAP7_75t_R _29807_ (.A1(net251),
    .A2(_10608_),
    .B(_10633_),
    .Y(_03616_));
 NOR2x1_ASAP7_75t_R _29808_ (.A(_00905_),
    .B(_10608_),
    .Y(_10634_));
 AO21x1_ASAP7_75t_R _29809_ (.A1(_08187_),
    .A2(_10608_),
    .B(_10634_),
    .Y(_03617_));
 TAPCELL_ASAP7_75t_R PHY_335 ();
 NOR2x1_ASAP7_75t_R _29811_ (.A(_00937_),
    .B(_10608_),
    .Y(_10636_));
 AO21x1_ASAP7_75t_R _29812_ (.A1(_08219_),
    .A2(_10608_),
    .B(_10636_),
    .Y(_03618_));
 NOR2x1_ASAP7_75t_R _29813_ (.A(_00970_),
    .B(_10608_),
    .Y(_10637_));
 AO21x1_ASAP7_75t_R _29814_ (.A1(_08254_),
    .A2(_10608_),
    .B(_10637_),
    .Y(_03619_));
 NOR2x1_ASAP7_75t_R _29815_ (.A(_01002_),
    .B(_10608_),
    .Y(_10638_));
 AO21x1_ASAP7_75t_R _29816_ (.A1(net250),
    .A2(_10608_),
    .B(_10638_),
    .Y(_03620_));
 NOR2x1_ASAP7_75t_R _29817_ (.A(_01036_),
    .B(_10608_),
    .Y(_10639_));
 AO21x1_ASAP7_75t_R _29818_ (.A1(_08319_),
    .A2(_10608_),
    .B(_10639_),
    .Y(_03621_));
 NOR2x1_ASAP7_75t_R _29819_ (.A(_01068_),
    .B(_10608_),
    .Y(_10640_));
 AO21x1_ASAP7_75t_R _29820_ (.A1(_08357_),
    .A2(_10608_),
    .B(_10640_),
    .Y(_03622_));
 NOR2x1_ASAP7_75t_R _29821_ (.A(_01101_),
    .B(_10608_),
    .Y(_10641_));
 AO21x1_ASAP7_75t_R _29822_ (.A1(_08388_),
    .A2(_10608_),
    .B(_10641_),
    .Y(_03623_));
 NOR2x1_ASAP7_75t_R _29823_ (.A(_01133_),
    .B(_10608_),
    .Y(_10642_));
 AO21x1_ASAP7_75t_R _29824_ (.A1(_08419_),
    .A2(_10608_),
    .B(_10642_),
    .Y(_03624_));
 NOR2x1_ASAP7_75t_R _29825_ (.A(_01167_),
    .B(_10608_),
    .Y(_10643_));
 AO21x1_ASAP7_75t_R _29826_ (.A1(_08451_),
    .A2(_10608_),
    .B(_10643_),
    .Y(_03625_));
 NOR2x1_ASAP7_75t_R _29827_ (.A(_01199_),
    .B(_10608_),
    .Y(_10644_));
 AO21x1_ASAP7_75t_R _29828_ (.A1(_08481_),
    .A2(_10608_),
    .B(_10644_),
    .Y(_03626_));
 NOR2x1_ASAP7_75t_R _29829_ (.A(_01233_),
    .B(_10608_),
    .Y(_10645_));
 AO21x1_ASAP7_75t_R _29830_ (.A1(_08512_),
    .A2(_10608_),
    .B(_10645_),
    .Y(_03627_));
 NOR2x1_ASAP7_75t_R _29831_ (.A(_01265_),
    .B(_10608_),
    .Y(_10646_));
 AO21x1_ASAP7_75t_R _29832_ (.A1(_08545_),
    .A2(_10608_),
    .B(_10646_),
    .Y(_03628_));
 NOR2x1_ASAP7_75t_R _29833_ (.A(_01299_),
    .B(_10608_),
    .Y(_10647_));
 AO21x1_ASAP7_75t_R _29834_ (.A1(_08573_),
    .A2(_10608_),
    .B(_10647_),
    .Y(_03629_));
 AND4x2_ASAP7_75t_R _29835_ (.A(_00323_),
    .B(_00184_),
    .C(_09940_),
    .D(_10334_),
    .Y(_10648_));
 TAPCELL_ASAP7_75t_R PHY_334 ();
 TAPCELL_ASAP7_75t_R PHY_333 ();
 TAPCELL_ASAP7_75t_R PHY_332 ();
 NOR2x1_ASAP7_75t_R _29839_ (.A(_00315_),
    .B(_10648_),
    .Y(_10652_));
 AO21x1_ASAP7_75t_R _29840_ (.A1(_07180_),
    .A2(_10648_),
    .B(_10652_),
    .Y(_03630_));
 NOR2x1_ASAP7_75t_R _29841_ (.A(_00269_),
    .B(net260),
    .Y(_10653_));
 AO21x1_ASAP7_75t_R _29842_ (.A1(_07313_),
    .A2(net260),
    .B(_10653_),
    .Y(_03631_));
 NOR2x1_ASAP7_75t_R _29843_ (.A(_00377_),
    .B(net260),
    .Y(_10654_));
 AO21x1_ASAP7_75t_R _29844_ (.A1(_07398_),
    .A2(net260),
    .B(_10654_),
    .Y(_03632_));
 NOR2x1_ASAP7_75t_R _29845_ (.A(_00408_),
    .B(net260),
    .Y(_10655_));
 AO21x1_ASAP7_75t_R _29846_ (.A1(_07469_),
    .A2(net260),
    .B(_10655_),
    .Y(_03633_));
 NOR2x1_ASAP7_75t_R _29847_ (.A(_00438_),
    .B(_10648_),
    .Y(_10656_));
 AO21x1_ASAP7_75t_R _29848_ (.A1(_07534_),
    .A2(_10648_),
    .B(_10656_),
    .Y(_03634_));
 NOR2x1_ASAP7_75t_R _29849_ (.A(_00468_),
    .B(net260),
    .Y(_10657_));
 AO21x1_ASAP7_75t_R _29850_ (.A1(_07581_),
    .A2(net260),
    .B(_10657_),
    .Y(_03635_));
 NOR2x1_ASAP7_75t_R _29851_ (.A(_00498_),
    .B(_10648_),
    .Y(_10658_));
 AO21x1_ASAP7_75t_R _29852_ (.A1(net253),
    .A2(_10648_),
    .B(_10658_),
    .Y(_03636_));
 NOR2x1_ASAP7_75t_R _29853_ (.A(_00528_),
    .B(net260),
    .Y(_10659_));
 AO21x1_ASAP7_75t_R _29854_ (.A1(_07676_),
    .A2(net260),
    .B(_10659_),
    .Y(_03637_));
 TAPCELL_ASAP7_75t_R PHY_331 ();
 NOR2x1_ASAP7_75t_R _29856_ (.A(_00558_),
    .B(net260),
    .Y(_10661_));
 AO21x1_ASAP7_75t_R _29857_ (.A1(net252),
    .A2(net260),
    .B(_10661_),
    .Y(_03638_));
 NOR2x1_ASAP7_75t_R _29858_ (.A(_00588_),
    .B(_10648_),
    .Y(_10662_));
 AO21x1_ASAP7_75t_R _29859_ (.A1(_07780_),
    .A2(_10648_),
    .B(_10662_),
    .Y(_03639_));
 TAPCELL_ASAP7_75t_R PHY_330 ();
 NOR2x1_ASAP7_75t_R _29861_ (.A(_00618_),
    .B(net260),
    .Y(_10664_));
 AO21x1_ASAP7_75t_R _29862_ (.A1(_07817_),
    .A2(net260),
    .B(_10664_),
    .Y(_03640_));
 NOR2x1_ASAP7_75t_R _29863_ (.A(_00648_),
    .B(net260),
    .Y(_10665_));
 AO21x1_ASAP7_75t_R _29864_ (.A1(_07865_),
    .A2(net260),
    .B(_10665_),
    .Y(_03641_));
 NOR2x1_ASAP7_75t_R _29865_ (.A(_00347_),
    .B(_10648_),
    .Y(_10666_));
 AO21x1_ASAP7_75t_R _29866_ (.A1(_07908_),
    .A2(_10648_),
    .B(_10666_),
    .Y(_03642_));
 NOR2x1_ASAP7_75t_R _29867_ (.A(_00710_),
    .B(net261),
    .Y(_10667_));
 AO21x1_ASAP7_75t_R _29868_ (.A1(_07950_),
    .A2(net261),
    .B(_10667_),
    .Y(_03643_));
 NOR2x1_ASAP7_75t_R _29869_ (.A(_00742_),
    .B(_10648_),
    .Y(_10668_));
 AO21x1_ASAP7_75t_R _29870_ (.A1(_07990_),
    .A2(_10648_),
    .B(_10668_),
    .Y(_03644_));
 NOR2x1_ASAP7_75t_R _29871_ (.A(_00775_),
    .B(net261),
    .Y(_10669_));
 AO21x1_ASAP7_75t_R _29872_ (.A1(_08034_),
    .A2(net261),
    .B(_10669_),
    .Y(_03645_));
 NOR2x1_ASAP7_75t_R _29873_ (.A(_00808_),
    .B(net260),
    .Y(_10670_));
 AO21x1_ASAP7_75t_R _29874_ (.A1(_08073_),
    .A2(net260),
    .B(_10670_),
    .Y(_03646_));
 NOR2x1_ASAP7_75t_R _29875_ (.A(_00841_),
    .B(net260),
    .Y(_10671_));
 AO21x1_ASAP7_75t_R _29876_ (.A1(_08116_),
    .A2(net260),
    .B(_10671_),
    .Y(_03647_));
 TAPCELL_ASAP7_75t_R PHY_329 ();
 NOR2x1_ASAP7_75t_R _29878_ (.A(_00873_),
    .B(net261),
    .Y(_10673_));
 AO21x1_ASAP7_75t_R _29879_ (.A1(net251),
    .A2(net261),
    .B(_10673_),
    .Y(_03648_));
 NOR2x1_ASAP7_75t_R _29880_ (.A(_00906_),
    .B(net261),
    .Y(_10674_));
 AO21x1_ASAP7_75t_R _29881_ (.A1(_08187_),
    .A2(net261),
    .B(_10674_),
    .Y(_03649_));
 TAPCELL_ASAP7_75t_R PHY_328 ();
 NOR2x1_ASAP7_75t_R _29883_ (.A(_00938_),
    .B(net260),
    .Y(_10676_));
 AO21x1_ASAP7_75t_R _29884_ (.A1(_08219_),
    .A2(net260),
    .B(_10676_),
    .Y(_03650_));
 NOR2x1_ASAP7_75t_R _29885_ (.A(_00971_),
    .B(net261),
    .Y(_10677_));
 AO21x1_ASAP7_75t_R _29886_ (.A1(_08254_),
    .A2(net261),
    .B(_10677_),
    .Y(_03651_));
 NOR2x1_ASAP7_75t_R _29887_ (.A(_01003_),
    .B(_10648_),
    .Y(_10678_));
 AO21x1_ASAP7_75t_R _29888_ (.A1(net250),
    .A2(_10648_),
    .B(_10678_),
    .Y(_03652_));
 NOR2x1_ASAP7_75t_R _29889_ (.A(_01037_),
    .B(net261),
    .Y(_10679_));
 AO21x1_ASAP7_75t_R _29890_ (.A1(_08319_),
    .A2(net261),
    .B(_10679_),
    .Y(_03653_));
 NOR2x1_ASAP7_75t_R _29891_ (.A(_01069_),
    .B(net261),
    .Y(_10680_));
 AO21x1_ASAP7_75t_R _29892_ (.A1(_08357_),
    .A2(net261),
    .B(_10680_),
    .Y(_03654_));
 NOR2x1_ASAP7_75t_R _29893_ (.A(_01102_),
    .B(net261),
    .Y(_10681_));
 AO21x1_ASAP7_75t_R _29894_ (.A1(_08388_),
    .A2(net261),
    .B(_10681_),
    .Y(_03655_));
 NOR2x1_ASAP7_75t_R _29895_ (.A(_01134_),
    .B(net261),
    .Y(_10682_));
 AO21x1_ASAP7_75t_R _29896_ (.A1(_08419_),
    .A2(net261),
    .B(_10682_),
    .Y(_03656_));
 NOR2x1_ASAP7_75t_R _29897_ (.A(_01168_),
    .B(net261),
    .Y(_10683_));
 AO21x1_ASAP7_75t_R _29898_ (.A1(_08451_),
    .A2(net261),
    .B(_10683_),
    .Y(_03657_));
 NOR2x1_ASAP7_75t_R _29899_ (.A(_01200_),
    .B(_10648_),
    .Y(_10684_));
 AO21x1_ASAP7_75t_R _29900_ (.A1(_08481_),
    .A2(_10648_),
    .B(_10684_),
    .Y(_03658_));
 NOR2x1_ASAP7_75t_R _29901_ (.A(_01234_),
    .B(net261),
    .Y(_10685_));
 AO21x1_ASAP7_75t_R _29902_ (.A1(_08512_),
    .A2(net261),
    .B(_10685_),
    .Y(_03659_));
 NOR2x1_ASAP7_75t_R _29903_ (.A(_01266_),
    .B(net260),
    .Y(_10686_));
 AO21x1_ASAP7_75t_R _29904_ (.A1(_08545_),
    .A2(net260),
    .B(_10686_),
    .Y(_03660_));
 NOR2x1_ASAP7_75t_R _29905_ (.A(_01300_),
    .B(net260),
    .Y(_10687_));
 AO21x1_ASAP7_75t_R _29906_ (.A1(_08573_),
    .A2(net260),
    .B(_10687_),
    .Y(_03661_));
 AND3x4_ASAP7_75t_R _29907_ (.A(_06882_),
    .B(_09940_),
    .C(_10334_),
    .Y(_10688_));
 TAPCELL_ASAP7_75t_R PHY_327 ();
 TAPCELL_ASAP7_75t_R PHY_326 ();
 TAPCELL_ASAP7_75t_R PHY_325 ();
 NOR2x1_ASAP7_75t_R _29911_ (.A(_00316_),
    .B(_10688_),
    .Y(_10692_));
 AO21x1_ASAP7_75t_R _29912_ (.A1(_07180_),
    .A2(_10688_),
    .B(_10692_),
    .Y(_03662_));
 NOR2x1_ASAP7_75t_R _29913_ (.A(_00270_),
    .B(_10688_),
    .Y(_10693_));
 AO21x1_ASAP7_75t_R _29914_ (.A1(_07313_),
    .A2(_10688_),
    .B(_10693_),
    .Y(_03663_));
 NOR2x1_ASAP7_75t_R _29915_ (.A(_00378_),
    .B(_10688_),
    .Y(_10694_));
 AO21x1_ASAP7_75t_R _29916_ (.A1(_07398_),
    .A2(_10688_),
    .B(_10694_),
    .Y(_03664_));
 NOR2x1_ASAP7_75t_R _29917_ (.A(_00409_),
    .B(_10688_),
    .Y(_10695_));
 AO21x1_ASAP7_75t_R _29918_ (.A1(_07469_),
    .A2(_10688_),
    .B(_10695_),
    .Y(_03665_));
 NOR2x1_ASAP7_75t_R _29919_ (.A(_00439_),
    .B(_10688_),
    .Y(_10696_));
 AO21x1_ASAP7_75t_R _29920_ (.A1(_07534_),
    .A2(_10688_),
    .B(_10696_),
    .Y(_03666_));
 NOR2x1_ASAP7_75t_R _29921_ (.A(_00469_),
    .B(_10688_),
    .Y(_10697_));
 AO21x1_ASAP7_75t_R _29922_ (.A1(_07581_),
    .A2(_10688_),
    .B(_10697_),
    .Y(_03667_));
 NOR2x1_ASAP7_75t_R _29923_ (.A(_00499_),
    .B(_10688_),
    .Y(_10698_));
 AO21x1_ASAP7_75t_R _29924_ (.A1(net253),
    .A2(_10688_),
    .B(_10698_),
    .Y(_03668_));
 NOR2x1_ASAP7_75t_R _29925_ (.A(_00529_),
    .B(_10688_),
    .Y(_10699_));
 AO21x1_ASAP7_75t_R _29926_ (.A1(_07676_),
    .A2(_10688_),
    .B(_10699_),
    .Y(_03669_));
 TAPCELL_ASAP7_75t_R PHY_324 ();
 NOR2x1_ASAP7_75t_R _29928_ (.A(_00559_),
    .B(_10688_),
    .Y(_10701_));
 AO21x1_ASAP7_75t_R _29929_ (.A1(net252),
    .A2(_10688_),
    .B(_10701_),
    .Y(_03670_));
 NOR2x1_ASAP7_75t_R _29930_ (.A(_00589_),
    .B(_10688_),
    .Y(_10702_));
 AO21x1_ASAP7_75t_R _29931_ (.A1(_07780_),
    .A2(_10688_),
    .B(_10702_),
    .Y(_03671_));
 TAPCELL_ASAP7_75t_R PHY_323 ();
 NOR2x1_ASAP7_75t_R _29933_ (.A(_00619_),
    .B(_10688_),
    .Y(_10704_));
 AO21x1_ASAP7_75t_R _29934_ (.A1(_07817_),
    .A2(_10688_),
    .B(_10704_),
    .Y(_03672_));
 NOR2x1_ASAP7_75t_R _29935_ (.A(_00649_),
    .B(_10688_),
    .Y(_10705_));
 AO21x1_ASAP7_75t_R _29936_ (.A1(_07865_),
    .A2(_10688_),
    .B(_10705_),
    .Y(_03673_));
 NOR2x1_ASAP7_75t_R _29937_ (.A(_00348_),
    .B(_10688_),
    .Y(_10706_));
 AO21x1_ASAP7_75t_R _29938_ (.A1(_07908_),
    .A2(_10688_),
    .B(_10706_),
    .Y(_03674_));
 NOR2x1_ASAP7_75t_R _29939_ (.A(_00711_),
    .B(_10688_),
    .Y(_10707_));
 AO21x1_ASAP7_75t_R _29940_ (.A1(_07950_),
    .A2(_10688_),
    .B(_10707_),
    .Y(_03675_));
 NOR2x1_ASAP7_75t_R _29941_ (.A(_00743_),
    .B(_10688_),
    .Y(_10708_));
 AO21x1_ASAP7_75t_R _29942_ (.A1(_07990_),
    .A2(_10688_),
    .B(_10708_),
    .Y(_03676_));
 NOR2x1_ASAP7_75t_R _29943_ (.A(_00776_),
    .B(_10688_),
    .Y(_10709_));
 AO21x1_ASAP7_75t_R _29944_ (.A1(_08034_),
    .A2(_10688_),
    .B(_10709_),
    .Y(_03677_));
 NOR2x1_ASAP7_75t_R _29945_ (.A(_00809_),
    .B(_10688_),
    .Y(_10710_));
 AO21x1_ASAP7_75t_R _29946_ (.A1(_08073_),
    .A2(_10688_),
    .B(_10710_),
    .Y(_03678_));
 NOR2x1_ASAP7_75t_R _29947_ (.A(_00842_),
    .B(_10688_),
    .Y(_10711_));
 AO21x1_ASAP7_75t_R _29948_ (.A1(_08116_),
    .A2(_10688_),
    .B(_10711_),
    .Y(_03679_));
 TAPCELL_ASAP7_75t_R PHY_322 ();
 NOR2x1_ASAP7_75t_R _29950_ (.A(_00874_),
    .B(_10688_),
    .Y(_10713_));
 AO21x1_ASAP7_75t_R _29951_ (.A1(net251),
    .A2(_10688_),
    .B(_10713_),
    .Y(_03680_));
 NOR2x1_ASAP7_75t_R _29952_ (.A(_00907_),
    .B(_10688_),
    .Y(_10714_));
 AO21x1_ASAP7_75t_R _29953_ (.A1(_08187_),
    .A2(_10688_),
    .B(_10714_),
    .Y(_03681_));
 TAPCELL_ASAP7_75t_R PHY_321 ();
 NOR2x1_ASAP7_75t_R _29955_ (.A(_00939_),
    .B(_10688_),
    .Y(_10716_));
 AO21x1_ASAP7_75t_R _29956_ (.A1(_08219_),
    .A2(_10688_),
    .B(_10716_),
    .Y(_03682_));
 NOR2x1_ASAP7_75t_R _29957_ (.A(_00972_),
    .B(_10688_),
    .Y(_10717_));
 AO21x1_ASAP7_75t_R _29958_ (.A1(_08254_),
    .A2(_10688_),
    .B(_10717_),
    .Y(_03683_));
 NOR2x1_ASAP7_75t_R _29959_ (.A(_01004_),
    .B(_10688_),
    .Y(_10718_));
 AO21x1_ASAP7_75t_R _29960_ (.A1(net250),
    .A2(_10688_),
    .B(_10718_),
    .Y(_03684_));
 NOR2x1_ASAP7_75t_R _29961_ (.A(_01038_),
    .B(_10688_),
    .Y(_10719_));
 AO21x1_ASAP7_75t_R _29962_ (.A1(_08319_),
    .A2(_10688_),
    .B(_10719_),
    .Y(_03685_));
 NOR2x1_ASAP7_75t_R _29963_ (.A(_01070_),
    .B(_10688_),
    .Y(_10720_));
 AO21x1_ASAP7_75t_R _29964_ (.A1(_08357_),
    .A2(_10688_),
    .B(_10720_),
    .Y(_03686_));
 NOR2x1_ASAP7_75t_R _29965_ (.A(_01103_),
    .B(_10688_),
    .Y(_10721_));
 AO21x1_ASAP7_75t_R _29966_ (.A1(_08388_),
    .A2(_10688_),
    .B(_10721_),
    .Y(_03687_));
 NOR2x1_ASAP7_75t_R _29967_ (.A(_01135_),
    .B(_10688_),
    .Y(_10722_));
 AO21x1_ASAP7_75t_R _29968_ (.A1(_08419_),
    .A2(_10688_),
    .B(_10722_),
    .Y(_03688_));
 NOR2x1_ASAP7_75t_R _29969_ (.A(_01169_),
    .B(_10688_),
    .Y(_10723_));
 AO21x1_ASAP7_75t_R _29970_ (.A1(_08451_),
    .A2(_10688_),
    .B(_10723_),
    .Y(_03689_));
 NOR2x1_ASAP7_75t_R _29971_ (.A(_01201_),
    .B(_10688_),
    .Y(_10724_));
 AO21x1_ASAP7_75t_R _29972_ (.A1(_08481_),
    .A2(_10688_),
    .B(_10724_),
    .Y(_03690_));
 NOR2x1_ASAP7_75t_R _29973_ (.A(_01235_),
    .B(_10688_),
    .Y(_10725_));
 AO21x1_ASAP7_75t_R _29974_ (.A1(_08512_),
    .A2(_10688_),
    .B(_10725_),
    .Y(_03691_));
 NOR2x1_ASAP7_75t_R _29975_ (.A(_01267_),
    .B(_10688_),
    .Y(_10726_));
 AO21x1_ASAP7_75t_R _29976_ (.A1(_08545_),
    .A2(_10688_),
    .B(_10726_),
    .Y(_03692_));
 NOR2x1_ASAP7_75t_R _29977_ (.A(_01301_),
    .B(_10688_),
    .Y(_10727_));
 AO21x1_ASAP7_75t_R _29978_ (.A1(_08573_),
    .A2(_10688_),
    .B(_10727_),
    .Y(_03693_));
 AND3x4_ASAP7_75t_R _29979_ (.A(_09663_),
    .B(_09940_),
    .C(_10334_),
    .Y(_10728_));
 TAPCELL_ASAP7_75t_R PHY_320 ();
 TAPCELL_ASAP7_75t_R PHY_319 ();
 TAPCELL_ASAP7_75t_R PHY_318 ();
 NOR2x1_ASAP7_75t_R _29983_ (.A(_00317_),
    .B(_10728_),
    .Y(_10732_));
 AO21x1_ASAP7_75t_R _29984_ (.A1(_07180_),
    .A2(_10728_),
    .B(_10732_),
    .Y(_03694_));
 NOR2x1_ASAP7_75t_R _29985_ (.A(_00271_),
    .B(_10728_),
    .Y(_10733_));
 AO21x1_ASAP7_75t_R _29986_ (.A1(_07313_),
    .A2(_10728_),
    .B(_10733_),
    .Y(_03695_));
 NOR2x1_ASAP7_75t_R _29987_ (.A(_00379_),
    .B(_10728_),
    .Y(_10734_));
 AO21x1_ASAP7_75t_R _29988_ (.A1(_07398_),
    .A2(_10728_),
    .B(_10734_),
    .Y(_03696_));
 NOR2x1_ASAP7_75t_R _29989_ (.A(_00410_),
    .B(_10728_),
    .Y(_10735_));
 AO21x1_ASAP7_75t_R _29990_ (.A1(_07469_),
    .A2(_10728_),
    .B(_10735_),
    .Y(_03697_));
 NOR2x1_ASAP7_75t_R _29991_ (.A(_00440_),
    .B(_10728_),
    .Y(_10736_));
 AO21x1_ASAP7_75t_R _29992_ (.A1(_07534_),
    .A2(_10728_),
    .B(_10736_),
    .Y(_03698_));
 NOR2x1_ASAP7_75t_R _29993_ (.A(_00470_),
    .B(_10728_),
    .Y(_10737_));
 AO21x1_ASAP7_75t_R _29994_ (.A1(_07581_),
    .A2(_10728_),
    .B(_10737_),
    .Y(_03699_));
 NOR2x1_ASAP7_75t_R _29995_ (.A(_00500_),
    .B(_10728_),
    .Y(_10738_));
 AO21x1_ASAP7_75t_R _29996_ (.A1(net253),
    .A2(_10728_),
    .B(_10738_),
    .Y(_03700_));
 NOR2x1_ASAP7_75t_R _29997_ (.A(_00530_),
    .B(_10728_),
    .Y(_10739_));
 AO21x1_ASAP7_75t_R _29998_ (.A1(_07676_),
    .A2(_10728_),
    .B(_10739_),
    .Y(_03701_));
 TAPCELL_ASAP7_75t_R PHY_317 ();
 NOR2x1_ASAP7_75t_R _30000_ (.A(_00560_),
    .B(_10728_),
    .Y(_10741_));
 AO21x1_ASAP7_75t_R _30001_ (.A1(net252),
    .A2(_10728_),
    .B(_10741_),
    .Y(_03702_));
 NOR2x1_ASAP7_75t_R _30002_ (.A(_00590_),
    .B(_10728_),
    .Y(_10742_));
 AO21x1_ASAP7_75t_R _30003_ (.A1(_07780_),
    .A2(_10728_),
    .B(_10742_),
    .Y(_03703_));
 TAPCELL_ASAP7_75t_R PHY_316 ();
 NOR2x1_ASAP7_75t_R _30005_ (.A(_00620_),
    .B(_10728_),
    .Y(_10744_));
 AO21x1_ASAP7_75t_R _30006_ (.A1(_07817_),
    .A2(_10728_),
    .B(_10744_),
    .Y(_03704_));
 NOR2x1_ASAP7_75t_R _30007_ (.A(_00650_),
    .B(_10728_),
    .Y(_10745_));
 AO21x1_ASAP7_75t_R _30008_ (.A1(_07865_),
    .A2(_10728_),
    .B(_10745_),
    .Y(_03705_));
 NOR2x1_ASAP7_75t_R _30009_ (.A(_00349_),
    .B(_10728_),
    .Y(_10746_));
 AO21x1_ASAP7_75t_R _30010_ (.A1(_07908_),
    .A2(_10728_),
    .B(_10746_),
    .Y(_03706_));
 NOR2x1_ASAP7_75t_R _30011_ (.A(_00712_),
    .B(_10728_),
    .Y(_10747_));
 AO21x1_ASAP7_75t_R _30012_ (.A1(_07950_),
    .A2(_10728_),
    .B(_10747_),
    .Y(_03707_));
 NOR2x1_ASAP7_75t_R _30013_ (.A(_00744_),
    .B(_10728_),
    .Y(_10748_));
 AO21x1_ASAP7_75t_R _30014_ (.A1(_07990_),
    .A2(_10728_),
    .B(_10748_),
    .Y(_03708_));
 NOR2x1_ASAP7_75t_R _30015_ (.A(_00777_),
    .B(_10728_),
    .Y(_10749_));
 AO21x1_ASAP7_75t_R _30016_ (.A1(_08034_),
    .A2(_10728_),
    .B(_10749_),
    .Y(_03709_));
 NOR2x1_ASAP7_75t_R _30017_ (.A(_00810_),
    .B(_10728_),
    .Y(_10750_));
 AO21x1_ASAP7_75t_R _30018_ (.A1(_08073_),
    .A2(_10728_),
    .B(_10750_),
    .Y(_03710_));
 NOR2x1_ASAP7_75t_R _30019_ (.A(_00843_),
    .B(_10728_),
    .Y(_10751_));
 AO21x1_ASAP7_75t_R _30020_ (.A1(_08116_),
    .A2(_10728_),
    .B(_10751_),
    .Y(_03711_));
 TAPCELL_ASAP7_75t_R PHY_315 ();
 NOR2x1_ASAP7_75t_R _30022_ (.A(_00875_),
    .B(_10728_),
    .Y(_10753_));
 AO21x1_ASAP7_75t_R _30023_ (.A1(net251),
    .A2(_10728_),
    .B(_10753_),
    .Y(_03712_));
 NOR2x1_ASAP7_75t_R _30024_ (.A(_00908_),
    .B(_10728_),
    .Y(_10754_));
 AO21x1_ASAP7_75t_R _30025_ (.A1(_08187_),
    .A2(_10728_),
    .B(_10754_),
    .Y(_03713_));
 TAPCELL_ASAP7_75t_R PHY_314 ();
 NOR2x1_ASAP7_75t_R _30027_ (.A(_00940_),
    .B(_10728_),
    .Y(_10756_));
 AO21x1_ASAP7_75t_R _30028_ (.A1(_08219_),
    .A2(_10728_),
    .B(_10756_),
    .Y(_03714_));
 NOR2x1_ASAP7_75t_R _30029_ (.A(_00973_),
    .B(_10728_),
    .Y(_10757_));
 AO21x1_ASAP7_75t_R _30030_ (.A1(_08254_),
    .A2(_10728_),
    .B(_10757_),
    .Y(_03715_));
 NOR2x1_ASAP7_75t_R _30031_ (.A(_01005_),
    .B(_10728_),
    .Y(_10758_));
 AO21x1_ASAP7_75t_R _30032_ (.A1(net250),
    .A2(_10728_),
    .B(_10758_),
    .Y(_03716_));
 NOR2x1_ASAP7_75t_R _30033_ (.A(_01039_),
    .B(_10728_),
    .Y(_10759_));
 AO21x1_ASAP7_75t_R _30034_ (.A1(_08319_),
    .A2(_10728_),
    .B(_10759_),
    .Y(_03717_));
 NOR2x1_ASAP7_75t_R _30035_ (.A(_01071_),
    .B(_10728_),
    .Y(_10760_));
 AO21x1_ASAP7_75t_R _30036_ (.A1(_08357_),
    .A2(_10728_),
    .B(_10760_),
    .Y(_03718_));
 NOR2x1_ASAP7_75t_R _30037_ (.A(_01104_),
    .B(_10728_),
    .Y(_10761_));
 AO21x1_ASAP7_75t_R _30038_ (.A1(_08388_),
    .A2(_10728_),
    .B(_10761_),
    .Y(_03719_));
 NOR2x1_ASAP7_75t_R _30039_ (.A(_01136_),
    .B(_10728_),
    .Y(_10762_));
 AO21x1_ASAP7_75t_R _30040_ (.A1(_08419_),
    .A2(_10728_),
    .B(_10762_),
    .Y(_03720_));
 NOR2x1_ASAP7_75t_R _30041_ (.A(_01170_),
    .B(_10728_),
    .Y(_10763_));
 AO21x1_ASAP7_75t_R _30042_ (.A1(_08451_),
    .A2(_10728_),
    .B(_10763_),
    .Y(_03721_));
 NOR2x1_ASAP7_75t_R _30043_ (.A(_01202_),
    .B(_10728_),
    .Y(_10764_));
 AO21x1_ASAP7_75t_R _30044_ (.A1(_08481_),
    .A2(_10728_),
    .B(_10764_),
    .Y(_03722_));
 NOR2x1_ASAP7_75t_R _30045_ (.A(_01236_),
    .B(_10728_),
    .Y(_10765_));
 AO21x1_ASAP7_75t_R _30046_ (.A1(_08512_),
    .A2(_10728_),
    .B(_10765_),
    .Y(_03723_));
 NOR2x1_ASAP7_75t_R _30047_ (.A(_01268_),
    .B(_10728_),
    .Y(_10766_));
 AO21x1_ASAP7_75t_R _30048_ (.A1(_08545_),
    .A2(_10728_),
    .B(_10766_),
    .Y(_03724_));
 NOR2x1_ASAP7_75t_R _30049_ (.A(_01302_),
    .B(_10728_),
    .Y(_10767_));
 AO21x1_ASAP7_75t_R _30050_ (.A1(_08573_),
    .A2(_10728_),
    .B(_10767_),
    .Y(_03725_));
 AND3x4_ASAP7_75t_R _30051_ (.A(_09736_),
    .B(_09940_),
    .C(_10334_),
    .Y(_10768_));
 TAPCELL_ASAP7_75t_R PHY_313 ();
 TAPCELL_ASAP7_75t_R PHY_312 ();
 TAPCELL_ASAP7_75t_R PHY_311 ();
 NOR2x1_ASAP7_75t_R _30055_ (.A(_00318_),
    .B(_10768_),
    .Y(_10772_));
 AO21x1_ASAP7_75t_R _30056_ (.A1(_07180_),
    .A2(_10768_),
    .B(_10772_),
    .Y(_03726_));
 NOR2x1_ASAP7_75t_R _30057_ (.A(_00272_),
    .B(_10768_),
    .Y(_10773_));
 AO21x1_ASAP7_75t_R _30058_ (.A1(_07313_),
    .A2(_10768_),
    .B(_10773_),
    .Y(_03727_));
 NOR2x1_ASAP7_75t_R _30059_ (.A(_00380_),
    .B(_10768_),
    .Y(_10774_));
 AO21x1_ASAP7_75t_R _30060_ (.A1(_07398_),
    .A2(_10768_),
    .B(_10774_),
    .Y(_03728_));
 NOR2x1_ASAP7_75t_R _30061_ (.A(_00411_),
    .B(_10768_),
    .Y(_10775_));
 AO21x1_ASAP7_75t_R _30062_ (.A1(_07469_),
    .A2(_10768_),
    .B(_10775_),
    .Y(_03729_));
 NOR2x1_ASAP7_75t_R _30063_ (.A(_00441_),
    .B(_10768_),
    .Y(_10776_));
 AO21x1_ASAP7_75t_R _30064_ (.A1(_07534_),
    .A2(_10768_),
    .B(_10776_),
    .Y(_03730_));
 NOR2x1_ASAP7_75t_R _30065_ (.A(_00471_),
    .B(_10768_),
    .Y(_10777_));
 AO21x1_ASAP7_75t_R _30066_ (.A1(_07581_),
    .A2(_10768_),
    .B(_10777_),
    .Y(_03731_));
 NOR2x1_ASAP7_75t_R _30067_ (.A(_00501_),
    .B(_10768_),
    .Y(_10778_));
 AO21x1_ASAP7_75t_R _30068_ (.A1(net253),
    .A2(_10768_),
    .B(_10778_),
    .Y(_03732_));
 NOR2x1_ASAP7_75t_R _30069_ (.A(_00531_),
    .B(_10768_),
    .Y(_10779_));
 AO21x1_ASAP7_75t_R _30070_ (.A1(_07676_),
    .A2(_10768_),
    .B(_10779_),
    .Y(_03733_));
 TAPCELL_ASAP7_75t_R PHY_310 ();
 NOR2x1_ASAP7_75t_R _30072_ (.A(_00561_),
    .B(_10768_),
    .Y(_10781_));
 AO21x1_ASAP7_75t_R _30073_ (.A1(net252),
    .A2(_10768_),
    .B(_10781_),
    .Y(_03734_));
 NOR2x1_ASAP7_75t_R _30074_ (.A(_00591_),
    .B(_10768_),
    .Y(_10782_));
 AO21x1_ASAP7_75t_R _30075_ (.A1(_07780_),
    .A2(_10768_),
    .B(_10782_),
    .Y(_03735_));
 TAPCELL_ASAP7_75t_R PHY_309 ();
 NOR2x1_ASAP7_75t_R _30077_ (.A(_00621_),
    .B(_10768_),
    .Y(_10784_));
 AO21x1_ASAP7_75t_R _30078_ (.A1(_07817_),
    .A2(_10768_),
    .B(_10784_),
    .Y(_03736_));
 NOR2x1_ASAP7_75t_R _30079_ (.A(_00651_),
    .B(_10768_),
    .Y(_10785_));
 AO21x1_ASAP7_75t_R _30080_ (.A1(_07865_),
    .A2(_10768_),
    .B(_10785_),
    .Y(_03737_));
 NOR2x1_ASAP7_75t_R _30081_ (.A(_00350_),
    .B(_10768_),
    .Y(_10786_));
 AO21x1_ASAP7_75t_R _30082_ (.A1(_07908_),
    .A2(_10768_),
    .B(_10786_),
    .Y(_03738_));
 NOR2x1_ASAP7_75t_R _30083_ (.A(_00713_),
    .B(_10768_),
    .Y(_10787_));
 AO21x1_ASAP7_75t_R _30084_ (.A1(_07950_),
    .A2(_10768_),
    .B(_10787_),
    .Y(_03739_));
 NOR2x1_ASAP7_75t_R _30085_ (.A(_00745_),
    .B(_10768_),
    .Y(_10788_));
 AO21x1_ASAP7_75t_R _30086_ (.A1(_07990_),
    .A2(_10768_),
    .B(_10788_),
    .Y(_03740_));
 NOR2x1_ASAP7_75t_R _30087_ (.A(_00778_),
    .B(_10768_),
    .Y(_10789_));
 AO21x1_ASAP7_75t_R _30088_ (.A1(_08034_),
    .A2(_10768_),
    .B(_10789_),
    .Y(_03741_));
 NOR2x1_ASAP7_75t_R _30089_ (.A(_00811_),
    .B(_10768_),
    .Y(_10790_));
 AO21x1_ASAP7_75t_R _30090_ (.A1(_08073_),
    .A2(_10768_),
    .B(_10790_),
    .Y(_03742_));
 NOR2x1_ASAP7_75t_R _30091_ (.A(_00844_),
    .B(_10768_),
    .Y(_10791_));
 AO21x1_ASAP7_75t_R _30092_ (.A1(_08116_),
    .A2(_10768_),
    .B(_10791_),
    .Y(_03743_));
 TAPCELL_ASAP7_75t_R PHY_308 ();
 NOR2x1_ASAP7_75t_R _30094_ (.A(_00876_),
    .B(_10768_),
    .Y(_10793_));
 AO21x1_ASAP7_75t_R _30095_ (.A1(net251),
    .A2(_10768_),
    .B(_10793_),
    .Y(_03744_));
 NOR2x1_ASAP7_75t_R _30096_ (.A(_00909_),
    .B(_10768_),
    .Y(_10794_));
 AO21x1_ASAP7_75t_R _30097_ (.A1(_08187_),
    .A2(_10768_),
    .B(_10794_),
    .Y(_03745_));
 TAPCELL_ASAP7_75t_R PHY_307 ();
 NOR2x1_ASAP7_75t_R _30099_ (.A(_00941_),
    .B(_10768_),
    .Y(_10796_));
 AO21x1_ASAP7_75t_R _30100_ (.A1(_08219_),
    .A2(_10768_),
    .B(_10796_),
    .Y(_03746_));
 NOR2x1_ASAP7_75t_R _30101_ (.A(_00974_),
    .B(_10768_),
    .Y(_10797_));
 AO21x1_ASAP7_75t_R _30102_ (.A1(_08254_),
    .A2(_10768_),
    .B(_10797_),
    .Y(_03747_));
 NOR2x1_ASAP7_75t_R _30103_ (.A(_01006_),
    .B(_10768_),
    .Y(_10798_));
 AO21x1_ASAP7_75t_R _30104_ (.A1(net250),
    .A2(_10768_),
    .B(_10798_),
    .Y(_03748_));
 NOR2x1_ASAP7_75t_R _30105_ (.A(_01040_),
    .B(_10768_),
    .Y(_10799_));
 AO21x1_ASAP7_75t_R _30106_ (.A1(_08319_),
    .A2(_10768_),
    .B(_10799_),
    .Y(_03749_));
 NOR2x1_ASAP7_75t_R _30107_ (.A(_01072_),
    .B(_10768_),
    .Y(_10800_));
 AO21x1_ASAP7_75t_R _30108_ (.A1(_08357_),
    .A2(_10768_),
    .B(_10800_),
    .Y(_03750_));
 NOR2x1_ASAP7_75t_R _30109_ (.A(_01105_),
    .B(_10768_),
    .Y(_10801_));
 AO21x1_ASAP7_75t_R _30110_ (.A1(_08388_),
    .A2(_10768_),
    .B(_10801_),
    .Y(_03751_));
 NOR2x1_ASAP7_75t_R _30111_ (.A(_01137_),
    .B(_10768_),
    .Y(_10802_));
 AO21x1_ASAP7_75t_R _30112_ (.A1(_08419_),
    .A2(_10768_),
    .B(_10802_),
    .Y(_03752_));
 NOR2x1_ASAP7_75t_R _30113_ (.A(_01171_),
    .B(_10768_),
    .Y(_10803_));
 AO21x1_ASAP7_75t_R _30114_ (.A1(_08451_),
    .A2(_10768_),
    .B(_10803_),
    .Y(_03753_));
 NOR2x1_ASAP7_75t_R _30115_ (.A(_01203_),
    .B(_10768_),
    .Y(_10804_));
 AO21x1_ASAP7_75t_R _30116_ (.A1(_08481_),
    .A2(_10768_),
    .B(_10804_),
    .Y(_03754_));
 NOR2x1_ASAP7_75t_R _30117_ (.A(_01237_),
    .B(_10768_),
    .Y(_10805_));
 AO21x1_ASAP7_75t_R _30118_ (.A1(_08512_),
    .A2(_10768_),
    .B(_10805_),
    .Y(_03755_));
 NOR2x1_ASAP7_75t_R _30119_ (.A(_01269_),
    .B(_10768_),
    .Y(_10806_));
 AO21x1_ASAP7_75t_R _30120_ (.A1(_08545_),
    .A2(_10768_),
    .B(_10806_),
    .Y(_03756_));
 NOR2x1_ASAP7_75t_R _30121_ (.A(_01303_),
    .B(_10768_),
    .Y(_10807_));
 AO21x1_ASAP7_75t_R _30122_ (.A1(_08573_),
    .A2(_10768_),
    .B(_10807_),
    .Y(_03757_));
 AND4x2_ASAP7_75t_R _30123_ (.A(_00323_),
    .B(_00184_),
    .C(_10102_),
    .D(_10334_),
    .Y(_10808_));
 TAPCELL_ASAP7_75t_R PHY_306 ();
 TAPCELL_ASAP7_75t_R PHY_305 ();
 TAPCELL_ASAP7_75t_R PHY_304 ();
 NOR2x1_ASAP7_75t_R _30127_ (.A(_00319_),
    .B(_10808_),
    .Y(_10812_));
 AO21x1_ASAP7_75t_R _30128_ (.A1(_07180_),
    .A2(_10808_),
    .B(_10812_),
    .Y(_03758_));
 NOR2x1_ASAP7_75t_R _30129_ (.A(_00273_),
    .B(net258),
    .Y(_10813_));
 AO21x1_ASAP7_75t_R _30130_ (.A1(_07313_),
    .A2(net258),
    .B(_10813_),
    .Y(_03759_));
 NOR2x1_ASAP7_75t_R _30131_ (.A(_00381_),
    .B(net259),
    .Y(_10814_));
 AO21x1_ASAP7_75t_R _30132_ (.A1(_07398_),
    .A2(net259),
    .B(_10814_),
    .Y(_03760_));
 NOR2x1_ASAP7_75t_R _30133_ (.A(_00412_),
    .B(net258),
    .Y(_10815_));
 AO21x1_ASAP7_75t_R _30134_ (.A1(_07469_),
    .A2(net258),
    .B(_10815_),
    .Y(_03761_));
 NOR2x1_ASAP7_75t_R _30135_ (.A(_00442_),
    .B(_10808_),
    .Y(_10816_));
 AO21x1_ASAP7_75t_R _30136_ (.A1(_07534_),
    .A2(_10808_),
    .B(_10816_),
    .Y(_03762_));
 NOR2x1_ASAP7_75t_R _30137_ (.A(_00472_),
    .B(net259),
    .Y(_10817_));
 AO21x1_ASAP7_75t_R _30138_ (.A1(_07581_),
    .A2(net259),
    .B(_10817_),
    .Y(_03763_));
 NOR2x1_ASAP7_75t_R _30139_ (.A(_00502_),
    .B(_10808_),
    .Y(_10818_));
 AO21x1_ASAP7_75t_R _30140_ (.A1(net253),
    .A2(_10808_),
    .B(_10818_),
    .Y(_03764_));
 NOR2x1_ASAP7_75t_R _30141_ (.A(_00532_),
    .B(net258),
    .Y(_10819_));
 AO21x1_ASAP7_75t_R _30142_ (.A1(_07676_),
    .A2(net258),
    .B(_10819_),
    .Y(_03765_));
 TAPCELL_ASAP7_75t_R PHY_303 ();
 NOR2x1_ASAP7_75t_R _30144_ (.A(_00562_),
    .B(net259),
    .Y(_10821_));
 AO21x1_ASAP7_75t_R _30145_ (.A1(net252),
    .A2(net259),
    .B(_10821_),
    .Y(_03766_));
 NOR2x1_ASAP7_75t_R _30146_ (.A(_00592_),
    .B(_10808_),
    .Y(_10822_));
 AO21x1_ASAP7_75t_R _30147_ (.A1(_07780_),
    .A2(_10808_),
    .B(_10822_),
    .Y(_03767_));
 TAPCELL_ASAP7_75t_R PHY_302 ();
 NOR2x1_ASAP7_75t_R _30149_ (.A(_00622_),
    .B(net258),
    .Y(_10824_));
 AO21x1_ASAP7_75t_R _30150_ (.A1(_07817_),
    .A2(net258),
    .B(_10824_),
    .Y(_03768_));
 NOR2x1_ASAP7_75t_R _30151_ (.A(_00652_),
    .B(net259),
    .Y(_10825_));
 AO21x1_ASAP7_75t_R _30152_ (.A1(_07865_),
    .A2(net259),
    .B(_10825_),
    .Y(_03769_));
 NOR2x1_ASAP7_75t_R _30153_ (.A(_00351_),
    .B(_10808_),
    .Y(_10826_));
 AO21x1_ASAP7_75t_R _30154_ (.A1(_07908_),
    .A2(_10808_),
    .B(_10826_),
    .Y(_03770_));
 NOR2x1_ASAP7_75t_R _30155_ (.A(_00714_),
    .B(net258),
    .Y(_10827_));
 AO21x1_ASAP7_75t_R _30156_ (.A1(_07950_),
    .A2(net258),
    .B(_10827_),
    .Y(_03771_));
 NOR2x1_ASAP7_75t_R _30157_ (.A(_00746_),
    .B(_10808_),
    .Y(_10828_));
 AO21x1_ASAP7_75t_R _30158_ (.A1(_07990_),
    .A2(_10808_),
    .B(_10828_),
    .Y(_03772_));
 NOR2x1_ASAP7_75t_R _30159_ (.A(_00779_),
    .B(net258),
    .Y(_10829_));
 AO21x1_ASAP7_75t_R _30160_ (.A1(_08034_),
    .A2(net258),
    .B(_10829_),
    .Y(_03773_));
 NOR2x1_ASAP7_75t_R _30161_ (.A(_00812_),
    .B(net258),
    .Y(_10830_));
 AO21x1_ASAP7_75t_R _30162_ (.A1(_08073_),
    .A2(net258),
    .B(_10830_),
    .Y(_03774_));
 NOR2x1_ASAP7_75t_R _30163_ (.A(_00845_),
    .B(net258),
    .Y(_10831_));
 AO21x1_ASAP7_75t_R _30164_ (.A1(_08116_),
    .A2(net258),
    .B(_10831_),
    .Y(_03775_));
 TAPCELL_ASAP7_75t_R PHY_301 ();
 NOR2x1_ASAP7_75t_R _30166_ (.A(_00877_),
    .B(net259),
    .Y(_10833_));
 AO21x1_ASAP7_75t_R _30167_ (.A1(net251),
    .A2(net259),
    .B(_10833_),
    .Y(_03776_));
 NOR2x1_ASAP7_75t_R _30168_ (.A(_00910_),
    .B(net259),
    .Y(_10834_));
 AO21x1_ASAP7_75t_R _30169_ (.A1(_08187_),
    .A2(net259),
    .B(_10834_),
    .Y(_03777_));
 TAPCELL_ASAP7_75t_R PHY_300 ();
 NOR2x1_ASAP7_75t_R _30171_ (.A(_00942_),
    .B(net258),
    .Y(_10836_));
 AO21x1_ASAP7_75t_R _30172_ (.A1(_08219_),
    .A2(net258),
    .B(_10836_),
    .Y(_03778_));
 NOR2x1_ASAP7_75t_R _30173_ (.A(_00975_),
    .B(net259),
    .Y(_10837_));
 AO21x1_ASAP7_75t_R _30174_ (.A1(_08254_),
    .A2(net259),
    .B(_10837_),
    .Y(_03779_));
 NOR2x1_ASAP7_75t_R _30175_ (.A(_01007_),
    .B(_10808_),
    .Y(_10838_));
 AO21x1_ASAP7_75t_R _30176_ (.A1(net250),
    .A2(_10808_),
    .B(_10838_),
    .Y(_03780_));
 NOR2x1_ASAP7_75t_R _30177_ (.A(_01041_),
    .B(net259),
    .Y(_10839_));
 AO21x1_ASAP7_75t_R _30178_ (.A1(_08319_),
    .A2(net259),
    .B(_10839_),
    .Y(_03781_));
 NOR2x1_ASAP7_75t_R _30179_ (.A(_01073_),
    .B(net258),
    .Y(_10840_));
 AO21x1_ASAP7_75t_R _30180_ (.A1(_08357_),
    .A2(net258),
    .B(_10840_),
    .Y(_03782_));
 NOR2x1_ASAP7_75t_R _30181_ (.A(_01106_),
    .B(net258),
    .Y(_10841_));
 AO21x1_ASAP7_75t_R _30182_ (.A1(_08388_),
    .A2(net258),
    .B(_10841_),
    .Y(_03783_));
 NOR2x1_ASAP7_75t_R _30183_ (.A(_01138_),
    .B(net258),
    .Y(_10842_));
 AO21x1_ASAP7_75t_R _30184_ (.A1(_08419_),
    .A2(net258),
    .B(_10842_),
    .Y(_03784_));
 NOR2x1_ASAP7_75t_R _30185_ (.A(_01172_),
    .B(net259),
    .Y(_10843_));
 AO21x1_ASAP7_75t_R _30186_ (.A1(_08451_),
    .A2(net259),
    .B(_10843_),
    .Y(_03785_));
 NOR2x1_ASAP7_75t_R _30187_ (.A(_01204_),
    .B(_10808_),
    .Y(_10844_));
 AO21x1_ASAP7_75t_R _30188_ (.A1(_08481_),
    .A2(_10808_),
    .B(_10844_),
    .Y(_03786_));
 NOR2x1_ASAP7_75t_R _30189_ (.A(_01238_),
    .B(net259),
    .Y(_10845_));
 AO21x1_ASAP7_75t_R _30190_ (.A1(_08512_),
    .A2(net259),
    .B(_10845_),
    .Y(_03787_));
 NOR2x1_ASAP7_75t_R _30191_ (.A(_01270_),
    .B(net258),
    .Y(_10846_));
 AO21x1_ASAP7_75t_R _30192_ (.A1(_08545_),
    .A2(net258),
    .B(_10846_),
    .Y(_03788_));
 NOR2x1_ASAP7_75t_R _30193_ (.A(_01304_),
    .B(net259),
    .Y(_10847_));
 AO21x1_ASAP7_75t_R _30194_ (.A1(_08573_),
    .A2(net259),
    .B(_10847_),
    .Y(_03789_));
 AND3x4_ASAP7_75t_R _30195_ (.A(_06882_),
    .B(_10102_),
    .C(_10334_),
    .Y(_10848_));
 TAPCELL_ASAP7_75t_R PHY_299 ();
 TAPCELL_ASAP7_75t_R PHY_298 ();
 TAPCELL_ASAP7_75t_R PHY_297 ();
 NOR2x1_ASAP7_75t_R _30199_ (.A(_00320_),
    .B(_10848_),
    .Y(_10852_));
 AO21x1_ASAP7_75t_R _30200_ (.A1(_07180_),
    .A2(_10848_),
    .B(_10852_),
    .Y(_03790_));
 NOR2x1_ASAP7_75t_R _30201_ (.A(_00274_),
    .B(_10848_),
    .Y(_10853_));
 AO21x1_ASAP7_75t_R _30202_ (.A1(_07313_),
    .A2(_10848_),
    .B(_10853_),
    .Y(_03791_));
 NOR2x1_ASAP7_75t_R _30203_ (.A(_00382_),
    .B(_10848_),
    .Y(_10854_));
 AO21x1_ASAP7_75t_R _30204_ (.A1(_07398_),
    .A2(_10848_),
    .B(_10854_),
    .Y(_03792_));
 NOR2x1_ASAP7_75t_R _30205_ (.A(_00413_),
    .B(_10848_),
    .Y(_10855_));
 AO21x1_ASAP7_75t_R _30206_ (.A1(_07469_),
    .A2(_10848_),
    .B(_10855_),
    .Y(_03793_));
 NOR2x1_ASAP7_75t_R _30207_ (.A(_00443_),
    .B(_10848_),
    .Y(_10856_));
 AO21x1_ASAP7_75t_R _30208_ (.A1(_07534_),
    .A2(_10848_),
    .B(_10856_),
    .Y(_03794_));
 NOR2x1_ASAP7_75t_R _30209_ (.A(_00473_),
    .B(_10848_),
    .Y(_10857_));
 AO21x1_ASAP7_75t_R _30210_ (.A1(_07581_),
    .A2(_10848_),
    .B(_10857_),
    .Y(_03795_));
 NOR2x1_ASAP7_75t_R _30211_ (.A(_00503_),
    .B(_10848_),
    .Y(_10858_));
 AO21x1_ASAP7_75t_R _30212_ (.A1(net253),
    .A2(_10848_),
    .B(_10858_),
    .Y(_03796_));
 NOR2x1_ASAP7_75t_R _30213_ (.A(_00533_),
    .B(_10848_),
    .Y(_10859_));
 AO21x1_ASAP7_75t_R _30214_ (.A1(_07676_),
    .A2(_10848_),
    .B(_10859_),
    .Y(_03797_));
 TAPCELL_ASAP7_75t_R PHY_296 ();
 NOR2x1_ASAP7_75t_R _30216_ (.A(_00563_),
    .B(_10848_),
    .Y(_10861_));
 AO21x1_ASAP7_75t_R _30217_ (.A1(net252),
    .A2(_10848_),
    .B(_10861_),
    .Y(_03798_));
 NOR2x1_ASAP7_75t_R _30218_ (.A(_00593_),
    .B(_10848_),
    .Y(_10862_));
 AO21x1_ASAP7_75t_R _30219_ (.A1(_07780_),
    .A2(_10848_),
    .B(_10862_),
    .Y(_03799_));
 TAPCELL_ASAP7_75t_R PHY_295 ();
 NOR2x1_ASAP7_75t_R _30221_ (.A(_00623_),
    .B(_10848_),
    .Y(_10864_));
 AO21x1_ASAP7_75t_R _30222_ (.A1(_07817_),
    .A2(_10848_),
    .B(_10864_),
    .Y(_03800_));
 NOR2x1_ASAP7_75t_R _30223_ (.A(_00653_),
    .B(_10848_),
    .Y(_10865_));
 AO21x1_ASAP7_75t_R _30224_ (.A1(_07865_),
    .A2(_10848_),
    .B(_10865_),
    .Y(_03801_));
 NOR2x1_ASAP7_75t_R _30225_ (.A(_00352_),
    .B(_10848_),
    .Y(_10866_));
 AO21x1_ASAP7_75t_R _30226_ (.A1(_07908_),
    .A2(_10848_),
    .B(_10866_),
    .Y(_03802_));
 NOR2x1_ASAP7_75t_R _30227_ (.A(_00715_),
    .B(_10848_),
    .Y(_10867_));
 AO21x1_ASAP7_75t_R _30228_ (.A1(_07950_),
    .A2(_10848_),
    .B(_10867_),
    .Y(_03803_));
 NOR2x1_ASAP7_75t_R _30229_ (.A(_00747_),
    .B(_10848_),
    .Y(_10868_));
 AO21x1_ASAP7_75t_R _30230_ (.A1(_07990_),
    .A2(_10848_),
    .B(_10868_),
    .Y(_03804_));
 NOR2x1_ASAP7_75t_R _30231_ (.A(_00780_),
    .B(_10848_),
    .Y(_10869_));
 AO21x1_ASAP7_75t_R _30232_ (.A1(_08034_),
    .A2(_10848_),
    .B(_10869_),
    .Y(_03805_));
 NOR2x1_ASAP7_75t_R _30233_ (.A(_00813_),
    .B(_10848_),
    .Y(_10870_));
 AO21x1_ASAP7_75t_R _30234_ (.A1(_08073_),
    .A2(_10848_),
    .B(_10870_),
    .Y(_03806_));
 NOR2x1_ASAP7_75t_R _30235_ (.A(_00846_),
    .B(_10848_),
    .Y(_10871_));
 AO21x1_ASAP7_75t_R _30236_ (.A1(_08116_),
    .A2(_10848_),
    .B(_10871_),
    .Y(_03807_));
 TAPCELL_ASAP7_75t_R PHY_294 ();
 NOR2x1_ASAP7_75t_R _30238_ (.A(_00878_),
    .B(_10848_),
    .Y(_10873_));
 AO21x1_ASAP7_75t_R _30239_ (.A1(net251),
    .A2(_10848_),
    .B(_10873_),
    .Y(_03808_));
 NOR2x1_ASAP7_75t_R _30240_ (.A(_00911_),
    .B(_10848_),
    .Y(_10874_));
 AO21x1_ASAP7_75t_R _30241_ (.A1(_08187_),
    .A2(_10848_),
    .B(_10874_),
    .Y(_03809_));
 TAPCELL_ASAP7_75t_R PHY_293 ();
 NOR2x1_ASAP7_75t_R _30243_ (.A(_00943_),
    .B(_10848_),
    .Y(_10876_));
 AO21x1_ASAP7_75t_R _30244_ (.A1(_08219_),
    .A2(_10848_),
    .B(_10876_),
    .Y(_03810_));
 NOR2x1_ASAP7_75t_R _30245_ (.A(_00976_),
    .B(_10848_),
    .Y(_10877_));
 AO21x1_ASAP7_75t_R _30246_ (.A1(_08254_),
    .A2(_10848_),
    .B(_10877_),
    .Y(_03811_));
 NOR2x1_ASAP7_75t_R _30247_ (.A(_01008_),
    .B(_10848_),
    .Y(_10878_));
 AO21x1_ASAP7_75t_R _30248_ (.A1(net250),
    .A2(_10848_),
    .B(_10878_),
    .Y(_03812_));
 NOR2x1_ASAP7_75t_R _30249_ (.A(_01042_),
    .B(_10848_),
    .Y(_10879_));
 AO21x1_ASAP7_75t_R _30250_ (.A1(_08319_),
    .A2(_10848_),
    .B(_10879_),
    .Y(_03813_));
 NOR2x1_ASAP7_75t_R _30251_ (.A(_01074_),
    .B(_10848_),
    .Y(_10880_));
 AO21x1_ASAP7_75t_R _30252_ (.A1(_08357_),
    .A2(_10848_),
    .B(_10880_),
    .Y(_03814_));
 NOR2x1_ASAP7_75t_R _30253_ (.A(_01107_),
    .B(_10848_),
    .Y(_10881_));
 AO21x1_ASAP7_75t_R _30254_ (.A1(_08388_),
    .A2(_10848_),
    .B(_10881_),
    .Y(_03815_));
 NOR2x1_ASAP7_75t_R _30255_ (.A(_01139_),
    .B(_10848_),
    .Y(_10882_));
 AO21x1_ASAP7_75t_R _30256_ (.A1(_08419_),
    .A2(_10848_),
    .B(_10882_),
    .Y(_03816_));
 NOR2x1_ASAP7_75t_R _30257_ (.A(_01173_),
    .B(_10848_),
    .Y(_10883_));
 AO21x1_ASAP7_75t_R _30258_ (.A1(_08451_),
    .A2(_10848_),
    .B(_10883_),
    .Y(_03817_));
 NOR2x1_ASAP7_75t_R _30259_ (.A(_01205_),
    .B(_10848_),
    .Y(_10884_));
 AO21x1_ASAP7_75t_R _30260_ (.A1(_08481_),
    .A2(_10848_),
    .B(_10884_),
    .Y(_03818_));
 NOR2x1_ASAP7_75t_R _30261_ (.A(_01239_),
    .B(_10848_),
    .Y(_10885_));
 AO21x1_ASAP7_75t_R _30262_ (.A1(_08512_),
    .A2(_10848_),
    .B(_10885_),
    .Y(_03819_));
 NOR2x1_ASAP7_75t_R _30263_ (.A(_01271_),
    .B(_10848_),
    .Y(_10886_));
 AO21x1_ASAP7_75t_R _30264_ (.A1(_08545_),
    .A2(_10848_),
    .B(_10886_),
    .Y(_03820_));
 NOR2x1_ASAP7_75t_R _30265_ (.A(_01305_),
    .B(_10848_),
    .Y(_10887_));
 AO21x1_ASAP7_75t_R _30266_ (.A1(_08573_),
    .A2(_10848_),
    .B(_10887_),
    .Y(_03821_));
 AND3x4_ASAP7_75t_R _30267_ (.A(_09663_),
    .B(_10102_),
    .C(_10334_),
    .Y(_10888_));
 TAPCELL_ASAP7_75t_R PHY_292 ();
 TAPCELL_ASAP7_75t_R PHY_291 ();
 TAPCELL_ASAP7_75t_R PHY_290 ();
 NOR2x1_ASAP7_75t_R _30271_ (.A(_00321_),
    .B(_10888_),
    .Y(_10892_));
 AO21x1_ASAP7_75t_R _30272_ (.A1(_07180_),
    .A2(_10888_),
    .B(_10892_),
    .Y(_03822_));
 NOR2x1_ASAP7_75t_R _30273_ (.A(_00275_),
    .B(_10888_),
    .Y(_10893_));
 AO21x1_ASAP7_75t_R _30274_ (.A1(_07313_),
    .A2(_10888_),
    .B(_10893_),
    .Y(_03823_));
 NOR2x1_ASAP7_75t_R _30275_ (.A(_00383_),
    .B(_10888_),
    .Y(_10894_));
 AO21x1_ASAP7_75t_R _30276_ (.A1(_07398_),
    .A2(_10888_),
    .B(_10894_),
    .Y(_03824_));
 NOR2x1_ASAP7_75t_R _30277_ (.A(_00414_),
    .B(_10888_),
    .Y(_10895_));
 AO21x1_ASAP7_75t_R _30278_ (.A1(_07469_),
    .A2(_10888_),
    .B(_10895_),
    .Y(_03825_));
 NOR2x1_ASAP7_75t_R _30279_ (.A(_00444_),
    .B(_10888_),
    .Y(_10896_));
 AO21x1_ASAP7_75t_R _30280_ (.A1(_07534_),
    .A2(_10888_),
    .B(_10896_),
    .Y(_03826_));
 NOR2x1_ASAP7_75t_R _30281_ (.A(_00474_),
    .B(_10888_),
    .Y(_10897_));
 AO21x1_ASAP7_75t_R _30282_ (.A1(_07581_),
    .A2(_10888_),
    .B(_10897_),
    .Y(_03827_));
 NOR2x1_ASAP7_75t_R _30283_ (.A(_00504_),
    .B(_10888_),
    .Y(_10898_));
 AO21x1_ASAP7_75t_R _30284_ (.A1(net253),
    .A2(_10888_),
    .B(_10898_),
    .Y(_03828_));
 NOR2x1_ASAP7_75t_R _30285_ (.A(_00534_),
    .B(_10888_),
    .Y(_10899_));
 AO21x1_ASAP7_75t_R _30286_ (.A1(_07676_),
    .A2(_10888_),
    .B(_10899_),
    .Y(_03829_));
 TAPCELL_ASAP7_75t_R PHY_289 ();
 NOR2x1_ASAP7_75t_R _30288_ (.A(_00564_),
    .B(_10888_),
    .Y(_10901_));
 AO21x1_ASAP7_75t_R _30289_ (.A1(net252),
    .A2(_10888_),
    .B(_10901_),
    .Y(_03830_));
 NOR2x1_ASAP7_75t_R _30290_ (.A(_00594_),
    .B(_10888_),
    .Y(_10902_));
 AO21x1_ASAP7_75t_R _30291_ (.A1(_07780_),
    .A2(_10888_),
    .B(_10902_),
    .Y(_03831_));
 TAPCELL_ASAP7_75t_R PHY_288 ();
 NOR2x1_ASAP7_75t_R _30293_ (.A(_00624_),
    .B(_10888_),
    .Y(_10904_));
 AO21x1_ASAP7_75t_R _30294_ (.A1(_07817_),
    .A2(_10888_),
    .B(_10904_),
    .Y(_03832_));
 NOR2x1_ASAP7_75t_R _30295_ (.A(_00654_),
    .B(_10888_),
    .Y(_10905_));
 AO21x1_ASAP7_75t_R _30296_ (.A1(_07865_),
    .A2(_10888_),
    .B(_10905_),
    .Y(_03833_));
 NOR2x1_ASAP7_75t_R _30297_ (.A(_00353_),
    .B(_10888_),
    .Y(_10906_));
 AO21x1_ASAP7_75t_R _30298_ (.A1(_07908_),
    .A2(_10888_),
    .B(_10906_),
    .Y(_03834_));
 NOR2x1_ASAP7_75t_R _30299_ (.A(_00716_),
    .B(_10888_),
    .Y(_10907_));
 AO21x1_ASAP7_75t_R _30300_ (.A1(_07950_),
    .A2(_10888_),
    .B(_10907_),
    .Y(_03835_));
 NOR2x1_ASAP7_75t_R _30301_ (.A(_00748_),
    .B(_10888_),
    .Y(_10908_));
 AO21x1_ASAP7_75t_R _30302_ (.A1(_07990_),
    .A2(_10888_),
    .B(_10908_),
    .Y(_03836_));
 NOR2x1_ASAP7_75t_R _30303_ (.A(_00781_),
    .B(_10888_),
    .Y(_10909_));
 AO21x1_ASAP7_75t_R _30304_ (.A1(_08034_),
    .A2(_10888_),
    .B(_10909_),
    .Y(_03837_));
 NOR2x1_ASAP7_75t_R _30305_ (.A(_00814_),
    .B(_10888_),
    .Y(_10910_));
 AO21x1_ASAP7_75t_R _30306_ (.A1(_08073_),
    .A2(_10888_),
    .B(_10910_),
    .Y(_03838_));
 NOR2x1_ASAP7_75t_R _30307_ (.A(_00847_),
    .B(_10888_),
    .Y(_10911_));
 AO21x1_ASAP7_75t_R _30308_ (.A1(_08116_),
    .A2(_10888_),
    .B(_10911_),
    .Y(_03839_));
 TAPCELL_ASAP7_75t_R PHY_287 ();
 NOR2x1_ASAP7_75t_R _30310_ (.A(_00879_),
    .B(_10888_),
    .Y(_10913_));
 AO21x1_ASAP7_75t_R _30311_ (.A1(net251),
    .A2(_10888_),
    .B(_10913_),
    .Y(_03840_));
 NOR2x1_ASAP7_75t_R _30312_ (.A(_00912_),
    .B(_10888_),
    .Y(_10914_));
 AO21x1_ASAP7_75t_R _30313_ (.A1(_08187_),
    .A2(_10888_),
    .B(_10914_),
    .Y(_03841_));
 TAPCELL_ASAP7_75t_R PHY_286 ();
 NOR2x1_ASAP7_75t_R _30315_ (.A(_00944_),
    .B(_10888_),
    .Y(_10916_));
 AO21x1_ASAP7_75t_R _30316_ (.A1(_08219_),
    .A2(_10888_),
    .B(_10916_),
    .Y(_03842_));
 NOR2x1_ASAP7_75t_R _30317_ (.A(_00977_),
    .B(_10888_),
    .Y(_10917_));
 AO21x1_ASAP7_75t_R _30318_ (.A1(_08254_),
    .A2(_10888_),
    .B(_10917_),
    .Y(_03843_));
 NOR2x1_ASAP7_75t_R _30319_ (.A(_01009_),
    .B(_10888_),
    .Y(_10918_));
 AO21x1_ASAP7_75t_R _30320_ (.A1(net250),
    .A2(_10888_),
    .B(_10918_),
    .Y(_03844_));
 NOR2x1_ASAP7_75t_R _30321_ (.A(_01043_),
    .B(_10888_),
    .Y(_10919_));
 AO21x1_ASAP7_75t_R _30322_ (.A1(_08319_),
    .A2(_10888_),
    .B(_10919_),
    .Y(_03845_));
 NOR2x1_ASAP7_75t_R _30323_ (.A(_01075_),
    .B(_10888_),
    .Y(_10920_));
 AO21x1_ASAP7_75t_R _30324_ (.A1(_08357_),
    .A2(_10888_),
    .B(_10920_),
    .Y(_03846_));
 NOR2x1_ASAP7_75t_R _30325_ (.A(_01108_),
    .B(_10888_),
    .Y(_10921_));
 AO21x1_ASAP7_75t_R _30326_ (.A1(_08388_),
    .A2(_10888_),
    .B(_10921_),
    .Y(_03847_));
 NOR2x1_ASAP7_75t_R _30327_ (.A(_01140_),
    .B(_10888_),
    .Y(_10922_));
 AO21x1_ASAP7_75t_R _30328_ (.A1(_08419_),
    .A2(_10888_),
    .B(_10922_),
    .Y(_03848_));
 NOR2x1_ASAP7_75t_R _30329_ (.A(_01174_),
    .B(_10888_),
    .Y(_10923_));
 AO21x1_ASAP7_75t_R _30330_ (.A1(_08451_),
    .A2(_10888_),
    .B(_10923_),
    .Y(_03849_));
 NOR2x1_ASAP7_75t_R _30331_ (.A(_01206_),
    .B(_10888_),
    .Y(_10924_));
 AO21x1_ASAP7_75t_R _30332_ (.A1(_08481_),
    .A2(_10888_),
    .B(_10924_),
    .Y(_03850_));
 NOR2x1_ASAP7_75t_R _30333_ (.A(_01240_),
    .B(_10888_),
    .Y(_10925_));
 AO21x1_ASAP7_75t_R _30334_ (.A1(_08512_),
    .A2(_10888_),
    .B(_10925_),
    .Y(_03851_));
 NOR2x1_ASAP7_75t_R _30335_ (.A(_01272_),
    .B(_10888_),
    .Y(_10926_));
 AO21x1_ASAP7_75t_R _30336_ (.A1(_08545_),
    .A2(_10888_),
    .B(_10926_),
    .Y(_03852_));
 NOR2x1_ASAP7_75t_R _30337_ (.A(_01306_),
    .B(_10888_),
    .Y(_10927_));
 AO21x1_ASAP7_75t_R _30338_ (.A1(_08573_),
    .A2(_10888_),
    .B(_10927_),
    .Y(_03853_));
 AND3x4_ASAP7_75t_R _30339_ (.A(_09736_),
    .B(_10102_),
    .C(_10334_),
    .Y(_10928_));
 TAPCELL_ASAP7_75t_R PHY_285 ();
 TAPCELL_ASAP7_75t_R PHY_284 ();
 TAPCELL_ASAP7_75t_R PHY_283 ();
 NOR2x1_ASAP7_75t_R _30343_ (.A(_00322_),
    .B(_10928_),
    .Y(_10932_));
 AO21x1_ASAP7_75t_R _30344_ (.A1(_07180_),
    .A2(_10928_),
    .B(_10932_),
    .Y(_03854_));
 NOR2x1_ASAP7_75t_R _30345_ (.A(_00276_),
    .B(_10928_),
    .Y(_10933_));
 AO21x1_ASAP7_75t_R _30346_ (.A1(_07313_),
    .A2(_10928_),
    .B(_10933_),
    .Y(_03855_));
 NOR2x1_ASAP7_75t_R _30347_ (.A(_00384_),
    .B(_10928_),
    .Y(_10934_));
 AO21x1_ASAP7_75t_R _30348_ (.A1(_07398_),
    .A2(_10928_),
    .B(_10934_),
    .Y(_03856_));
 NOR2x1_ASAP7_75t_R _30349_ (.A(_00415_),
    .B(_10928_),
    .Y(_10935_));
 AO21x1_ASAP7_75t_R _30350_ (.A1(_07469_),
    .A2(_10928_),
    .B(_10935_),
    .Y(_03857_));
 NOR2x1_ASAP7_75t_R _30351_ (.A(_00445_),
    .B(_10928_),
    .Y(_10936_));
 AO21x1_ASAP7_75t_R _30352_ (.A1(_07534_),
    .A2(_10928_),
    .B(_10936_),
    .Y(_03858_));
 NOR2x1_ASAP7_75t_R _30353_ (.A(_00475_),
    .B(_10928_),
    .Y(_10937_));
 AO21x1_ASAP7_75t_R _30354_ (.A1(_07581_),
    .A2(_10928_),
    .B(_10937_),
    .Y(_03859_));
 NOR2x1_ASAP7_75t_R _30355_ (.A(_00505_),
    .B(_10928_),
    .Y(_10938_));
 AO21x1_ASAP7_75t_R _30356_ (.A1(net253),
    .A2(_10928_),
    .B(_10938_),
    .Y(_03860_));
 NOR2x1_ASAP7_75t_R _30357_ (.A(_00535_),
    .B(_10928_),
    .Y(_10939_));
 AO21x1_ASAP7_75t_R _30358_ (.A1(_07676_),
    .A2(_10928_),
    .B(_10939_),
    .Y(_03861_));
 TAPCELL_ASAP7_75t_R PHY_282 ();
 NOR2x1_ASAP7_75t_R _30360_ (.A(_00565_),
    .B(_10928_),
    .Y(_10941_));
 AO21x1_ASAP7_75t_R _30361_ (.A1(net252),
    .A2(_10928_),
    .B(_10941_),
    .Y(_03862_));
 NOR2x1_ASAP7_75t_R _30362_ (.A(_00595_),
    .B(_10928_),
    .Y(_10942_));
 AO21x1_ASAP7_75t_R _30363_ (.A1(_07780_),
    .A2(_10928_),
    .B(_10942_),
    .Y(_03863_));
 TAPCELL_ASAP7_75t_R PHY_281 ();
 NOR2x1_ASAP7_75t_R _30365_ (.A(_00625_),
    .B(_10928_),
    .Y(_10944_));
 AO21x1_ASAP7_75t_R _30366_ (.A1(_07817_),
    .A2(_10928_),
    .B(_10944_),
    .Y(_03864_));
 NOR2x1_ASAP7_75t_R _30367_ (.A(_00655_),
    .B(_10928_),
    .Y(_10945_));
 AO21x1_ASAP7_75t_R _30368_ (.A1(_07865_),
    .A2(_10928_),
    .B(_10945_),
    .Y(_03865_));
 NOR2x1_ASAP7_75t_R _30369_ (.A(_00354_),
    .B(_10928_),
    .Y(_10946_));
 AO21x1_ASAP7_75t_R _30370_ (.A1(_07908_),
    .A2(_10928_),
    .B(_10946_),
    .Y(_03866_));
 NOR2x1_ASAP7_75t_R _30371_ (.A(_00717_),
    .B(_10928_),
    .Y(_10947_));
 AO21x1_ASAP7_75t_R _30372_ (.A1(_07950_),
    .A2(_10928_),
    .B(_10947_),
    .Y(_03867_));
 NOR2x1_ASAP7_75t_R _30373_ (.A(_00749_),
    .B(_10928_),
    .Y(_10948_));
 AO21x1_ASAP7_75t_R _30374_ (.A1(_07990_),
    .A2(_10928_),
    .B(_10948_),
    .Y(_03868_));
 NOR2x1_ASAP7_75t_R _30375_ (.A(_00782_),
    .B(_10928_),
    .Y(_10949_));
 AO21x1_ASAP7_75t_R _30376_ (.A1(_08034_),
    .A2(_10928_),
    .B(_10949_),
    .Y(_03869_));
 NOR2x1_ASAP7_75t_R _30377_ (.A(_00815_),
    .B(_10928_),
    .Y(_10950_));
 AO21x1_ASAP7_75t_R _30378_ (.A1(_08073_),
    .A2(_10928_),
    .B(_10950_),
    .Y(_03870_));
 NOR2x1_ASAP7_75t_R _30379_ (.A(_00848_),
    .B(_10928_),
    .Y(_10951_));
 AO21x1_ASAP7_75t_R _30380_ (.A1(_08116_),
    .A2(_10928_),
    .B(_10951_),
    .Y(_03871_));
 TAPCELL_ASAP7_75t_R PHY_280 ();
 NOR2x1_ASAP7_75t_R _30382_ (.A(_00880_),
    .B(_10928_),
    .Y(_10953_));
 AO21x1_ASAP7_75t_R _30383_ (.A1(net251),
    .A2(_10928_),
    .B(_10953_),
    .Y(_03872_));
 NOR2x1_ASAP7_75t_R _30384_ (.A(_00913_),
    .B(_10928_),
    .Y(_10954_));
 AO21x1_ASAP7_75t_R _30385_ (.A1(_08187_),
    .A2(_10928_),
    .B(_10954_),
    .Y(_03873_));
 TAPCELL_ASAP7_75t_R PHY_279 ();
 NOR2x1_ASAP7_75t_R _30387_ (.A(_00945_),
    .B(_10928_),
    .Y(_10956_));
 AO21x1_ASAP7_75t_R _30388_ (.A1(_08219_),
    .A2(_10928_),
    .B(_10956_),
    .Y(_03874_));
 NOR2x1_ASAP7_75t_R _30389_ (.A(_00978_),
    .B(_10928_),
    .Y(_10957_));
 AO21x1_ASAP7_75t_R _30390_ (.A1(_08254_),
    .A2(_10928_),
    .B(_10957_),
    .Y(_03875_));
 NOR2x1_ASAP7_75t_R _30391_ (.A(_01010_),
    .B(_10928_),
    .Y(_10958_));
 AO21x1_ASAP7_75t_R _30392_ (.A1(net250),
    .A2(_10928_),
    .B(_10958_),
    .Y(_03876_));
 NOR2x1_ASAP7_75t_R _30393_ (.A(_01044_),
    .B(_10928_),
    .Y(_10959_));
 AO21x1_ASAP7_75t_R _30394_ (.A1(_08319_),
    .A2(_10928_),
    .B(_10959_),
    .Y(_03877_));
 NOR2x1_ASAP7_75t_R _30395_ (.A(_01076_),
    .B(_10928_),
    .Y(_10960_));
 AO21x1_ASAP7_75t_R _30396_ (.A1(_08357_),
    .A2(_10928_),
    .B(_10960_),
    .Y(_03878_));
 NOR2x1_ASAP7_75t_R _30397_ (.A(_01109_),
    .B(_10928_),
    .Y(_10961_));
 AO21x1_ASAP7_75t_R _30398_ (.A1(_08388_),
    .A2(_10928_),
    .B(_10961_),
    .Y(_03879_));
 NOR2x1_ASAP7_75t_R _30399_ (.A(_01141_),
    .B(_10928_),
    .Y(_10962_));
 AO21x1_ASAP7_75t_R _30400_ (.A1(_08419_),
    .A2(_10928_),
    .B(_10962_),
    .Y(_03880_));
 NOR2x1_ASAP7_75t_R _30401_ (.A(_01175_),
    .B(_10928_),
    .Y(_10963_));
 AO21x1_ASAP7_75t_R _30402_ (.A1(_08451_),
    .A2(_10928_),
    .B(_10963_),
    .Y(_03881_));
 NOR2x1_ASAP7_75t_R _30403_ (.A(_01207_),
    .B(_10928_),
    .Y(_10964_));
 AO21x1_ASAP7_75t_R _30404_ (.A1(_08481_),
    .A2(_10928_),
    .B(_10964_),
    .Y(_03882_));
 NOR2x1_ASAP7_75t_R _30405_ (.A(_01241_),
    .B(_10928_),
    .Y(_10965_));
 AO21x1_ASAP7_75t_R _30406_ (.A1(_08512_),
    .A2(_10928_),
    .B(_10965_),
    .Y(_03883_));
 NOR2x1_ASAP7_75t_R _30407_ (.A(_01273_),
    .B(_10928_),
    .Y(_10966_));
 AO21x1_ASAP7_75t_R _30408_ (.A1(_08545_),
    .A2(_10928_),
    .B(_10966_),
    .Y(_03884_));
 NOR2x1_ASAP7_75t_R _30409_ (.A(_01307_),
    .B(_10928_),
    .Y(_10967_));
 AO21x1_ASAP7_75t_R _30410_ (.A1(_08573_),
    .A2(_10928_),
    .B(_10967_),
    .Y(_03885_));
 AND5x1_ASAP7_75t_R _30411_ (.A(_13325_),
    .B(_00282_),
    .C(_05778_),
    .D(_13313_),
    .E(_05517_),
    .Y(_10968_));
 NAND2x1_ASAP7_75t_R _30412_ (.A(_05757_),
    .B(_10968_),
    .Y(_10969_));
 NAND2x1_ASAP7_75t_R _30413_ (.A(_01519_),
    .B(_10969_),
    .Y(_10970_));
 OA21x2_ASAP7_75t_R _30414_ (.A1(_05777_),
    .A2(_10969_),
    .B(_10970_),
    .Y(_03886_));
 AND2x2_ASAP7_75t_R _30415_ (.A(_13777_),
    .B(_14501_),
    .Y(_10971_));
 AO21x1_ASAP7_75t_R _30416_ (.A1(_02289_),
    .A2(_18108_),
    .B(_10971_),
    .Y(_10972_));
 AO22x2_ASAP7_75t_R _30417_ (.A1(_18108_),
    .A2(_07176_),
    .B1(_10972_),
    .B2(_02286_),
    .Y(_10973_));
 INVx3_ASAP7_75t_R _30418_ (.A(_10973_),
    .Y(_10974_));
 AND2x4_ASAP7_75t_R _30419_ (.A(_05667_),
    .B(_05661_),
    .Y(_10975_));
 OR2x6_ASAP7_75t_R _30420_ (.A(_05668_),
    .B(_10975_),
    .Y(_10976_));
 TAPCELL_ASAP7_75t_R PHY_278 ();
 AND3x4_ASAP7_75t_R _30422_ (.A(_05582_),
    .B(_09353_),
    .C(_10976_),
    .Y(_10978_));
 TAPCELL_ASAP7_75t_R PHY_277 ();
 TAPCELL_ASAP7_75t_R PHY_276 ();
 AND2x2_ASAP7_75t_R _30425_ (.A(_05586_),
    .B(_05600_),
    .Y(_10981_));
 AND3x4_ASAP7_75t_R _30426_ (.A(_05582_),
    .B(_09364_),
    .C(_09351_),
    .Y(_10982_));
 OAI21x1_ASAP7_75t_R _30427_ (.A1(_10981_),
    .A2(_10975_),
    .B(_10982_),
    .Y(_10983_));
 AOI22x1_ASAP7_75t_R _30428_ (.A1(_10981_),
    .A2(_10982_),
    .B1(_10983_),
    .B2(_00661_),
    .Y(_10984_));
 AO21x1_ASAP7_75t_R _30429_ (.A1(_10974_),
    .A2(_10978_),
    .B(_10984_),
    .Y(_10985_));
 NAND3x2_ASAP7_75t_R _30430_ (.B(_09353_),
    .C(_10976_),
    .Y(_10986_),
    .A(_05582_));
 TAPCELL_ASAP7_75t_R PHY_275 ();
 AO22x2_ASAP7_75t_R _30432_ (.A1(_10981_),
    .A2(_10982_),
    .B1(_10983_),
    .B2(_00661_),
    .Y(_10988_));
 OA211x2_ASAP7_75t_R _30433_ (.A1(_10974_),
    .A2(_10986_),
    .B(_00659_),
    .C(_10988_),
    .Y(_10989_));
 AO21x1_ASAP7_75t_R _30434_ (.A1(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .A2(_10985_),
    .B(_10989_),
    .Y(_03887_));
 TAPCELL_ASAP7_75t_R PHY_274 ();
 NAND2x1_ASAP7_75t_R _30436_ (.A(_02456_),
    .B(_10983_),
    .Y(_10991_));
 OA211x2_ASAP7_75t_R _30437_ (.A1(_09363_),
    .A2(_10986_),
    .B(_10991_),
    .C(_10988_),
    .Y(_10992_));
 AO21x1_ASAP7_75t_R _30438_ (.A1(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .A2(_10984_),
    .B(_10992_),
    .Y(_03888_));
 TAPCELL_ASAP7_75t_R PHY_273 ();
 TAPCELL_ASAP7_75t_R PHY_272 ();
 NAND2x1_ASAP7_75t_R _30441_ (.A(_09390_),
    .B(_10978_),
    .Y(_10995_));
 TAPCELL_ASAP7_75t_R PHY_271 ();
 OA211x2_ASAP7_75t_R _30443_ (.A1(_02458_),
    .A2(_10978_),
    .B(_10995_),
    .C(_10988_),
    .Y(_10997_));
 AOI21x1_ASAP7_75t_R _30444_ (.A1(_01517_),
    .A2(_10984_),
    .B(_10997_),
    .Y(_03889_));
 TAPCELL_ASAP7_75t_R PHY_270 ();
 TAPCELL_ASAP7_75t_R PHY_269 ();
 AO21x1_ASAP7_75t_R _30447_ (.A1(_02457_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11000_));
 TAPCELL_ASAP7_75t_R PHY_268 ();
 OR3x1_ASAP7_75t_R _30449_ (.A(_01516_),
    .B(_02457_),
    .C(_10978_),
    .Y(_11002_));
 OR2x2_ASAP7_75t_R _30450_ (.A(_09397_),
    .B(_10986_),
    .Y(_11003_));
 AOI21x1_ASAP7_75t_R _30451_ (.A1(_11002_),
    .A2(_11003_),
    .B(_10984_),
    .Y(_11004_));
 AOI21x1_ASAP7_75t_R _30452_ (.A1(_01516_),
    .A2(_11000_),
    .B(_11004_),
    .Y(_03890_));
 NAND2x1_ASAP7_75t_R _30453_ (.A(_09408_),
    .B(_10978_),
    .Y(_11005_));
 OA211x2_ASAP7_75t_R _30454_ (.A1(_02460_),
    .A2(_10978_),
    .B(_11005_),
    .C(_10988_),
    .Y(_11006_));
 AOI21x1_ASAP7_75t_R _30455_ (.A1(_01515_),
    .A2(_10984_),
    .B(_11006_),
    .Y(_03891_));
 TAPCELL_ASAP7_75t_R PHY_267 ();
 AO21x1_ASAP7_75t_R _30457_ (.A1(_02459_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11008_));
 OR3x1_ASAP7_75t_R _30458_ (.A(_01514_),
    .B(_02459_),
    .C(_10978_),
    .Y(_11009_));
 INVx2_ASAP7_75t_R _30459_ (.A(_09417_),
    .Y(_11010_));
 NAND2x1_ASAP7_75t_R _30460_ (.A(_11010_),
    .B(_10978_),
    .Y(_11011_));
 AOI21x1_ASAP7_75t_R _30461_ (.A1(_11009_),
    .A2(_11011_),
    .B(_10984_),
    .Y(_11012_));
 AOI21x1_ASAP7_75t_R _30462_ (.A1(_01514_),
    .A2(_11008_),
    .B(_11012_),
    .Y(_03892_));
 NAND2x1_ASAP7_75t_R _30463_ (.A(_09426_),
    .B(_10978_),
    .Y(_11013_));
 OA211x2_ASAP7_75t_R _30464_ (.A1(_02462_),
    .A2(_10978_),
    .B(_11013_),
    .C(_10988_),
    .Y(_11014_));
 AOI21x1_ASAP7_75t_R _30465_ (.A1(_01513_),
    .A2(_10984_),
    .B(_11014_),
    .Y(_03893_));
 TAPCELL_ASAP7_75t_R PHY_266 ();
 TAPCELL_ASAP7_75t_R PHY_265 ();
 OR3x1_ASAP7_75t_R _30468_ (.A(_01512_),
    .B(_02461_),
    .C(_10978_),
    .Y(_11017_));
 OAI21x1_ASAP7_75t_R _30469_ (.A1(_09432_),
    .A2(_10986_),
    .B(_11017_),
    .Y(_11018_));
 AO21x1_ASAP7_75t_R _30470_ (.A1(_02461_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11019_));
 AOI22x1_ASAP7_75t_R _30471_ (.A1(_10988_),
    .A2(_11018_),
    .B1(_11019_),
    .B2(_01512_),
    .Y(_03894_));
 NAND3x2_ASAP7_75t_R _30472_ (.B(_09365_),
    .C(_10976_),
    .Y(_11020_),
    .A(_05582_));
 INVx2_ASAP7_75t_R _30473_ (.A(_11020_),
    .Y(_11021_));
 NAND2x1_ASAP7_75t_R _30474_ (.A(_09438_),
    .B(_11021_),
    .Y(_11022_));
 OA211x2_ASAP7_75t_R _30475_ (.A1(_02464_),
    .A2(_10978_),
    .B(_11022_),
    .C(_10988_),
    .Y(_11023_));
 AOI21x1_ASAP7_75t_R _30476_ (.A1(_01511_),
    .A2(_10984_),
    .B(_11023_),
    .Y(_03895_));
 AO21x1_ASAP7_75t_R _30477_ (.A1(_02463_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11024_));
 OR3x1_ASAP7_75t_R _30478_ (.A(_01510_),
    .B(_02463_),
    .C(_10978_),
    .Y(_11025_));
 OR2x2_ASAP7_75t_R _30479_ (.A(_09445_),
    .B(_10986_),
    .Y(_11026_));
 AOI21x1_ASAP7_75t_R _30480_ (.A1(_11025_),
    .A2(_11026_),
    .B(_10984_),
    .Y(_11027_));
 AOI21x1_ASAP7_75t_R _30481_ (.A1(_01510_),
    .A2(_11024_),
    .B(_11027_),
    .Y(_03896_));
 NAND2x1_ASAP7_75t_R _30482_ (.A(_09452_),
    .B(_10978_),
    .Y(_11028_));
 OA211x2_ASAP7_75t_R _30483_ (.A1(_02466_),
    .A2(_10978_),
    .B(_11028_),
    .C(_10988_),
    .Y(_11029_));
 AOI21x1_ASAP7_75t_R _30484_ (.A1(_01509_),
    .A2(_10984_),
    .B(_11029_),
    .Y(_03897_));
 TAPCELL_ASAP7_75t_R PHY_264 ();
 OR3x1_ASAP7_75t_R _30486_ (.A(_01508_),
    .B(_02465_),
    .C(_10978_),
    .Y(_11031_));
 OAI21x1_ASAP7_75t_R _30487_ (.A1(_09458_),
    .A2(_10986_),
    .B(_11031_),
    .Y(_11032_));
 AO21x1_ASAP7_75t_R _30488_ (.A1(_02465_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11033_));
 AOI22x1_ASAP7_75t_R _30489_ (.A1(_10988_),
    .A2(_11032_),
    .B1(_11033_),
    .B2(_01508_),
    .Y(_03898_));
 TAPCELL_ASAP7_75t_R PHY_263 ();
 NAND2x1_ASAP7_75t_R _30491_ (.A(_09465_),
    .B(_10978_),
    .Y(_11035_));
 OA211x2_ASAP7_75t_R _30492_ (.A1(_02468_),
    .A2(_10978_),
    .B(_11035_),
    .C(_10988_),
    .Y(_11036_));
 AOI21x1_ASAP7_75t_R _30493_ (.A1(_01507_),
    .A2(_10984_),
    .B(_11036_),
    .Y(_03899_));
 OR3x1_ASAP7_75t_R _30494_ (.A(_01506_),
    .B(_02467_),
    .C(_10978_),
    .Y(_11037_));
 OAI21x1_ASAP7_75t_R _30495_ (.A1(_09473_),
    .A2(_10986_),
    .B(_11037_),
    .Y(_11038_));
 AO21x1_ASAP7_75t_R _30496_ (.A1(_02467_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11039_));
 AOI22x1_ASAP7_75t_R _30497_ (.A1(_10988_),
    .A2(_11038_),
    .B1(_11039_),
    .B2(_01506_),
    .Y(_03900_));
 NAND2x1_ASAP7_75t_R _30498_ (.A(_09481_),
    .B(_10978_),
    .Y(_11040_));
 OA211x2_ASAP7_75t_R _30499_ (.A1(_02470_),
    .A2(_10978_),
    .B(_11040_),
    .C(_10988_),
    .Y(_11041_));
 AOI21x1_ASAP7_75t_R _30500_ (.A1(_01505_),
    .A2(_10984_),
    .B(_11041_),
    .Y(_03901_));
 AO21x1_ASAP7_75t_R _30501_ (.A1(_02469_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11042_));
 OR3x1_ASAP7_75t_R _30502_ (.A(_01504_),
    .B(_02469_),
    .C(_10978_),
    .Y(_11043_));
 OR2x2_ASAP7_75t_R _30503_ (.A(_09488_),
    .B(_10986_),
    .Y(_11044_));
 AOI21x1_ASAP7_75t_R _30504_ (.A1(_11043_),
    .A2(_11044_),
    .B(_10984_),
    .Y(_11045_));
 AOI21x1_ASAP7_75t_R _30505_ (.A1(_01504_),
    .A2(_11042_),
    .B(_11045_),
    .Y(_03902_));
 NAND2x1_ASAP7_75t_R _30506_ (.A(_09496_),
    .B(_10978_),
    .Y(_11046_));
 OA211x2_ASAP7_75t_R _30507_ (.A1(_02472_),
    .A2(_10978_),
    .B(_11046_),
    .C(_10988_),
    .Y(_11047_));
 AOI21x1_ASAP7_75t_R _30508_ (.A1(_01503_),
    .A2(_10984_),
    .B(_11047_),
    .Y(_03903_));
 OR3x1_ASAP7_75t_R _30509_ (.A(_01502_),
    .B(_02471_),
    .C(_10978_),
    .Y(_11048_));
 OAI21x1_ASAP7_75t_R _30510_ (.A1(_09503_),
    .A2(_10986_),
    .B(_11048_),
    .Y(_11049_));
 TAPCELL_ASAP7_75t_R PHY_262 ();
 AO21x1_ASAP7_75t_R _30512_ (.A1(_02471_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11051_));
 AOI22x1_ASAP7_75t_R _30513_ (.A1(_10988_),
    .A2(_11049_),
    .B1(_11051_),
    .B2(_01502_),
    .Y(_03904_));
 NAND2x1_ASAP7_75t_R _30514_ (.A(_09512_),
    .B(_10978_),
    .Y(_11052_));
 OA211x2_ASAP7_75t_R _30515_ (.A1(_02474_),
    .A2(_10978_),
    .B(_11052_),
    .C(_10988_),
    .Y(_11053_));
 AOI21x1_ASAP7_75t_R _30516_ (.A1(_01501_),
    .A2(_10984_),
    .B(_11053_),
    .Y(_03905_));
 TAPCELL_ASAP7_75t_R PHY_261 ();
 NOR2x1_ASAP7_75t_R _30518_ (.A(_01500_),
    .B(_02473_),
    .Y(_11055_));
 NOR2x1_ASAP7_75t_R _30519_ (.A(_09519_),
    .B(_10986_),
    .Y(_11056_));
 AO21x1_ASAP7_75t_R _30520_ (.A1(_10986_),
    .A2(_11055_),
    .B(_11056_),
    .Y(_11057_));
 AO21x1_ASAP7_75t_R _30521_ (.A1(_02473_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11058_));
 AOI22x1_ASAP7_75t_R _30522_ (.A1(_10988_),
    .A2(_11057_),
    .B1(_11058_),
    .B2(_01500_),
    .Y(_03906_));
 TAPCELL_ASAP7_75t_R PHY_260 ();
 NAND2x1_ASAP7_75t_R _30524_ (.A(_09526_),
    .B(_10978_),
    .Y(_11060_));
 OA211x2_ASAP7_75t_R _30525_ (.A1(_02476_),
    .A2(_10978_),
    .B(_11060_),
    .C(_10988_),
    .Y(_11061_));
 AOI21x1_ASAP7_75t_R _30526_ (.A1(_01499_),
    .A2(_10984_),
    .B(_11061_),
    .Y(_03907_));
 NOR2x1_ASAP7_75t_R _30527_ (.A(_01498_),
    .B(_02475_),
    .Y(_11062_));
 NOR2x1_ASAP7_75t_R _30528_ (.A(_09532_),
    .B(_10986_),
    .Y(_11063_));
 AO21x1_ASAP7_75t_R _30529_ (.A1(_10986_),
    .A2(_11062_),
    .B(_11063_),
    .Y(_11064_));
 AO21x1_ASAP7_75t_R _30530_ (.A1(_02475_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11065_));
 AOI22x1_ASAP7_75t_R _30531_ (.A1(_10988_),
    .A2(_11064_),
    .B1(_11065_),
    .B2(_01498_),
    .Y(_03908_));
 NAND2x1_ASAP7_75t_R _30532_ (.A(_09539_),
    .B(_11021_),
    .Y(_11066_));
 OA211x2_ASAP7_75t_R _30533_ (.A1(_02478_),
    .A2(_10978_),
    .B(_11066_),
    .C(_10988_),
    .Y(_11067_));
 AOI21x1_ASAP7_75t_R _30534_ (.A1(_01497_),
    .A2(_10984_),
    .B(_11067_),
    .Y(_03909_));
 OR3x1_ASAP7_75t_R _30535_ (.A(_01496_),
    .B(_02477_),
    .C(_10978_),
    .Y(_11068_));
 OAI21x1_ASAP7_75t_R _30536_ (.A1(_09545_),
    .A2(_10986_),
    .B(_11068_),
    .Y(_11069_));
 AO21x1_ASAP7_75t_R _30537_ (.A1(_02477_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11070_));
 AOI22x1_ASAP7_75t_R _30538_ (.A1(_10988_),
    .A2(_11069_),
    .B1(_11070_),
    .B2(_01496_),
    .Y(_03910_));
 OR2x2_ASAP7_75t_R _30539_ (.A(_02480_),
    .B(_10978_),
    .Y(_11071_));
 OA211x2_ASAP7_75t_R _30540_ (.A1(_09560_),
    .A2(_11020_),
    .B(_11071_),
    .C(_10988_),
    .Y(_11072_));
 AOI21x1_ASAP7_75t_R _30541_ (.A1(_01495_),
    .A2(_10984_),
    .B(_11072_),
    .Y(_03911_));
 OR3x1_ASAP7_75t_R _30542_ (.A(_01494_),
    .B(_02479_),
    .C(_10978_),
    .Y(_11073_));
 OAI21x1_ASAP7_75t_R _30543_ (.A1(_09565_),
    .A2(_10986_),
    .B(_11073_),
    .Y(_11074_));
 AO21x1_ASAP7_75t_R _30544_ (.A1(_02479_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11075_));
 AOI22x1_ASAP7_75t_R _30545_ (.A1(_10988_),
    .A2(_11074_),
    .B1(_11075_),
    .B2(_01494_),
    .Y(_03912_));
 NAND2x1_ASAP7_75t_R _30546_ (.A(_09572_),
    .B(_11021_),
    .Y(_11076_));
 OA211x2_ASAP7_75t_R _30547_ (.A1(_02482_),
    .A2(_10978_),
    .B(_11076_),
    .C(_10988_),
    .Y(_11077_));
 AOI21x1_ASAP7_75t_R _30548_ (.A1(_01493_),
    .A2(_10984_),
    .B(_11077_),
    .Y(_03913_));
 OR3x1_ASAP7_75t_R _30549_ (.A(_01492_),
    .B(_02481_),
    .C(_10978_),
    .Y(_11078_));
 OAI21x1_ASAP7_75t_R _30550_ (.A1(_09578_),
    .A2(_10986_),
    .B(_11078_),
    .Y(_11079_));
 AO21x1_ASAP7_75t_R _30551_ (.A1(_02481_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11080_));
 AOI22x1_ASAP7_75t_R _30552_ (.A1(_10988_),
    .A2(_11079_),
    .B1(_11080_),
    .B2(_01492_),
    .Y(_03914_));
 NAND2x1_ASAP7_75t_R _30553_ (.A(_09585_),
    .B(_10978_),
    .Y(_11081_));
 OA211x2_ASAP7_75t_R _30554_ (.A1(_02484_),
    .A2(_10978_),
    .B(_11081_),
    .C(_10988_),
    .Y(_11082_));
 AOI21x1_ASAP7_75t_R _30555_ (.A1(_01491_),
    .A2(_10984_),
    .B(_11082_),
    .Y(_03915_));
 AO21x1_ASAP7_75t_R _30556_ (.A1(_02483_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11083_));
 OR3x1_ASAP7_75t_R _30557_ (.A(_01490_),
    .B(_02483_),
    .C(_10978_),
    .Y(_11084_));
 OR2x2_ASAP7_75t_R _30558_ (.A(_09591_),
    .B(_10986_),
    .Y(_11085_));
 AOI21x1_ASAP7_75t_R _30559_ (.A1(_11084_),
    .A2(_11085_),
    .B(_10984_),
    .Y(_11086_));
 AOI21x1_ASAP7_75t_R _30560_ (.A1(_01490_),
    .A2(_11083_),
    .B(_11086_),
    .Y(_03916_));
 NAND2x1_ASAP7_75t_R _30561_ (.A(_09598_),
    .B(_10978_),
    .Y(_11087_));
 OA211x2_ASAP7_75t_R _30562_ (.A1(_02486_),
    .A2(_10978_),
    .B(_11087_),
    .C(_10988_),
    .Y(_11088_));
 AOI21x1_ASAP7_75t_R _30563_ (.A1(_01489_),
    .A2(_10984_),
    .B(_11088_),
    .Y(_03917_));
 OR3x1_ASAP7_75t_R _30564_ (.A(_01488_),
    .B(_02485_),
    .C(_10978_),
    .Y(_11089_));
 OAI21x1_ASAP7_75t_R _30565_ (.A1(_09605_),
    .A2(_10986_),
    .B(_11089_),
    .Y(_11090_));
 AO21x1_ASAP7_75t_R _30566_ (.A1(_02485_),
    .A2(_10986_),
    .B(_10984_),
    .Y(_11091_));
 AOI22x1_ASAP7_75t_R _30567_ (.A1(_10988_),
    .A2(_11090_),
    .B1(_11091_),
    .B2(_01488_),
    .Y(_03918_));
 AND5x2_ASAP7_75t_R _30568_ (.A(_13302_),
    .B(net289),
    .C(_13955_),
    .D(_05542_),
    .E(_09351_),
    .Y(_11092_));
 AND3x1_ASAP7_75t_R _30569_ (.A(_14083_),
    .B(_06884_),
    .C(_11092_),
    .Y(_11093_));
 AND4x1_ASAP7_75t_R _30570_ (.A(_01315_),
    .B(_05729_),
    .C(_05525_),
    .D(_05723_),
    .Y(_11094_));
 OA211x2_ASAP7_75t_R _30571_ (.A1(_05558_),
    .A2(_06915_),
    .B(_11094_),
    .C(_06594_),
    .Y(_11095_));
 NAND2x1_ASAP7_75t_R _30572_ (.A(_10975_),
    .B(_11092_),
    .Y(_11096_));
 OA21x2_ASAP7_75t_R _30573_ (.A1(_11093_),
    .A2(_11095_),
    .B(_11096_),
    .Y(_11097_));
 TAPCELL_ASAP7_75t_R PHY_259 ();
 NAND2x2_ASAP7_75t_R _30575_ (.A(_10976_),
    .B(_11092_),
    .Y(_11099_));
 OR2x2_ASAP7_75t_R _30576_ (.A(_10973_),
    .B(_11099_),
    .Y(_11100_));
 NAND2x1_ASAP7_75t_R _30577_ (.A(_11097_),
    .B(_11100_),
    .Y(_11101_));
 OAI21x1_ASAP7_75t_R _30578_ (.A1(_11093_),
    .A2(_11095_),
    .B(_11096_),
    .Y(_11102_));
 TAPCELL_ASAP7_75t_R PHY_258 ();
 AND4x1_ASAP7_75t_R _30580_ (.A(_07504_),
    .B(_09351_),
    .C(_10973_),
    .D(_10976_),
    .Y(_11104_));
 OAI21x1_ASAP7_75t_R _30581_ (.A1(_11102_),
    .A2(_11104_),
    .B(_00660_),
    .Y(_11105_));
 OA21x2_ASAP7_75t_R _30582_ (.A1(_00660_),
    .A2(_11101_),
    .B(_11105_),
    .Y(_03919_));
 TAPCELL_ASAP7_75t_R PHY_257 ();
 AO21x2_ASAP7_75t_R _30584_ (.A1(_18114_),
    .A2(_07311_),
    .B(_09362_),
    .Y(_11107_));
 NAND3x2_ASAP7_75t_R _30585_ (.B(_09351_),
    .C(_10976_),
    .Y(_11108_),
    .A(_07170_));
 TAPCELL_ASAP7_75t_R PHY_256 ();
 AO32x1_ASAP7_75t_R _30587_ (.A1(_11107_),
    .A2(_10976_),
    .A3(_11092_),
    .B1(_11108_),
    .B2(_02392_),
    .Y(_11110_));
 NAND2x1_ASAP7_75t_R _30588_ (.A(_11097_),
    .B(_11110_),
    .Y(_11111_));
 OA21x2_ASAP7_75t_R _30589_ (.A1(\cs_registers_i.mhpmcounter[2][1] ),
    .A2(_11097_),
    .B(_11111_),
    .Y(_03920_));
 AND2x6_ASAP7_75t_R _30590_ (.A(_10976_),
    .B(_11092_),
    .Y(_11112_));
 TAPCELL_ASAP7_75t_R PHY_255 ();
 TAPCELL_ASAP7_75t_R PHY_254 ();
 NAND2x1_ASAP7_75t_R _30593_ (.A(_09390_),
    .B(_11112_),
    .Y(_11115_));
 OA211x2_ASAP7_75t_R _30594_ (.A1(_02394_),
    .A2(_11112_),
    .B(_11115_),
    .C(_11097_),
    .Y(_11116_));
 AOI21x1_ASAP7_75t_R _30595_ (.A1(_01486_),
    .A2(_11102_),
    .B(_11116_),
    .Y(_03921_));
 TAPCELL_ASAP7_75t_R PHY_253 ();
 TAPCELL_ASAP7_75t_R PHY_252 ();
 AO21x1_ASAP7_75t_R _30598_ (.A1(_02393_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11119_));
 TAPCELL_ASAP7_75t_R PHY_251 ();
 TAPCELL_ASAP7_75t_R PHY_250 ();
 TAPCELL_ASAP7_75t_R PHY_249 ();
 OR3x1_ASAP7_75t_R _30602_ (.A(_01485_),
    .B(_02393_),
    .C(_11112_),
    .Y(_11123_));
 OAI21x1_ASAP7_75t_R _30603_ (.A1(_09397_),
    .A2(_11099_),
    .B(_11123_),
    .Y(_11124_));
 AOI22x1_ASAP7_75t_R _30604_ (.A1(_01485_),
    .A2(_11119_),
    .B1(_11124_),
    .B2(_11097_),
    .Y(_03922_));
 NAND2x1_ASAP7_75t_R _30605_ (.A(_09408_),
    .B(_11112_),
    .Y(_11125_));
 OA211x2_ASAP7_75t_R _30606_ (.A1(_02396_),
    .A2(_11112_),
    .B(_11125_),
    .C(_11097_),
    .Y(_11126_));
 AOI21x1_ASAP7_75t_R _30607_ (.A1(_01484_),
    .A2(_11102_),
    .B(_11126_),
    .Y(_03923_));
 TAPCELL_ASAP7_75t_R PHY_248 ();
 OR3x1_ASAP7_75t_R _30609_ (.A(_01483_),
    .B(_02395_),
    .C(_11112_),
    .Y(_11128_));
 OAI21x1_ASAP7_75t_R _30610_ (.A1(_09417_),
    .A2(_11099_),
    .B(_11128_),
    .Y(_11129_));
 AO21x1_ASAP7_75t_R _30611_ (.A1(_02395_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11130_));
 AOI22x1_ASAP7_75t_R _30612_ (.A1(_11097_),
    .A2(_11129_),
    .B1(_11130_),
    .B2(_01483_),
    .Y(_03924_));
 TAPCELL_ASAP7_75t_R PHY_247 ();
 TAPCELL_ASAP7_75t_R PHY_246 ();
 NOR2x1_ASAP7_75t_R _30615_ (.A(_09426_),
    .B(_11099_),
    .Y(_11133_));
 AO21x1_ASAP7_75t_R _30616_ (.A1(_02398_),
    .A2(_11099_),
    .B(_11133_),
    .Y(_11134_));
 TAPCELL_ASAP7_75t_R PHY_245 ();
 AND2x2_ASAP7_75t_R _30618_ (.A(_01482_),
    .B(_11102_),
    .Y(_11136_));
 AOI21x1_ASAP7_75t_R _30619_ (.A1(_11097_),
    .A2(_11134_),
    .B(_11136_),
    .Y(_03925_));
 OR3x1_ASAP7_75t_R _30620_ (.A(_01481_),
    .B(_02397_),
    .C(_11112_),
    .Y(_11137_));
 OAI21x1_ASAP7_75t_R _30621_ (.A1(_09432_),
    .A2(_11099_),
    .B(_11137_),
    .Y(_11138_));
 AO21x1_ASAP7_75t_R _30622_ (.A1(_02397_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11139_));
 AOI22x1_ASAP7_75t_R _30623_ (.A1(_11097_),
    .A2(_11138_),
    .B1(_11139_),
    .B2(_01481_),
    .Y(_03926_));
 NOR2x1_ASAP7_75t_R _30624_ (.A(_09438_),
    .B(_11099_),
    .Y(_11140_));
 AO21x1_ASAP7_75t_R _30625_ (.A1(_02400_),
    .A2(_11099_),
    .B(_11140_),
    .Y(_11141_));
 AND2x2_ASAP7_75t_R _30626_ (.A(_01480_),
    .B(_11102_),
    .Y(_11142_));
 AOI21x1_ASAP7_75t_R _30627_ (.A1(_11097_),
    .A2(_11141_),
    .B(_11142_),
    .Y(_03927_));
 OR3x1_ASAP7_75t_R _30628_ (.A(_01479_),
    .B(_02399_),
    .C(_11112_),
    .Y(_11143_));
 OAI21x1_ASAP7_75t_R _30629_ (.A1(_09445_),
    .A2(_11099_),
    .B(_11143_),
    .Y(_11144_));
 AO21x1_ASAP7_75t_R _30630_ (.A1(_02399_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11145_));
 AOI22x1_ASAP7_75t_R _30631_ (.A1(_11097_),
    .A2(_11144_),
    .B1(_11145_),
    .B2(_01479_),
    .Y(_03928_));
 NOR2x1_ASAP7_75t_R _30632_ (.A(_09452_),
    .B(_11099_),
    .Y(_11146_));
 AO21x1_ASAP7_75t_R _30633_ (.A1(_02402_),
    .A2(_11099_),
    .B(_11146_),
    .Y(_11147_));
 AND2x2_ASAP7_75t_R _30634_ (.A(_01478_),
    .B(_11102_),
    .Y(_11148_));
 AOI21x1_ASAP7_75t_R _30635_ (.A1(_11097_),
    .A2(_11147_),
    .B(_11148_),
    .Y(_03929_));
 AO21x1_ASAP7_75t_R _30636_ (.A1(_02401_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11149_));
 OR3x1_ASAP7_75t_R _30637_ (.A(_01477_),
    .B(_02401_),
    .C(_11112_),
    .Y(_11150_));
 OAI21x1_ASAP7_75t_R _30638_ (.A1(_09458_),
    .A2(_11099_),
    .B(_11150_),
    .Y(_11151_));
 AOI22x1_ASAP7_75t_R _30639_ (.A1(_01477_),
    .A2(_11149_),
    .B1(_11151_),
    .B2(_11097_),
    .Y(_03930_));
 NOR2x1_ASAP7_75t_R _30640_ (.A(_09465_),
    .B(_11099_),
    .Y(_11152_));
 AO21x1_ASAP7_75t_R _30641_ (.A1(_02404_),
    .A2(_11099_),
    .B(_11152_),
    .Y(_11153_));
 AND2x2_ASAP7_75t_R _30642_ (.A(_01476_),
    .B(_11102_),
    .Y(_11154_));
 AOI21x1_ASAP7_75t_R _30643_ (.A1(_11097_),
    .A2(_11153_),
    .B(_11154_),
    .Y(_03931_));
 TAPCELL_ASAP7_75t_R PHY_244 ();
 AO21x1_ASAP7_75t_R _30645_ (.A1(_02403_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11156_));
 OR3x1_ASAP7_75t_R _30646_ (.A(_01475_),
    .B(_02403_),
    .C(_11112_),
    .Y(_11157_));
 OAI21x1_ASAP7_75t_R _30647_ (.A1(_09473_),
    .A2(_11099_),
    .B(_11157_),
    .Y(_11158_));
 AOI22x1_ASAP7_75t_R _30648_ (.A1(_01475_),
    .A2(_11156_),
    .B1(_11158_),
    .B2(_11097_),
    .Y(_03932_));
 NOR2x1_ASAP7_75t_R _30649_ (.A(_09481_),
    .B(_11099_),
    .Y(_11159_));
 AO21x1_ASAP7_75t_R _30650_ (.A1(_02406_),
    .A2(_11099_),
    .B(_11159_),
    .Y(_11160_));
 AND2x2_ASAP7_75t_R _30651_ (.A(_01474_),
    .B(_11102_),
    .Y(_11161_));
 AOI21x1_ASAP7_75t_R _30652_ (.A1(_11097_),
    .A2(_11160_),
    .B(_11161_),
    .Y(_03933_));
 AO21x1_ASAP7_75t_R _30653_ (.A1(_02405_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11162_));
 OR3x1_ASAP7_75t_R _30654_ (.A(_01473_),
    .B(_02405_),
    .C(_11112_),
    .Y(_11163_));
 OAI21x1_ASAP7_75t_R _30655_ (.A1(_09488_),
    .A2(_11099_),
    .B(_11163_),
    .Y(_11164_));
 AOI22x1_ASAP7_75t_R _30656_ (.A1(_01473_),
    .A2(_11162_),
    .B1(_11164_),
    .B2(_11097_),
    .Y(_03934_));
 NAND2x1_ASAP7_75t_R _30657_ (.A(_09496_),
    .B(_11112_),
    .Y(_11165_));
 OA211x2_ASAP7_75t_R _30658_ (.A1(_02408_),
    .A2(_11112_),
    .B(_11165_),
    .C(_11097_),
    .Y(_11166_));
 AOI21x1_ASAP7_75t_R _30659_ (.A1(_01472_),
    .A2(_11102_),
    .B(_11166_),
    .Y(_03935_));
 OR3x1_ASAP7_75t_R _30660_ (.A(_01471_),
    .B(_02407_),
    .C(_11112_),
    .Y(_11167_));
 OAI21x1_ASAP7_75t_R _30661_ (.A1(_09503_),
    .A2(_11099_),
    .B(_11167_),
    .Y(_11168_));
 AO21x1_ASAP7_75t_R _30662_ (.A1(_02407_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11169_));
 AOI22x1_ASAP7_75t_R _30663_ (.A1(_11097_),
    .A2(_11168_),
    .B1(_11169_),
    .B2(_01471_),
    .Y(_03936_));
 NAND2x1_ASAP7_75t_R _30664_ (.A(_09512_),
    .B(_11112_),
    .Y(_11170_));
 OA211x2_ASAP7_75t_R _30665_ (.A1(_02410_),
    .A2(_11112_),
    .B(_11170_),
    .C(_11097_),
    .Y(_11171_));
 AOI21x1_ASAP7_75t_R _30666_ (.A1(_01470_),
    .A2(_11102_),
    .B(_11171_),
    .Y(_03937_));
 INVx1_ASAP7_75t_R _30667_ (.A(_01469_),
    .Y(_11172_));
 AO21x1_ASAP7_75t_R _30668_ (.A1(_02409_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11173_));
 AND3x4_ASAP7_75t_R _30669_ (.A(_07170_),
    .B(_09351_),
    .C(_10976_),
    .Y(_11174_));
 TAPCELL_ASAP7_75t_R PHY_243 ();
 INVx1_ASAP7_75t_R _30671_ (.A(_02409_),
    .Y(_11176_));
 AND3x1_ASAP7_75t_R _30672_ (.A(_01469_),
    .B(_11176_),
    .C(_11108_),
    .Y(_11177_));
 AO21x1_ASAP7_75t_R _30673_ (.A1(_09519_),
    .A2(_11174_),
    .B(_11177_),
    .Y(_11178_));
 AO22x1_ASAP7_75t_R _30674_ (.A1(_11172_),
    .A2(_11173_),
    .B1(_11178_),
    .B2(_11097_),
    .Y(_03938_));
 NOR2x1_ASAP7_75t_R _30675_ (.A(_09526_),
    .B(_11099_),
    .Y(_11179_));
 AO21x1_ASAP7_75t_R _30676_ (.A1(_02412_),
    .A2(_11099_),
    .B(_11179_),
    .Y(_11180_));
 AND2x2_ASAP7_75t_R _30677_ (.A(_01468_),
    .B(_11102_),
    .Y(_11181_));
 AOI21x1_ASAP7_75t_R _30678_ (.A1(_11097_),
    .A2(_11180_),
    .B(_11181_),
    .Y(_03939_));
 INVx1_ASAP7_75t_R _30679_ (.A(_02411_),
    .Y(_11182_));
 AND3x1_ASAP7_75t_R _30680_ (.A(_01467_),
    .B(_11182_),
    .C(_11108_),
    .Y(_11183_));
 AO21x1_ASAP7_75t_R _30681_ (.A1(_09532_),
    .A2(_11174_),
    .B(_11183_),
    .Y(_11184_));
 AO21x1_ASAP7_75t_R _30682_ (.A1(_02411_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11185_));
 AO22x1_ASAP7_75t_R _30683_ (.A1(_11097_),
    .A2(_11184_),
    .B1(_11185_),
    .B2(_05985_),
    .Y(_03940_));
 NOR2x2_ASAP7_75t_R _30684_ (.A(_09539_),
    .B(_11099_),
    .Y(_11186_));
 AOI21x1_ASAP7_75t_R _30685_ (.A1(_02414_),
    .A2(_11099_),
    .B(_11186_),
    .Y(_11187_));
 NAND2x1_ASAP7_75t_R _30686_ (.A(_01466_),
    .B(_11102_),
    .Y(_11188_));
 OA21x2_ASAP7_75t_R _30687_ (.A1(_11102_),
    .A2(_11187_),
    .B(_11188_),
    .Y(_03941_));
 AO21x1_ASAP7_75t_R _30688_ (.A1(_02413_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11189_));
 OR3x1_ASAP7_75t_R _30689_ (.A(_01465_),
    .B(_02413_),
    .C(_11112_),
    .Y(_11190_));
 OAI21x1_ASAP7_75t_R _30690_ (.A1(_09545_),
    .A2(_11099_),
    .B(_11190_),
    .Y(_11191_));
 AOI22x1_ASAP7_75t_R _30691_ (.A1(_01465_),
    .A2(_11189_),
    .B1(_11191_),
    .B2(_11097_),
    .Y(_03942_));
 AOI21x1_ASAP7_75t_R _30692_ (.A1(net292),
    .A2(_09553_),
    .B(_09559_),
    .Y(_11192_));
 INVx1_ASAP7_75t_R _30693_ (.A(_02416_),
    .Y(_11193_));
 AO221x1_ASAP7_75t_R _30694_ (.A1(_11192_),
    .A2(_11174_),
    .B1(_11099_),
    .B2(_11193_),
    .C(_11102_),
    .Y(_11194_));
 OA21x2_ASAP7_75t_R _30695_ (.A1(\cs_registers_i.mhpmcounter[2][24] ),
    .A2(_11097_),
    .B(_11194_),
    .Y(_03943_));
 AO21x1_ASAP7_75t_R _30696_ (.A1(_02415_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11195_));
 OR3x1_ASAP7_75t_R _30697_ (.A(_01463_),
    .B(_02415_),
    .C(_11112_),
    .Y(_11196_));
 OAI21x1_ASAP7_75t_R _30698_ (.A1(_09565_),
    .A2(_11099_),
    .B(_11196_),
    .Y(_11197_));
 AOI22x1_ASAP7_75t_R _30699_ (.A1(_01463_),
    .A2(_11195_),
    .B1(_11197_),
    .B2(_11097_),
    .Y(_03944_));
 NOR2x1_ASAP7_75t_R _30700_ (.A(_09572_),
    .B(_11099_),
    .Y(_11198_));
 AO21x1_ASAP7_75t_R _30701_ (.A1(_02418_),
    .A2(_11099_),
    .B(_11198_),
    .Y(_11199_));
 AND2x2_ASAP7_75t_R _30702_ (.A(_01462_),
    .B(_11102_),
    .Y(_11200_));
 AOI21x1_ASAP7_75t_R _30703_ (.A1(_11097_),
    .A2(_11199_),
    .B(_11200_),
    .Y(_03945_));
 INVx1_ASAP7_75t_R _30704_ (.A(_01461_),
    .Y(_11201_));
 AO21x1_ASAP7_75t_R _30705_ (.A1(_02417_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11202_));
 INVx2_ASAP7_75t_R _30706_ (.A(_09578_),
    .Y(_11203_));
 OR3x1_ASAP7_75t_R _30707_ (.A(_11201_),
    .B(_02417_),
    .C(_11174_),
    .Y(_11204_));
 OAI21x1_ASAP7_75t_R _30708_ (.A1(_11203_),
    .A2(_11108_),
    .B(_11204_),
    .Y(_11205_));
 AO22x1_ASAP7_75t_R _30709_ (.A1(_11201_),
    .A2(_11202_),
    .B1(_11205_),
    .B2(_11097_),
    .Y(_03946_));
 NAND2x1_ASAP7_75t_R _30710_ (.A(_09585_),
    .B(_11112_),
    .Y(_11206_));
 OAI21x1_ASAP7_75t_R _30711_ (.A1(_02420_),
    .A2(_11112_),
    .B(_11206_),
    .Y(_11207_));
 NAND2x1_ASAP7_75t_R _30712_ (.A(_01460_),
    .B(_11102_),
    .Y(_11208_));
 OA21x2_ASAP7_75t_R _30713_ (.A1(_11102_),
    .A2(_11207_),
    .B(_11208_),
    .Y(_03947_));
 INVx2_ASAP7_75t_R _30714_ (.A(_09591_),
    .Y(_11209_));
 OR3x1_ASAP7_75t_R _30715_ (.A(_05989_),
    .B(_02419_),
    .C(_11174_),
    .Y(_11210_));
 OAI21x1_ASAP7_75t_R _30716_ (.A1(_11209_),
    .A2(_11108_),
    .B(_11210_),
    .Y(_11211_));
 AO21x1_ASAP7_75t_R _30717_ (.A1(_02419_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11212_));
 AO22x1_ASAP7_75t_R _30718_ (.A1(_11097_),
    .A2(_11211_),
    .B1(_11212_),
    .B2(_05989_),
    .Y(_03948_));
 NAND2x1_ASAP7_75t_R _30719_ (.A(_09598_),
    .B(_11112_),
    .Y(_11213_));
 OA211x2_ASAP7_75t_R _30720_ (.A1(_02422_),
    .A2(_11112_),
    .B(_11213_),
    .C(_11097_),
    .Y(_11214_));
 AOI21x1_ASAP7_75t_R _30721_ (.A1(_01458_),
    .A2(_11102_),
    .B(_11214_),
    .Y(_03949_));
 INVx2_ASAP7_75t_R _30722_ (.A(_09605_),
    .Y(_11215_));
 INVx1_ASAP7_75t_R _30723_ (.A(_01457_),
    .Y(_11216_));
 OR3x1_ASAP7_75t_R _30724_ (.A(_11216_),
    .B(_02421_),
    .C(_11174_),
    .Y(_11217_));
 OAI21x1_ASAP7_75t_R _30725_ (.A1(_11215_),
    .A2(_11108_),
    .B(_11217_),
    .Y(_11218_));
 AO21x1_ASAP7_75t_R _30726_ (.A1(_02421_),
    .A2(_11108_),
    .B(_11102_),
    .Y(_11219_));
 AO22x1_ASAP7_75t_R _30727_ (.A1(_11097_),
    .A2(_11218_),
    .B1(_11219_),
    .B2(_11216_),
    .Y(_03950_));
 INVx1_ASAP7_75t_R _30728_ (.A(_07667_),
    .Y(_11220_));
 NAND2x2_ASAP7_75t_R _30729_ (.A(_11220_),
    .B(_09365_),
    .Y(_11221_));
 OR3x1_ASAP7_75t_R _30730_ (.A(_09458_),
    .B(_09465_),
    .C(_11221_),
    .Y(_11222_));
 OR3x1_ASAP7_75t_R _30731_ (.A(_06171_),
    .B(_06173_),
    .C(_06176_),
    .Y(_11223_));
 AO221x2_ASAP7_75t_R _30732_ (.A1(_11223_),
    .A2(_06340_),
    .B1(_06872_),
    .B2(_06327_),
    .C(_06251_),
    .Y(_11224_));
 INVx1_ASAP7_75t_R _30733_ (.A(_11224_),
    .Y(_11225_));
 OR3x4_ASAP7_75t_R _30734_ (.A(_05677_),
    .B(_06880_),
    .C(_11225_),
    .Y(_11226_));
 TAPCELL_ASAP7_75t_R PHY_242 ();
 NAND2x2_ASAP7_75t_R _30736_ (.A(_06262_),
    .B(_11226_),
    .Y(_11228_));
 AOI21x1_ASAP7_75t_R _30737_ (.A1(_01456_),
    .A2(_11221_),
    .B(_11228_),
    .Y(_11229_));
 TAPCELL_ASAP7_75t_R PHY_241 ();
 OR3x4_ASAP7_75t_R _30739_ (.A(_01718_),
    .B(_05712_),
    .C(_06257_),
    .Y(_11231_));
 TAPCELL_ASAP7_75t_R PHY_240 ();
 OAI22x1_ASAP7_75t_R _30741_ (.A1(_02140_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_02107_),
    .Y(_11233_));
 AO21x1_ASAP7_75t_R _30742_ (.A1(_11222_),
    .A2(_11229_),
    .B(_11233_),
    .Y(_03951_));
 AOI21x1_ASAP7_75t_R _30743_ (.A1(_01455_),
    .A2(_11221_),
    .B(_11228_),
    .Y(_11234_));
 OAI22x1_ASAP7_75t_R _30744_ (.A1(_17592_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_02106_),
    .Y(_11235_));
 AO21x1_ASAP7_75t_R _30745_ (.A1(_11222_),
    .A2(_11234_),
    .B(_11235_),
    .Y(_03952_));
 INVx2_ASAP7_75t_R _30746_ (.A(_09432_),
    .Y(_11236_));
 AND3x4_ASAP7_75t_R _30747_ (.A(_05632_),
    .B(_09364_),
    .C(_09351_),
    .Y(_11237_));
 TAPCELL_ASAP7_75t_R PHY_239 ();
 NAND2x2_ASAP7_75t_R _30749_ (.A(_05582_),
    .B(_11237_),
    .Y(_11239_));
 AO21x1_ASAP7_75t_R _30750_ (.A1(_06828_),
    .A2(_02105_),
    .B(_06262_),
    .Y(_11240_));
 INVx1_ASAP7_75t_R _30751_ (.A(_11221_),
    .Y(_11241_));
 AND3x4_ASAP7_75t_R _30752_ (.A(_01311_),
    .B(_06873_),
    .C(_11224_),
    .Y(_11242_));
 NOR2x2_ASAP7_75t_R _30753_ (.A(_01718_),
    .B(_06262_),
    .Y(_11243_));
 OR2x6_ASAP7_75t_R _30754_ (.A(_11242_),
    .B(_11243_),
    .Y(_11244_));
 TAPCELL_ASAP7_75t_R PHY_238 ();
 OA21x2_ASAP7_75t_R _30756_ (.A1(_02105_),
    .A2(_11224_),
    .B(_11244_),
    .Y(_11246_));
 OR3x1_ASAP7_75t_R _30757_ (.A(_01454_),
    .B(_11241_),
    .C(_11246_),
    .Y(_11247_));
 OA211x2_ASAP7_75t_R _30758_ (.A1(_01453_),
    .A2(_11226_),
    .B(_11240_),
    .C(_11247_),
    .Y(_11248_));
 OAI21x1_ASAP7_75t_R _30759_ (.A1(_11236_),
    .A2(_11239_),
    .B(_11248_),
    .Y(_03953_));
 NOR2x1_ASAP7_75t_R _30760_ (.A(_09397_),
    .B(_11239_),
    .Y(_11249_));
 AO21x1_ASAP7_75t_R _30761_ (.A1(_01453_),
    .A2(_11239_),
    .B(_11249_),
    .Y(_11250_));
 OAI22x1_ASAP7_75t_R _30762_ (.A1(_01454_),
    .A2(_06262_),
    .B1(_11228_),
    .B2(_11250_),
    .Y(_03954_));
 INVx1_ASAP7_75t_R _30763_ (.A(_01452_),
    .Y(_11251_));
 OR2x6_ASAP7_75t_R _30764_ (.A(_01873_),
    .B(_05747_),
    .Y(_11252_));
 TAPCELL_ASAP7_75t_R PHY_237 ();
 TAPCELL_ASAP7_75t_R PHY_236 ();
 AO21x1_ASAP7_75t_R _30767_ (.A1(_05420_),
    .A2(_05909_),
    .B(_13640_),
    .Y(_11255_));
 OA211x2_ASAP7_75t_R _30768_ (.A1(net280),
    .A2(_08581_),
    .B(_11255_),
    .C(_05755_),
    .Y(_11256_));
 AO21x1_ASAP7_75t_R _30769_ (.A1(_11251_),
    .A2(_11252_),
    .B(_11256_),
    .Y(_03955_));
 TAPCELL_ASAP7_75t_R PHY_235 ();
 TAPCELL_ASAP7_75t_R PHY_234 ();
 AOI22x1_ASAP7_75t_R _30772_ (.A1(_13217_),
    .A2(_05910_),
    .B1(_08580_),
    .B2(_16499_),
    .Y(_11259_));
 TAPCELL_ASAP7_75t_R PHY_233 ();
 NOR2x1_ASAP7_75t_R _30774_ (.A(_01451_),
    .B(_05755_),
    .Y(_11261_));
 AO21x1_ASAP7_75t_R _30775_ (.A1(_05755_),
    .A2(_11259_),
    .B(_11261_),
    .Y(_03956_));
 TAPCELL_ASAP7_75t_R PHY_232 ();
 AO21x1_ASAP7_75t_R _30777_ (.A1(_05420_),
    .A2(_05909_),
    .B(_06098_),
    .Y(_11263_));
 OA211x2_ASAP7_75t_R _30778_ (.A1(_05767_),
    .A2(_05910_),
    .B(_11263_),
    .C(_05755_),
    .Y(_11264_));
 AOI21x1_ASAP7_75t_R _30779_ (.A1(_01450_),
    .A2(_11252_),
    .B(_11264_),
    .Y(_03957_));
 TAPCELL_ASAP7_75t_R PHY_231 ();
 OR2x2_ASAP7_75t_R _30781_ (.A(_06102_),
    .B(_08580_),
    .Y(_11266_));
 OA211x2_ASAP7_75t_R _30782_ (.A1(_06277_),
    .A2(_08581_),
    .B(_11266_),
    .C(_05755_),
    .Y(_11267_));
 AOI21x1_ASAP7_75t_R _30783_ (.A1(_01449_),
    .A2(_11252_),
    .B(_11267_),
    .Y(_03958_));
 NAND2x1_ASAP7_75t_R _30784_ (.A(_14080_),
    .B(_05910_),
    .Y(_11268_));
 OA211x2_ASAP7_75t_R _30785_ (.A1(_05766_),
    .A2(_05910_),
    .B(_11268_),
    .C(_05755_),
    .Y(_11269_));
 AOI21x1_ASAP7_75t_R _30786_ (.A1(_01448_),
    .A2(_11252_),
    .B(_11269_),
    .Y(_03959_));
 AO221x1_ASAP7_75t_R _30787_ (.A1(_06108_),
    .A2(_05910_),
    .B1(_08580_),
    .B2(_08767_),
    .C(_11252_),
    .Y(_11270_));
 OAI21x1_ASAP7_75t_R _30788_ (.A1(_01447_),
    .A2(_05755_),
    .B(_11270_),
    .Y(_03960_));
 AO21x1_ASAP7_75t_R _30789_ (.A1(_05420_),
    .A2(_05909_),
    .B(_05605_),
    .Y(_11271_));
 OA211x2_ASAP7_75t_R _30790_ (.A1(_05768_),
    .A2(_05910_),
    .B(_11271_),
    .C(_05755_),
    .Y(_11272_));
 AOI21x1_ASAP7_75t_R _30791_ (.A1(_01446_),
    .A2(_11252_),
    .B(_11272_),
    .Y(_03961_));
 AO221x1_ASAP7_75t_R _30792_ (.A1(_05653_),
    .A2(_05910_),
    .B1(_08580_),
    .B2(_00676_),
    .C(_11252_),
    .Y(_11273_));
 OAI21x1_ASAP7_75t_R _30793_ (.A1(_01445_),
    .A2(_05755_),
    .B(_11273_),
    .Y(_03962_));
 AO221x1_ASAP7_75t_R _30794_ (.A1(_06060_),
    .A2(_05910_),
    .B1(_08580_),
    .B2(_05773_),
    .C(_11252_),
    .Y(_11274_));
 OAI21x1_ASAP7_75t_R _30795_ (.A1(_01444_),
    .A2(_05755_),
    .B(_11274_),
    .Y(_03963_));
 INVx1_ASAP7_75t_R _30796_ (.A(_14373_),
    .Y(_11275_));
 AO221x1_ASAP7_75t_R _30797_ (.A1(_11275_),
    .A2(_05910_),
    .B1(_08580_),
    .B2(_06350_),
    .C(_11252_),
    .Y(_11276_));
 OAI21x1_ASAP7_75t_R _30798_ (.A1(_01443_),
    .A2(_05755_),
    .B(_11276_),
    .Y(_03964_));
 AO21x1_ASAP7_75t_R _30799_ (.A1(_05420_),
    .A2(_05909_),
    .B(_05672_),
    .Y(_11277_));
 OA211x2_ASAP7_75t_R _30800_ (.A1(_05772_),
    .A2(_05910_),
    .B(_11277_),
    .C(_05755_),
    .Y(_11278_));
 AOI21x1_ASAP7_75t_R _30801_ (.A1(_01442_),
    .A2(_11252_),
    .B(_11278_),
    .Y(_03965_));
 AO221x1_ASAP7_75t_R _30802_ (.A1(_15160_),
    .A2(_05910_),
    .B1(_08580_),
    .B2(_06368_),
    .C(_11252_),
    .Y(_11279_));
 OAI21x1_ASAP7_75t_R _30803_ (.A1(_01441_),
    .A2(_05755_),
    .B(_11279_),
    .Y(_03966_));
 TAPCELL_ASAP7_75t_R PHY_230 ();
 OR2x2_ASAP7_75t_R _30805_ (.A(_15266_),
    .B(_08580_),
    .Y(_11281_));
 OA211x2_ASAP7_75t_R _30806_ (.A1(_05771_),
    .A2(_08581_),
    .B(_11281_),
    .C(_05755_),
    .Y(_11282_));
 AOI21x1_ASAP7_75t_R _30807_ (.A1(_02221_),
    .A2(_11252_),
    .B(_11282_),
    .Y(_03967_));
 OR2x2_ASAP7_75t_R _30808_ (.A(_15352_),
    .B(_08580_),
    .Y(_11283_));
 OA211x2_ASAP7_75t_R _30809_ (.A1(_06384_),
    .A2(_08581_),
    .B(_11283_),
    .C(_05755_),
    .Y(_11284_));
 AOI21x1_ASAP7_75t_R _30810_ (.A1(_02220_),
    .A2(_11252_),
    .B(_11284_),
    .Y(_03968_));
 INVx1_ASAP7_75t_R _30811_ (.A(_02219_),
    .Y(_11285_));
 AO221x1_ASAP7_75t_R _30812_ (.A1(_05887_),
    .A2(_05910_),
    .B1(_08580_),
    .B2(net155),
    .C(_11252_),
    .Y(_11286_));
 OA21x2_ASAP7_75t_R _30813_ (.A1(_11285_),
    .A2(_05755_),
    .B(_11286_),
    .Y(_03969_));
 NAND2x1_ASAP7_75t_R _30814_ (.A(_15617_),
    .B(_08581_),
    .Y(_11287_));
 OA211x2_ASAP7_75t_R _30815_ (.A1(_00785_),
    .A2(_08581_),
    .B(_11287_),
    .C(_05755_),
    .Y(_11288_));
 AOI21x1_ASAP7_75t_R _30816_ (.A1(_02218_),
    .A2(_11252_),
    .B(_11288_),
    .Y(_03970_));
 OR2x2_ASAP7_75t_R _30817_ (.A(_15731_),
    .B(_08580_),
    .Y(_11289_));
 OA211x2_ASAP7_75t_R _30818_ (.A1(_05770_),
    .A2(_08581_),
    .B(_11289_),
    .C(_05755_),
    .Y(_11290_));
 AOI21x1_ASAP7_75t_R _30819_ (.A1(_02217_),
    .A2(_11252_),
    .B(_11290_),
    .Y(_03971_));
 NAND2x1_ASAP7_75t_R _30820_ (.A(_15841_),
    .B(_08581_),
    .Y(_11291_));
 TAPCELL_ASAP7_75t_R PHY_229 ();
 OA211x2_ASAP7_75t_R _30822_ (.A1(_06412_),
    .A2(_08581_),
    .B(_11291_),
    .C(_05755_),
    .Y(_11293_));
 AOI21x1_ASAP7_75t_R _30823_ (.A1(_02216_),
    .A2(_11252_),
    .B(_11293_),
    .Y(_03972_));
 TAPCELL_ASAP7_75t_R PHY_228 ();
 OR2x2_ASAP7_75t_R _30825_ (.A(_15971_),
    .B(_08580_),
    .Y(_11295_));
 OA211x2_ASAP7_75t_R _30826_ (.A1(_16020_),
    .A2(_08581_),
    .B(_11295_),
    .C(_05755_),
    .Y(_11296_));
 AOI21x1_ASAP7_75t_R _30827_ (.A1(_02215_),
    .A2(_11252_),
    .B(_11296_),
    .Y(_03973_));
 INVx1_ASAP7_75t_R _30828_ (.A(_16083_),
    .Y(_11297_));
 AO221x1_ASAP7_75t_R _30829_ (.A1(_11297_),
    .A2(_05910_),
    .B1(_08580_),
    .B2(net257),
    .C(_11252_),
    .Y(_11298_));
 OA21x2_ASAP7_75t_R _30830_ (.A1(_16088_),
    .A2(_05755_),
    .B(_11298_),
    .Y(_03974_));
 NAND2x1_ASAP7_75t_R _30831_ (.A(_16204_),
    .B(_08581_),
    .Y(_11299_));
 OA211x2_ASAP7_75t_R _30832_ (.A1(_16260_),
    .A2(_08581_),
    .B(_11299_),
    .C(_05755_),
    .Y(_11300_));
 AOI21x1_ASAP7_75t_R _30833_ (.A1(_02213_),
    .A2(_11252_),
    .B(_11300_),
    .Y(_03975_));
 OR2x2_ASAP7_75t_R _30834_ (.A(_16324_),
    .B(_08580_),
    .Y(_11301_));
 OA211x2_ASAP7_75t_R _30835_ (.A1(_06440_),
    .A2(_08581_),
    .B(_11301_),
    .C(_05755_),
    .Y(_11302_));
 AOI21x1_ASAP7_75t_R _30836_ (.A1(_02212_),
    .A2(_11252_),
    .B(_11302_),
    .Y(_03976_));
 OR2x2_ASAP7_75t_R _30837_ (.A(_16433_),
    .B(_08580_),
    .Y(_11303_));
 OA211x2_ASAP7_75t_R _30838_ (.A1(_05760_),
    .A2(_08581_),
    .B(_11303_),
    .C(_05755_),
    .Y(_11304_));
 AOI21x1_ASAP7_75t_R _30839_ (.A1(_02211_),
    .A2(_11252_),
    .B(_11304_),
    .Y(_03977_));
 NAND2x1_ASAP7_75t_R _30840_ (.A(_04547_),
    .B(_08581_),
    .Y(_11305_));
 OA211x2_ASAP7_75t_R _30841_ (.A1(_06452_),
    .A2(_08581_),
    .B(_11305_),
    .C(_05755_),
    .Y(_11306_));
 AOI21x1_ASAP7_75t_R _30842_ (.A1(_02210_),
    .A2(_11252_),
    .B(_11306_),
    .Y(_03978_));
 INVx1_ASAP7_75t_R _30843_ (.A(_02209_),
    .Y(_11307_));
 AO221x1_ASAP7_75t_R _30844_ (.A1(_04667_),
    .A2(_05910_),
    .B1(_08580_),
    .B2(net165),
    .C(_11252_),
    .Y(_11308_));
 OA21x2_ASAP7_75t_R _30845_ (.A1(_11307_),
    .A2(_05755_),
    .B(_11308_),
    .Y(_03979_));
 OR2x2_ASAP7_75t_R _30846_ (.A(_04780_),
    .B(_08580_),
    .Y(_11309_));
 OA211x2_ASAP7_75t_R _30847_ (.A1(_06464_),
    .A2(_08581_),
    .B(_11309_),
    .C(_05755_),
    .Y(_11310_));
 AOI21x1_ASAP7_75t_R _30848_ (.A1(_02208_),
    .A2(_11252_),
    .B(_11310_),
    .Y(_03980_));
 OR2x2_ASAP7_75t_R _30849_ (.A(_04888_),
    .B(_08580_),
    .Y(_11311_));
 OA211x2_ASAP7_75t_R _30850_ (.A1(_04937_),
    .A2(_08581_),
    .B(_11311_),
    .C(_05755_),
    .Y(_11312_));
 AOI21x1_ASAP7_75t_R _30851_ (.A1(_02207_),
    .A2(_11252_),
    .B(_11312_),
    .Y(_03981_));
 OR2x2_ASAP7_75t_R _30852_ (.A(_04996_),
    .B(_08580_),
    .Y(_11313_));
 OA211x2_ASAP7_75t_R _30853_ (.A1(_06477_),
    .A2(_08581_),
    .B(_11313_),
    .C(_05755_),
    .Y(_11314_));
 AOI21x1_ASAP7_75t_R _30854_ (.A1(_02206_),
    .A2(_11252_),
    .B(_11314_),
    .Y(_03982_));
 OR2x2_ASAP7_75t_R _30855_ (.A(_05105_),
    .B(_08580_),
    .Y(_11315_));
 OA211x2_ASAP7_75t_R _30856_ (.A1(_05154_),
    .A2(_08581_),
    .B(_11315_),
    .C(_05755_),
    .Y(_11316_));
 AOI21x1_ASAP7_75t_R _30857_ (.A1(_02205_),
    .A2(_11252_),
    .B(_11316_),
    .Y(_03983_));
 OR2x2_ASAP7_75t_R _30858_ (.A(_05213_),
    .B(_08580_),
    .Y(_11317_));
 OA211x2_ASAP7_75t_R _30859_ (.A1(_06491_),
    .A2(_08581_),
    .B(_11317_),
    .C(_05755_),
    .Y(_11318_));
 AOI21x1_ASAP7_75t_R _30860_ (.A1(_02204_),
    .A2(_11252_),
    .B(_11318_),
    .Y(_03984_));
 OR2x2_ASAP7_75t_R _30861_ (.A(_05323_),
    .B(_08580_),
    .Y(_11319_));
 OA211x2_ASAP7_75t_R _30862_ (.A1(_05372_),
    .A2(_08581_),
    .B(_11319_),
    .C(_05755_),
    .Y(_11320_));
 AOI21x1_ASAP7_75t_R _30863_ (.A1(_02203_),
    .A2(_11252_),
    .B(_11320_),
    .Y(_03985_));
 AOI211x1_ASAP7_75t_R _30864_ (.A1(_05512_),
    .A2(_05909_),
    .B(_11252_),
    .C(_05484_),
    .Y(_11321_));
 AO21x1_ASAP7_75t_R _30865_ (.A1(_08606_),
    .A2(_11252_),
    .B(_11321_),
    .Y(_03986_));
 OR3x4_ASAP7_75t_R _30866_ (.A(_06312_),
    .B(net95),
    .C(_06516_),
    .Y(_11322_));
 TAPCELL_ASAP7_75t_R PHY_227 ();
 TAPCELL_ASAP7_75t_R PHY_226 ();
 TAPCELL_ASAP7_75t_R PHY_225 ();
 NAND2x1_ASAP7_75t_R _30870_ (.A(_02201_),
    .B(_11322_),
    .Y(_11326_));
 OA21x2_ASAP7_75t_R _30871_ (.A1(net239),
    .A2(_11322_),
    .B(_11326_),
    .Y(_03987_));
 NAND2x1_ASAP7_75t_R _30872_ (.A(_02200_),
    .B(_11322_),
    .Y(_11327_));
 OA21x2_ASAP7_75t_R _30873_ (.A1(net242),
    .A2(_11322_),
    .B(_11327_),
    .Y(_03988_));
 NAND2x1_ASAP7_75t_R _30874_ (.A(_02199_),
    .B(_11322_),
    .Y(_11328_));
 OA21x2_ASAP7_75t_R _30875_ (.A1(net243),
    .A2(_11322_),
    .B(_11328_),
    .Y(_03989_));
 NAND2x1_ASAP7_75t_R _30876_ (.A(_02198_),
    .B(_11322_),
    .Y(_11329_));
 OA21x2_ASAP7_75t_R _30877_ (.A1(net244),
    .A2(_11322_),
    .B(_11329_),
    .Y(_03990_));
 NAND2x1_ASAP7_75t_R _30878_ (.A(_02197_),
    .B(_11322_),
    .Y(_11330_));
 OA21x2_ASAP7_75t_R _30879_ (.A1(net245),
    .A2(_11322_),
    .B(_11330_),
    .Y(_03991_));
 NAND2x1_ASAP7_75t_R _30880_ (.A(_02196_),
    .B(_11322_),
    .Y(_11331_));
 OA21x2_ASAP7_75t_R _30881_ (.A1(net246),
    .A2(_11322_),
    .B(_11331_),
    .Y(_03992_));
 NOR2x1_ASAP7_75t_R _30882_ (.A(net247),
    .B(_11322_),
    .Y(_11332_));
 AOI21x1_ASAP7_75t_R _30883_ (.A1(_02195_),
    .A2(_11322_),
    .B(_11332_),
    .Y(_03993_));
 NAND2x1_ASAP7_75t_R _30884_ (.A(_02194_),
    .B(_11322_),
    .Y(_11333_));
 OA21x2_ASAP7_75t_R _30885_ (.A1(net248),
    .A2(_11322_),
    .B(_11333_),
    .Y(_03994_));
 NAND2x1_ASAP7_75t_R _30886_ (.A(_02193_),
    .B(_11322_),
    .Y(_11334_));
 OA21x2_ASAP7_75t_R _30887_ (.A1(net219),
    .A2(_11322_),
    .B(_11334_),
    .Y(_03995_));
 NAND2x1_ASAP7_75t_R _30888_ (.A(_02192_),
    .B(_11322_),
    .Y(_11335_));
 OA21x2_ASAP7_75t_R _30889_ (.A1(net220),
    .A2(_11322_),
    .B(_11335_),
    .Y(_03996_));
 TAPCELL_ASAP7_75t_R PHY_224 ();
 TAPCELL_ASAP7_75t_R PHY_223 ();
 NAND2x1_ASAP7_75t_R _30892_ (.A(_02191_),
    .B(_11322_),
    .Y(_11338_));
 OA21x2_ASAP7_75t_R _30893_ (.A1(net221),
    .A2(_11322_),
    .B(_11338_),
    .Y(_03997_));
 NAND2x1_ASAP7_75t_R _30894_ (.A(_02190_),
    .B(_11322_),
    .Y(_11339_));
 OA21x2_ASAP7_75t_R _30895_ (.A1(net222),
    .A2(_11322_),
    .B(_11339_),
    .Y(_03998_));
 NAND2x1_ASAP7_75t_R _30896_ (.A(_02189_),
    .B(_11322_),
    .Y(_11340_));
 OA21x2_ASAP7_75t_R _30897_ (.A1(net223),
    .A2(_11322_),
    .B(_11340_),
    .Y(_03999_));
 NAND2x1_ASAP7_75t_R _30898_ (.A(_02188_),
    .B(_11322_),
    .Y(_11341_));
 OA21x2_ASAP7_75t_R _30899_ (.A1(net224),
    .A2(_11322_),
    .B(_11341_),
    .Y(_04000_));
 NAND2x1_ASAP7_75t_R _30900_ (.A(_02187_),
    .B(_11322_),
    .Y(_11342_));
 OA21x2_ASAP7_75t_R _30901_ (.A1(net225),
    .A2(_11322_),
    .B(_11342_),
    .Y(_04001_));
 NAND2x1_ASAP7_75t_R _30902_ (.A(_02186_),
    .B(_11322_),
    .Y(_11343_));
 OA21x2_ASAP7_75t_R _30903_ (.A1(net226),
    .A2(_11322_),
    .B(_11343_),
    .Y(_04002_));
 NAND2x1_ASAP7_75t_R _30904_ (.A(_02185_),
    .B(_11322_),
    .Y(_11344_));
 OA21x2_ASAP7_75t_R _30905_ (.A1(net227),
    .A2(_11322_),
    .B(_11344_),
    .Y(_04003_));
 NAND2x1_ASAP7_75t_R _30906_ (.A(_02184_),
    .B(_11322_),
    .Y(_11345_));
 OA21x2_ASAP7_75t_R _30907_ (.A1(net228),
    .A2(_11322_),
    .B(_11345_),
    .Y(_04004_));
 NAND2x1_ASAP7_75t_R _30908_ (.A(_02183_),
    .B(_11322_),
    .Y(_11346_));
 OA21x2_ASAP7_75t_R _30909_ (.A1(net229),
    .A2(_11322_),
    .B(_11346_),
    .Y(_04005_));
 NAND2x1_ASAP7_75t_R _30910_ (.A(_02182_),
    .B(_11322_),
    .Y(_11347_));
 OA21x2_ASAP7_75t_R _30911_ (.A1(net230),
    .A2(_11322_),
    .B(_11347_),
    .Y(_04006_));
 TAPCELL_ASAP7_75t_R PHY_222 ();
 TAPCELL_ASAP7_75t_R PHY_221 ();
 NAND2x1_ASAP7_75t_R _30914_ (.A(_02181_),
    .B(_11322_),
    .Y(_11350_));
 OA21x2_ASAP7_75t_R _30915_ (.A1(net231),
    .A2(_11322_),
    .B(_11350_),
    .Y(_04007_));
 NAND2x1_ASAP7_75t_R _30916_ (.A(_02180_),
    .B(_11322_),
    .Y(_11351_));
 OA21x2_ASAP7_75t_R _30917_ (.A1(net232),
    .A2(_11322_),
    .B(_11351_),
    .Y(_04008_));
 NAND2x1_ASAP7_75t_R _30918_ (.A(_02179_),
    .B(_11322_),
    .Y(_11352_));
 OA21x2_ASAP7_75t_R _30919_ (.A1(net233),
    .A2(_11322_),
    .B(_11352_),
    .Y(_04009_));
 NAND2x1_ASAP7_75t_R _30920_ (.A(_02178_),
    .B(_11322_),
    .Y(_11353_));
 OA21x2_ASAP7_75t_R _30921_ (.A1(net234),
    .A2(_11322_),
    .B(_11353_),
    .Y(_04010_));
 NAND2x1_ASAP7_75t_R _30922_ (.A(_02177_),
    .B(_11322_),
    .Y(_11354_));
 OA21x2_ASAP7_75t_R _30923_ (.A1(net235),
    .A2(_11322_),
    .B(_11354_),
    .Y(_04011_));
 NAND2x1_ASAP7_75t_R _30924_ (.A(_02176_),
    .B(_11322_),
    .Y(_11355_));
 OA21x2_ASAP7_75t_R _30925_ (.A1(net236),
    .A2(_11322_),
    .B(_11355_),
    .Y(_04012_));
 NAND2x1_ASAP7_75t_R _30926_ (.A(_02175_),
    .B(_11322_),
    .Y(_11356_));
 OA21x2_ASAP7_75t_R _30927_ (.A1(net237),
    .A2(_11322_),
    .B(_11356_),
    .Y(_04013_));
 NAND2x1_ASAP7_75t_R _30928_ (.A(_02174_),
    .B(_11322_),
    .Y(_11357_));
 OA21x2_ASAP7_75t_R _30929_ (.A1(net238),
    .A2(_11322_),
    .B(_11357_),
    .Y(_04014_));
 NAND2x1_ASAP7_75t_R _30930_ (.A(_02173_),
    .B(_11322_),
    .Y(_11358_));
 OA21x2_ASAP7_75t_R _30931_ (.A1(net240),
    .A2(_11322_),
    .B(_11358_),
    .Y(_04015_));
 NAND2x1_ASAP7_75t_R _30932_ (.A(_01729_),
    .B(_11322_),
    .Y(_11359_));
 OA21x2_ASAP7_75t_R _30933_ (.A1(net241),
    .A2(_11322_),
    .B(_11359_),
    .Y(_04016_));
 AOI22x1_ASAP7_75t_R _30934_ (.A1(_10975_),
    .A2(_10982_),
    .B1(_10983_),
    .B2(_00661_),
    .Y(_11360_));
 TAPCELL_ASAP7_75t_R PHY_220 ();
 OR2x2_ASAP7_75t_R _30936_ (.A(_10983_),
    .B(_10973_),
    .Y(_11362_));
 AO22x2_ASAP7_75t_R _30937_ (.A1(_10975_),
    .A2(_10982_),
    .B1(_10983_),
    .B2(_00661_),
    .Y(_11363_));
 TAPCELL_ASAP7_75t_R PHY_219 ();
 OA211x2_ASAP7_75t_R _30939_ (.A1(_02488_),
    .A2(_10978_),
    .B(_11362_),
    .C(_11363_),
    .Y(_11365_));
 AOI21x1_ASAP7_75t_R _30940_ (.A1(_02172_),
    .A2(_11360_),
    .B(_11365_),
    .Y(_04017_));
 TAPCELL_ASAP7_75t_R PHY_218 ();
 OR3x1_ASAP7_75t_R _30942_ (.A(_02171_),
    .B(_02487_),
    .C(_10978_),
    .Y(_11367_));
 OAI21x1_ASAP7_75t_R _30943_ (.A1(_09363_),
    .A2(_10986_),
    .B(_11367_),
    .Y(_11368_));
 TAPCELL_ASAP7_75t_R PHY_217 ();
 AO21x1_ASAP7_75t_R _30945_ (.A1(_02487_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11370_));
 AOI22x1_ASAP7_75t_R _30946_ (.A1(_11363_),
    .A2(_11368_),
    .B1(_11370_),
    .B2(_02171_),
    .Y(_04018_));
 OA211x2_ASAP7_75t_R _30947_ (.A1(_02490_),
    .A2(_10978_),
    .B(_10995_),
    .C(_11363_),
    .Y(_11371_));
 AOI21x1_ASAP7_75t_R _30948_ (.A1(_02170_),
    .A2(_11360_),
    .B(_11371_),
    .Y(_04019_));
 AO21x1_ASAP7_75t_R _30949_ (.A1(_02489_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11372_));
 OR3x1_ASAP7_75t_R _30950_ (.A(_02169_),
    .B(_02489_),
    .C(_10978_),
    .Y(_11373_));
 TAPCELL_ASAP7_75t_R PHY_216 ();
 AOI21x1_ASAP7_75t_R _30952_ (.A1(_11003_),
    .A2(_11373_),
    .B(_11360_),
    .Y(_11375_));
 AOI21x1_ASAP7_75t_R _30953_ (.A1(_02169_),
    .A2(_11372_),
    .B(_11375_),
    .Y(_04020_));
 OA211x2_ASAP7_75t_R _30954_ (.A1(_02492_),
    .A2(_10978_),
    .B(_11005_),
    .C(_11363_),
    .Y(_11376_));
 AOI21x1_ASAP7_75t_R _30955_ (.A1(_02168_),
    .A2(_11360_),
    .B(_11376_),
    .Y(_04021_));
 AO21x1_ASAP7_75t_R _30956_ (.A1(_02491_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11377_));
 OR3x1_ASAP7_75t_R _30957_ (.A(_02167_),
    .B(_02491_),
    .C(_10978_),
    .Y(_11378_));
 AOI21x1_ASAP7_75t_R _30958_ (.A1(_11011_),
    .A2(_11378_),
    .B(_11360_),
    .Y(_11379_));
 AOI21x1_ASAP7_75t_R _30959_ (.A1(_02167_),
    .A2(_11377_),
    .B(_11379_),
    .Y(_04022_));
 OA211x2_ASAP7_75t_R _30960_ (.A1(_02494_),
    .A2(_10978_),
    .B(_11013_),
    .C(_11363_),
    .Y(_11380_));
 AOI21x1_ASAP7_75t_R _30961_ (.A1(_02166_),
    .A2(_11360_),
    .B(_11380_),
    .Y(_04023_));
 OR3x1_ASAP7_75t_R _30962_ (.A(_02165_),
    .B(_02493_),
    .C(_10978_),
    .Y(_11381_));
 OAI21x1_ASAP7_75t_R _30963_ (.A1(_09432_),
    .A2(_10986_),
    .B(_11381_),
    .Y(_11382_));
 AO21x1_ASAP7_75t_R _30964_ (.A1(_02493_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11383_));
 AOI22x1_ASAP7_75t_R _30965_ (.A1(_11363_),
    .A2(_11382_),
    .B1(_11383_),
    .B2(_02165_),
    .Y(_04024_));
 OA211x2_ASAP7_75t_R _30966_ (.A1(_02496_),
    .A2(_10978_),
    .B(_11022_),
    .C(_11363_),
    .Y(_11384_));
 AOI21x1_ASAP7_75t_R _30967_ (.A1(_02164_),
    .A2(_11360_),
    .B(_11384_),
    .Y(_04025_));
 AO21x1_ASAP7_75t_R _30968_ (.A1(_02495_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11385_));
 OR3x1_ASAP7_75t_R _30969_ (.A(_02163_),
    .B(_02495_),
    .C(_10978_),
    .Y(_11386_));
 AOI21x1_ASAP7_75t_R _30970_ (.A1(_11026_),
    .A2(_11386_),
    .B(_11360_),
    .Y(_11387_));
 AOI21x1_ASAP7_75t_R _30971_ (.A1(_02163_),
    .A2(_11385_),
    .B(_11387_),
    .Y(_04026_));
 TAPCELL_ASAP7_75t_R PHY_215 ();
 OA211x2_ASAP7_75t_R _30973_ (.A1(_02498_),
    .A2(_10978_),
    .B(_11028_),
    .C(_11363_),
    .Y(_11389_));
 AOI21x1_ASAP7_75t_R _30974_ (.A1(_02162_),
    .A2(_11360_),
    .B(_11389_),
    .Y(_04027_));
 OR3x1_ASAP7_75t_R _30975_ (.A(_02161_),
    .B(_02497_),
    .C(_10978_),
    .Y(_11390_));
 OAI21x1_ASAP7_75t_R _30976_ (.A1(_09458_),
    .A2(_10986_),
    .B(_11390_),
    .Y(_11391_));
 AO21x1_ASAP7_75t_R _30977_ (.A1(_02497_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11392_));
 AOI22x1_ASAP7_75t_R _30978_ (.A1(_11363_),
    .A2(_11391_),
    .B1(_11392_),
    .B2(_02161_),
    .Y(_04028_));
 OA211x2_ASAP7_75t_R _30979_ (.A1(_02500_),
    .A2(_10978_),
    .B(_11035_),
    .C(_11363_),
    .Y(_11393_));
 AOI21x1_ASAP7_75t_R _30980_ (.A1(_02160_),
    .A2(_11360_),
    .B(_11393_),
    .Y(_04029_));
 OR3x1_ASAP7_75t_R _30981_ (.A(_02159_),
    .B(_02499_),
    .C(_10978_),
    .Y(_11394_));
 OAI21x1_ASAP7_75t_R _30982_ (.A1(_09473_),
    .A2(_10986_),
    .B(_11394_),
    .Y(_11395_));
 AO21x1_ASAP7_75t_R _30983_ (.A1(_02499_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11396_));
 AOI22x1_ASAP7_75t_R _30984_ (.A1(_11363_),
    .A2(_11395_),
    .B1(_11396_),
    .B2(_02159_),
    .Y(_04030_));
 OA211x2_ASAP7_75t_R _30985_ (.A1(_02502_),
    .A2(_10978_),
    .B(_11040_),
    .C(_11363_),
    .Y(_11397_));
 AOI21x1_ASAP7_75t_R _30986_ (.A1(_02158_),
    .A2(_11360_),
    .B(_11397_),
    .Y(_04031_));
 AOI21x1_ASAP7_75t_R _30987_ (.A1(_02501_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11398_));
 OR3x1_ASAP7_75t_R _30988_ (.A(_02157_),
    .B(_02501_),
    .C(_10978_),
    .Y(_11399_));
 AO21x1_ASAP7_75t_R _30989_ (.A1(_11044_),
    .A2(_11399_),
    .B(_11360_),
    .Y(_11400_));
 OA21x2_ASAP7_75t_R _30990_ (.A1(_06033_),
    .A2(_11398_),
    .B(_11400_),
    .Y(_04032_));
 OA211x2_ASAP7_75t_R _30991_ (.A1(_02504_),
    .A2(_10978_),
    .B(_11046_),
    .C(_11363_),
    .Y(_11401_));
 AOI21x1_ASAP7_75t_R _30992_ (.A1(_02156_),
    .A2(_11360_),
    .B(_11401_),
    .Y(_04033_));
 OR3x1_ASAP7_75t_R _30993_ (.A(_02155_),
    .B(_02503_),
    .C(_10978_),
    .Y(_11402_));
 OAI21x1_ASAP7_75t_R _30994_ (.A1(_09503_),
    .A2(_10986_),
    .B(_11402_),
    .Y(_11403_));
 AO21x1_ASAP7_75t_R _30995_ (.A1(_02503_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11404_));
 AOI22x1_ASAP7_75t_R _30996_ (.A1(_11363_),
    .A2(_11403_),
    .B1(_11404_),
    .B2(_02155_),
    .Y(_04034_));
 OA211x2_ASAP7_75t_R _30997_ (.A1(_02506_),
    .A2(_10978_),
    .B(_11052_),
    .C(_11363_),
    .Y(_11405_));
 AOI21x1_ASAP7_75t_R _30998_ (.A1(_02154_),
    .A2(_11360_),
    .B(_11405_),
    .Y(_04035_));
 NOR2x1_ASAP7_75t_R _30999_ (.A(_02153_),
    .B(_02505_),
    .Y(_11406_));
 AO21x1_ASAP7_75t_R _31000_ (.A1(_10986_),
    .A2(_11406_),
    .B(_11056_),
    .Y(_11407_));
 AO21x1_ASAP7_75t_R _31001_ (.A1(_02505_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11408_));
 AOI22x1_ASAP7_75t_R _31002_ (.A1(_11363_),
    .A2(_11407_),
    .B1(_11408_),
    .B2(_02153_),
    .Y(_04036_));
 OA211x2_ASAP7_75t_R _31003_ (.A1(_02508_),
    .A2(_10978_),
    .B(_11060_),
    .C(_11363_),
    .Y(_11409_));
 AOI21x1_ASAP7_75t_R _31004_ (.A1(_02152_),
    .A2(_11360_),
    .B(_11409_),
    .Y(_04037_));
 NOR2x1_ASAP7_75t_R _31005_ (.A(_02151_),
    .B(_02507_),
    .Y(_11410_));
 AO21x1_ASAP7_75t_R _31006_ (.A1(_10986_),
    .A2(_11410_),
    .B(_11063_),
    .Y(_11411_));
 AO21x1_ASAP7_75t_R _31007_ (.A1(_02507_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11412_));
 AOI22x1_ASAP7_75t_R _31008_ (.A1(_11363_),
    .A2(_11411_),
    .B1(_11412_),
    .B2(_02151_),
    .Y(_04038_));
 OA211x2_ASAP7_75t_R _31009_ (.A1(_02510_),
    .A2(_10978_),
    .B(_11066_),
    .C(_11363_),
    .Y(_11413_));
 AOI21x1_ASAP7_75t_R _31010_ (.A1(_02150_),
    .A2(_11360_),
    .B(_11413_),
    .Y(_04039_));
 OR3x1_ASAP7_75t_R _31011_ (.A(_02149_),
    .B(_02509_),
    .C(_10978_),
    .Y(_11414_));
 OAI21x1_ASAP7_75t_R _31012_ (.A1(_09545_),
    .A2(_10986_),
    .B(_11414_),
    .Y(_11415_));
 AO21x1_ASAP7_75t_R _31013_ (.A1(_02509_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11416_));
 AOI22x1_ASAP7_75t_R _31014_ (.A1(_11363_),
    .A2(_11415_),
    .B1(_11416_),
    .B2(_02149_),
    .Y(_04040_));
 OR2x2_ASAP7_75t_R _31015_ (.A(_02512_),
    .B(_10978_),
    .Y(_11417_));
 OA211x2_ASAP7_75t_R _31016_ (.A1(_09560_),
    .A2(_11020_),
    .B(_11363_),
    .C(_11417_),
    .Y(_11418_));
 AOI21x1_ASAP7_75t_R _31017_ (.A1(_02148_),
    .A2(_11360_),
    .B(_11418_),
    .Y(_04041_));
 OR3x1_ASAP7_75t_R _31018_ (.A(_02147_),
    .B(_02511_),
    .C(_10978_),
    .Y(_11419_));
 OAI21x1_ASAP7_75t_R _31019_ (.A1(_09565_),
    .A2(_10986_),
    .B(_11419_),
    .Y(_11420_));
 AO21x1_ASAP7_75t_R _31020_ (.A1(_02511_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11421_));
 AOI22x1_ASAP7_75t_R _31021_ (.A1(_11363_),
    .A2(_11420_),
    .B1(_11421_),
    .B2(_02147_),
    .Y(_04042_));
 OA211x2_ASAP7_75t_R _31022_ (.A1(_02514_),
    .A2(_10978_),
    .B(_11076_),
    .C(_11363_),
    .Y(_11422_));
 AOI21x1_ASAP7_75t_R _31023_ (.A1(_02146_),
    .A2(_11360_),
    .B(_11422_),
    .Y(_04043_));
 OR3x1_ASAP7_75t_R _31024_ (.A(_02145_),
    .B(_02513_),
    .C(_10978_),
    .Y(_11423_));
 OAI21x1_ASAP7_75t_R _31025_ (.A1(_09578_),
    .A2(_10986_),
    .B(_11423_),
    .Y(_11424_));
 AO21x1_ASAP7_75t_R _31026_ (.A1(_02513_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11425_));
 AOI22x1_ASAP7_75t_R _31027_ (.A1(_11363_),
    .A2(_11424_),
    .B1(_11425_),
    .B2(_02145_),
    .Y(_04044_));
 OA211x2_ASAP7_75t_R _31028_ (.A1(_02516_),
    .A2(_10978_),
    .B(_11081_),
    .C(_11363_),
    .Y(_11426_));
 AOI21x1_ASAP7_75t_R _31029_ (.A1(_02144_),
    .A2(_11360_),
    .B(_11426_),
    .Y(_04045_));
 AOI21x1_ASAP7_75t_R _31030_ (.A1(_02515_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11427_));
 OR3x1_ASAP7_75t_R _31031_ (.A(_02143_),
    .B(_02515_),
    .C(_10978_),
    .Y(_11428_));
 AO21x1_ASAP7_75t_R _31032_ (.A1(_11085_),
    .A2(_11428_),
    .B(_11360_),
    .Y(_11429_));
 OA21x2_ASAP7_75t_R _31033_ (.A1(_06040_),
    .A2(_11427_),
    .B(_11429_),
    .Y(_04046_));
 OA211x2_ASAP7_75t_R _31034_ (.A1(_02518_),
    .A2(_10978_),
    .B(_11087_),
    .C(_11363_),
    .Y(_11430_));
 AOI21x1_ASAP7_75t_R _31035_ (.A1(_02142_),
    .A2(_11360_),
    .B(_11430_),
    .Y(_04047_));
 OR3x1_ASAP7_75t_R _31036_ (.A(_02141_),
    .B(_02517_),
    .C(_10978_),
    .Y(_11431_));
 OAI21x1_ASAP7_75t_R _31037_ (.A1(_09605_),
    .A2(_10986_),
    .B(_11431_),
    .Y(_11432_));
 AO21x1_ASAP7_75t_R _31038_ (.A1(_02517_),
    .A2(_10986_),
    .B(_11360_),
    .Y(_11433_));
 AOI22x1_ASAP7_75t_R _31039_ (.A1(_11363_),
    .A2(_11432_),
    .B1(_11433_),
    .B2(_02141_),
    .Y(_04048_));
 AOI21x1_ASAP7_75t_R _31040_ (.A1(_05705_),
    .A2(_05712_),
    .B(_06257_),
    .Y(_11434_));
 NOR2x1_ASAP7_75t_R _31041_ (.A(_02140_),
    .B(_11434_),
    .Y(_11435_));
 INVx1_ASAP7_75t_R _31042_ (.A(_01577_),
    .Y(_11436_));
 NAND2x1_ASAP7_75t_R _31043_ (.A(_01456_),
    .B(_06258_),
    .Y(_11437_));
 OA211x2_ASAP7_75t_R _31044_ (.A1(_11436_),
    .A2(_06258_),
    .B(_11434_),
    .C(_11437_),
    .Y(_11438_));
 OR3x1_ASAP7_75t_R _31045_ (.A(_11224_),
    .B(_11435_),
    .C(_11438_),
    .Y(_04049_));
 NOR2x1_ASAP7_75t_R _31046_ (.A(_17592_),
    .B(_11434_),
    .Y(_11439_));
 INVx1_ASAP7_75t_R _31047_ (.A(_01576_),
    .Y(_11440_));
 NAND2x1_ASAP7_75t_R _31048_ (.A(_01455_),
    .B(_06258_),
    .Y(_11441_));
 OA211x2_ASAP7_75t_R _31049_ (.A1(_11440_),
    .A2(_06258_),
    .B(_11434_),
    .C(_11441_),
    .Y(_11442_));
 OR3x1_ASAP7_75t_R _31050_ (.A(_11224_),
    .B(_11439_),
    .C(_11442_),
    .Y(_04050_));
 INVx1_ASAP7_75t_R _31051_ (.A(_09365_),
    .Y(_11443_));
 OR3x4_ASAP7_75t_R _31052_ (.A(_06908_),
    .B(_07507_),
    .C(_11443_),
    .Y(_11444_));
 TAPCELL_ASAP7_75t_R PHY_214 ();
 TAPCELL_ASAP7_75t_R PHY_213 ();
 TAPCELL_ASAP7_75t_R PHY_212 ();
 NAND2x1_ASAP7_75t_R _31056_ (.A(_02139_),
    .B(_11444_),
    .Y(_11448_));
 OA21x2_ASAP7_75t_R _31057_ (.A1(_10974_),
    .A2(_11444_),
    .B(_11448_),
    .Y(_04051_));
 NAND2x1_ASAP7_75t_R _31058_ (.A(_02138_),
    .B(_11444_),
    .Y(_11449_));
 OA21x2_ASAP7_75t_R _31059_ (.A1(_09363_),
    .A2(_11444_),
    .B(_11449_),
    .Y(_04052_));
 NAND2x1_ASAP7_75t_R _31060_ (.A(_02137_),
    .B(_11444_),
    .Y(_11450_));
 OA21x2_ASAP7_75t_R _31061_ (.A1(_09390_),
    .A2(_11444_),
    .B(_11450_),
    .Y(_04053_));
 NAND2x1_ASAP7_75t_R _31062_ (.A(_02136_),
    .B(_11444_),
    .Y(_11451_));
 OA21x2_ASAP7_75t_R _31063_ (.A1(_09397_),
    .A2(_11444_),
    .B(_11451_),
    .Y(_04054_));
 NAND2x1_ASAP7_75t_R _31064_ (.A(_02135_),
    .B(_11444_),
    .Y(_11452_));
 OA21x2_ASAP7_75t_R _31065_ (.A1(_09408_),
    .A2(_11444_),
    .B(_11452_),
    .Y(_04055_));
 NAND2x1_ASAP7_75t_R _31066_ (.A(_02134_),
    .B(_11444_),
    .Y(_11453_));
 OA21x2_ASAP7_75t_R _31067_ (.A1(_09417_),
    .A2(_11444_),
    .B(_11453_),
    .Y(_04056_));
 NAND2x1_ASAP7_75t_R _31068_ (.A(_02133_),
    .B(_11444_),
    .Y(_11454_));
 OA21x2_ASAP7_75t_R _31069_ (.A1(_09426_),
    .A2(_11444_),
    .B(_11454_),
    .Y(_04057_));
 NAND2x1_ASAP7_75t_R _31070_ (.A(_02132_),
    .B(_11444_),
    .Y(_11455_));
 OA21x2_ASAP7_75t_R _31071_ (.A1(_09432_),
    .A2(_11444_),
    .B(_11455_),
    .Y(_04058_));
 TAPCELL_ASAP7_75t_R PHY_211 ();
 NAND2x1_ASAP7_75t_R _31073_ (.A(_02131_),
    .B(_11444_),
    .Y(_11457_));
 OA21x2_ASAP7_75t_R _31074_ (.A1(_09438_),
    .A2(_11444_),
    .B(_11457_),
    .Y(_04059_));
 NAND2x1_ASAP7_75t_R _31075_ (.A(_02130_),
    .B(_11444_),
    .Y(_11458_));
 OA21x2_ASAP7_75t_R _31076_ (.A1(_09445_),
    .A2(_11444_),
    .B(_11458_),
    .Y(_04060_));
 TAPCELL_ASAP7_75t_R PHY_210 ();
 NAND2x1_ASAP7_75t_R _31078_ (.A(_02129_),
    .B(_11444_),
    .Y(_11460_));
 OA21x2_ASAP7_75t_R _31079_ (.A1(_09452_),
    .A2(_11444_),
    .B(_11460_),
    .Y(_04061_));
 NAND2x1_ASAP7_75t_R _31080_ (.A(_02128_),
    .B(_11444_),
    .Y(_11461_));
 OA21x2_ASAP7_75t_R _31081_ (.A1(_09458_),
    .A2(_11444_),
    .B(_11461_),
    .Y(_04062_));
 NAND2x1_ASAP7_75t_R _31082_ (.A(_02127_),
    .B(_11444_),
    .Y(_11462_));
 OA21x2_ASAP7_75t_R _31083_ (.A1(_09465_),
    .A2(_11444_),
    .B(_11462_),
    .Y(_04063_));
 NAND2x1_ASAP7_75t_R _31084_ (.A(_02126_),
    .B(_11444_),
    .Y(_11463_));
 OA21x2_ASAP7_75t_R _31085_ (.A1(_09473_),
    .A2(_11444_),
    .B(_11463_),
    .Y(_04064_));
 NAND2x1_ASAP7_75t_R _31086_ (.A(_02125_),
    .B(_11444_),
    .Y(_11464_));
 OA21x2_ASAP7_75t_R _31087_ (.A1(_09481_),
    .A2(_11444_),
    .B(_11464_),
    .Y(_04065_));
 NAND2x1_ASAP7_75t_R _31088_ (.A(_02124_),
    .B(_11444_),
    .Y(_11465_));
 OA21x2_ASAP7_75t_R _31089_ (.A1(_09488_),
    .A2(_11444_),
    .B(_11465_),
    .Y(_04066_));
 NAND2x1_ASAP7_75t_R _31090_ (.A(_02123_),
    .B(_11444_),
    .Y(_11466_));
 OA21x2_ASAP7_75t_R _31091_ (.A1(_09496_),
    .A2(_11444_),
    .B(_11466_),
    .Y(_04067_));
 NAND2x1_ASAP7_75t_R _31092_ (.A(_02122_),
    .B(_11444_),
    .Y(_11467_));
 OA21x2_ASAP7_75t_R _31093_ (.A1(_09503_),
    .A2(_11444_),
    .B(_11467_),
    .Y(_04068_));
 TAPCELL_ASAP7_75t_R PHY_209 ();
 NAND2x1_ASAP7_75t_R _31095_ (.A(_02121_),
    .B(_11444_),
    .Y(_11469_));
 OA21x2_ASAP7_75t_R _31096_ (.A1(_09512_),
    .A2(_11444_),
    .B(_11469_),
    .Y(_04069_));
 NAND2x1_ASAP7_75t_R _31097_ (.A(_02120_),
    .B(_11444_),
    .Y(_11470_));
 OA21x2_ASAP7_75t_R _31098_ (.A1(_09519_),
    .A2(_11444_),
    .B(_11470_),
    .Y(_04070_));
 TAPCELL_ASAP7_75t_R PHY_208 ();
 NAND2x1_ASAP7_75t_R _31100_ (.A(_02119_),
    .B(_11444_),
    .Y(_11472_));
 OA21x2_ASAP7_75t_R _31101_ (.A1(_09526_),
    .A2(_11444_),
    .B(_11472_),
    .Y(_04071_));
 NAND2x1_ASAP7_75t_R _31102_ (.A(_02118_),
    .B(_11444_),
    .Y(_11473_));
 OA21x2_ASAP7_75t_R _31103_ (.A1(_09532_),
    .A2(_11444_),
    .B(_11473_),
    .Y(_04072_));
 NAND2x1_ASAP7_75t_R _31104_ (.A(_02117_),
    .B(_11444_),
    .Y(_11474_));
 OA21x2_ASAP7_75t_R _31105_ (.A1(_09539_),
    .A2(_11444_),
    .B(_11474_),
    .Y(_04073_));
 NAND2x1_ASAP7_75t_R _31106_ (.A(_02116_),
    .B(_11444_),
    .Y(_11475_));
 OA21x2_ASAP7_75t_R _31107_ (.A1(_09545_),
    .A2(_11444_),
    .B(_11475_),
    .Y(_04074_));
 NAND2x1_ASAP7_75t_R _31108_ (.A(_02115_),
    .B(_11444_),
    .Y(_11476_));
 OA21x2_ASAP7_75t_R _31109_ (.A1(_11192_),
    .A2(_11444_),
    .B(_11476_),
    .Y(_04075_));
 NAND2x1_ASAP7_75t_R _31110_ (.A(_02114_),
    .B(_11444_),
    .Y(_11477_));
 OA21x2_ASAP7_75t_R _31111_ (.A1(_09565_),
    .A2(_11444_),
    .B(_11477_),
    .Y(_04076_));
 NAND2x1_ASAP7_75t_R _31112_ (.A(_02113_),
    .B(_11444_),
    .Y(_11478_));
 OA21x2_ASAP7_75t_R _31113_ (.A1(_09572_),
    .A2(_11444_),
    .B(_11478_),
    .Y(_04077_));
 NAND2x1_ASAP7_75t_R _31114_ (.A(_02112_),
    .B(_11444_),
    .Y(_11479_));
 OA21x2_ASAP7_75t_R _31115_ (.A1(_09578_),
    .A2(_11444_),
    .B(_11479_),
    .Y(_04078_));
 NAND2x1_ASAP7_75t_R _31116_ (.A(_02111_),
    .B(_11444_),
    .Y(_11480_));
 OA21x2_ASAP7_75t_R _31117_ (.A1(_09585_),
    .A2(_11444_),
    .B(_11480_),
    .Y(_04079_));
 NAND2x1_ASAP7_75t_R _31118_ (.A(_02110_),
    .B(_11444_),
    .Y(_11481_));
 OA21x2_ASAP7_75t_R _31119_ (.A1(_09591_),
    .A2(_11444_),
    .B(_11481_),
    .Y(_04080_));
 NAND2x1_ASAP7_75t_R _31120_ (.A(_02109_),
    .B(_11444_),
    .Y(_11482_));
 OA21x2_ASAP7_75t_R _31121_ (.A1(_09598_),
    .A2(_11444_),
    .B(_11482_),
    .Y(_04081_));
 NAND2x1_ASAP7_75t_R _31122_ (.A(_02108_),
    .B(_11444_),
    .Y(_11483_));
 OA21x2_ASAP7_75t_R _31123_ (.A1(_09605_),
    .A2(_11444_),
    .B(_11483_),
    .Y(_04082_));
 TAPCELL_ASAP7_75t_R PHY_207 ();
 TAPCELL_ASAP7_75t_R PHY_206 ();
 TAPCELL_ASAP7_75t_R PHY_205 ();
 AND2x2_ASAP7_75t_R _31127_ (.A(_01456_),
    .B(_11242_),
    .Y(_11487_));
 AOI21x1_ASAP7_75t_R _31128_ (.A1(_02107_),
    .A2(_11226_),
    .B(_11487_),
    .Y(_04083_));
 AND2x2_ASAP7_75t_R _31129_ (.A(_01455_),
    .B(_11242_),
    .Y(_11488_));
 AOI21x1_ASAP7_75t_R _31130_ (.A1(_02106_),
    .A2(_11226_),
    .B(_11488_),
    .Y(_04084_));
 AND2x2_ASAP7_75t_R _31131_ (.A(_01454_),
    .B(_11242_),
    .Y(_11489_));
 AOI21x1_ASAP7_75t_R _31132_ (.A1(_02105_),
    .A2(_11226_),
    .B(_11489_),
    .Y(_04085_));
 AND2x2_ASAP7_75t_R _31133_ (.A(_01913_),
    .B(_11242_),
    .Y(_11490_));
 AOI21x1_ASAP7_75t_R _31134_ (.A1(_02104_),
    .A2(_11226_),
    .B(_11490_),
    .Y(_04086_));
 AND2x2_ASAP7_75t_R _31135_ (.A(_01912_),
    .B(_11242_),
    .Y(_11491_));
 AOI21x1_ASAP7_75t_R _31136_ (.A1(_02103_),
    .A2(_11226_),
    .B(_11491_),
    .Y(_04087_));
 AND2x2_ASAP7_75t_R _31137_ (.A(_01911_),
    .B(_11242_),
    .Y(_11492_));
 AOI21x1_ASAP7_75t_R _31138_ (.A1(_02102_),
    .A2(_11226_),
    .B(_11492_),
    .Y(_04088_));
 INVx1_ASAP7_75t_R _31139_ (.A(_02101_),
    .Y(_11493_));
 NAND2x1_ASAP7_75t_R _31140_ (.A(_01910_),
    .B(_11242_),
    .Y(_11494_));
 OA21x2_ASAP7_75t_R _31141_ (.A1(_11493_),
    .A2(_11242_),
    .B(_11494_),
    .Y(_04089_));
 AND2x2_ASAP7_75t_R _31142_ (.A(_01909_),
    .B(_11242_),
    .Y(_11495_));
 AOI21x1_ASAP7_75t_R _31143_ (.A1(_02100_),
    .A2(_11226_),
    .B(_11495_),
    .Y(_04090_));
 AND2x2_ASAP7_75t_R _31144_ (.A(_01908_),
    .B(_11242_),
    .Y(_11496_));
 AOI21x1_ASAP7_75t_R _31145_ (.A1(_02099_),
    .A2(_11226_),
    .B(_11496_),
    .Y(_04091_));
 AND5x2_ASAP7_75t_R _31146_ (.A(_14497_),
    .B(_05572_),
    .C(_05606_),
    .D(_05611_),
    .E(_09365_),
    .Y(_11497_));
 INVx1_ASAP7_75t_R _31147_ (.A(_11497_),
    .Y(_11498_));
 OR4x2_ASAP7_75t_R _31148_ (.A(_13301_),
    .B(_05560_),
    .C(_05685_),
    .D(_11498_),
    .Y(_11499_));
 TAPCELL_ASAP7_75t_R PHY_204 ();
 TAPCELL_ASAP7_75t_R PHY_203 ();
 TAPCELL_ASAP7_75t_R PHY_202 ();
 NAND2x1_ASAP7_75t_R _31152_ (.A(_02098_),
    .B(_11499_),
    .Y(_11503_));
 OA21x2_ASAP7_75t_R _31153_ (.A1(_10974_),
    .A2(_11499_),
    .B(_11503_),
    .Y(_04092_));
 NAND2x1_ASAP7_75t_R _31154_ (.A(_02097_),
    .B(_11499_),
    .Y(_11504_));
 OA21x2_ASAP7_75t_R _31155_ (.A1(_09363_),
    .A2(_11499_),
    .B(_11504_),
    .Y(_04093_));
 NAND2x1_ASAP7_75t_R _31156_ (.A(_02096_),
    .B(_11499_),
    .Y(_11505_));
 OA21x2_ASAP7_75t_R _31157_ (.A1(_09390_),
    .A2(_11499_),
    .B(_11505_),
    .Y(_04094_));
 NAND2x1_ASAP7_75t_R _31158_ (.A(_02095_),
    .B(_11499_),
    .Y(_11506_));
 OA21x2_ASAP7_75t_R _31159_ (.A1(_09397_),
    .A2(_11499_),
    .B(_11506_),
    .Y(_04095_));
 NAND2x1_ASAP7_75t_R _31160_ (.A(_02094_),
    .B(_11499_),
    .Y(_11507_));
 OA21x2_ASAP7_75t_R _31161_ (.A1(_09408_),
    .A2(_11499_),
    .B(_11507_),
    .Y(_04096_));
 NAND2x1_ASAP7_75t_R _31162_ (.A(_02093_),
    .B(_11499_),
    .Y(_11508_));
 OA21x2_ASAP7_75t_R _31163_ (.A1(_09417_),
    .A2(_11499_),
    .B(_11508_),
    .Y(_04097_));
 NAND2x1_ASAP7_75t_R _31164_ (.A(_02092_),
    .B(_11499_),
    .Y(_11509_));
 OA21x2_ASAP7_75t_R _31165_ (.A1(_09426_),
    .A2(_11499_),
    .B(_11509_),
    .Y(_04098_));
 NAND2x1_ASAP7_75t_R _31166_ (.A(_02091_),
    .B(_11499_),
    .Y(_11510_));
 OA21x2_ASAP7_75t_R _31167_ (.A1(_09432_),
    .A2(_11499_),
    .B(_11510_),
    .Y(_04099_));
 TAPCELL_ASAP7_75t_R PHY_201 ();
 NAND2x1_ASAP7_75t_R _31169_ (.A(_02090_),
    .B(_11499_),
    .Y(_11512_));
 OA21x2_ASAP7_75t_R _31170_ (.A1(_09438_),
    .A2(_11499_),
    .B(_11512_),
    .Y(_04100_));
 NAND2x1_ASAP7_75t_R _31171_ (.A(_02089_),
    .B(_11499_),
    .Y(_11513_));
 OA21x2_ASAP7_75t_R _31172_ (.A1(_09445_),
    .A2(_11499_),
    .B(_11513_),
    .Y(_04101_));
 TAPCELL_ASAP7_75t_R PHY_200 ();
 NAND2x1_ASAP7_75t_R _31174_ (.A(_02088_),
    .B(_11499_),
    .Y(_11515_));
 OA21x2_ASAP7_75t_R _31175_ (.A1(_09452_),
    .A2(_11499_),
    .B(_11515_),
    .Y(_04102_));
 NAND2x1_ASAP7_75t_R _31176_ (.A(_02087_),
    .B(_11499_),
    .Y(_11516_));
 OA21x2_ASAP7_75t_R _31177_ (.A1(_09458_),
    .A2(_11499_),
    .B(_11516_),
    .Y(_04103_));
 NAND2x1_ASAP7_75t_R _31178_ (.A(_02086_),
    .B(_11499_),
    .Y(_11517_));
 OA21x2_ASAP7_75t_R _31179_ (.A1(_09465_),
    .A2(_11499_),
    .B(_11517_),
    .Y(_04104_));
 NAND2x1_ASAP7_75t_R _31180_ (.A(_02085_),
    .B(_11499_),
    .Y(_11518_));
 OA21x2_ASAP7_75t_R _31181_ (.A1(_09473_),
    .A2(_11499_),
    .B(_11518_),
    .Y(_04105_));
 NAND2x1_ASAP7_75t_R _31182_ (.A(_02084_),
    .B(_11499_),
    .Y(_11519_));
 OA21x2_ASAP7_75t_R _31183_ (.A1(_09481_),
    .A2(_11499_),
    .B(_11519_),
    .Y(_04106_));
 NAND2x1_ASAP7_75t_R _31184_ (.A(_02083_),
    .B(_11499_),
    .Y(_11520_));
 OA21x2_ASAP7_75t_R _31185_ (.A1(_09488_),
    .A2(_11499_),
    .B(_11520_),
    .Y(_04107_));
 NAND2x1_ASAP7_75t_R _31186_ (.A(_02082_),
    .B(_11499_),
    .Y(_11521_));
 OA21x2_ASAP7_75t_R _31187_ (.A1(_09496_),
    .A2(_11499_),
    .B(_11521_),
    .Y(_04108_));
 NAND2x1_ASAP7_75t_R _31188_ (.A(_02081_),
    .B(_11499_),
    .Y(_11522_));
 OA21x2_ASAP7_75t_R _31189_ (.A1(_09503_),
    .A2(_11499_),
    .B(_11522_),
    .Y(_04109_));
 TAPCELL_ASAP7_75t_R PHY_199 ();
 NAND2x1_ASAP7_75t_R _31191_ (.A(_02080_),
    .B(_11499_),
    .Y(_11524_));
 OA21x2_ASAP7_75t_R _31192_ (.A1(_09512_),
    .A2(_11499_),
    .B(_11524_),
    .Y(_04110_));
 NAND2x1_ASAP7_75t_R _31193_ (.A(_02079_),
    .B(_11499_),
    .Y(_11525_));
 OA21x2_ASAP7_75t_R _31194_ (.A1(_09519_),
    .A2(_11499_),
    .B(_11525_),
    .Y(_04111_));
 TAPCELL_ASAP7_75t_R PHY_198 ();
 NAND2x1_ASAP7_75t_R _31196_ (.A(_02078_),
    .B(_11499_),
    .Y(_11527_));
 OA21x2_ASAP7_75t_R _31197_ (.A1(_09526_),
    .A2(_11499_),
    .B(_11527_),
    .Y(_04112_));
 NAND2x1_ASAP7_75t_R _31198_ (.A(_02077_),
    .B(_11499_),
    .Y(_11528_));
 OA21x2_ASAP7_75t_R _31199_ (.A1(_09532_),
    .A2(_11499_),
    .B(_11528_),
    .Y(_04113_));
 NAND2x1_ASAP7_75t_R _31200_ (.A(_02076_),
    .B(_11499_),
    .Y(_11529_));
 OA21x2_ASAP7_75t_R _31201_ (.A1(_09539_),
    .A2(_11499_),
    .B(_11529_),
    .Y(_04114_));
 NAND2x1_ASAP7_75t_R _31202_ (.A(_02075_),
    .B(_11499_),
    .Y(_11530_));
 OA21x2_ASAP7_75t_R _31203_ (.A1(_09545_),
    .A2(_11499_),
    .B(_11530_),
    .Y(_04115_));
 NAND2x1_ASAP7_75t_R _31204_ (.A(_02074_),
    .B(_11499_),
    .Y(_11531_));
 OA21x2_ASAP7_75t_R _31205_ (.A1(_11192_),
    .A2(_11499_),
    .B(_11531_),
    .Y(_04116_));
 NAND2x1_ASAP7_75t_R _31206_ (.A(_02073_),
    .B(_11499_),
    .Y(_11532_));
 OA21x2_ASAP7_75t_R _31207_ (.A1(_09565_),
    .A2(_11499_),
    .B(_11532_),
    .Y(_04117_));
 NAND2x1_ASAP7_75t_R _31208_ (.A(_02072_),
    .B(_11499_),
    .Y(_11533_));
 OA21x2_ASAP7_75t_R _31209_ (.A1(_09572_),
    .A2(_11499_),
    .B(_11533_),
    .Y(_04118_));
 NAND2x1_ASAP7_75t_R _31210_ (.A(_02071_),
    .B(_11499_),
    .Y(_11534_));
 OA21x2_ASAP7_75t_R _31211_ (.A1(_09578_),
    .A2(_11499_),
    .B(_11534_),
    .Y(_04119_));
 NAND2x1_ASAP7_75t_R _31212_ (.A(_02070_),
    .B(_11499_),
    .Y(_11535_));
 OA21x2_ASAP7_75t_R _31213_ (.A1(_09585_),
    .A2(_11499_),
    .B(_11535_),
    .Y(_04120_));
 NAND2x1_ASAP7_75t_R _31214_ (.A(_02069_),
    .B(_11499_),
    .Y(_11536_));
 OA21x2_ASAP7_75t_R _31215_ (.A1(_09591_),
    .A2(_11499_),
    .B(_11536_),
    .Y(_04121_));
 NAND2x1_ASAP7_75t_R _31216_ (.A(_02068_),
    .B(_11499_),
    .Y(_11537_));
 OA21x2_ASAP7_75t_R _31217_ (.A1(_09598_),
    .A2(_11499_),
    .B(_11537_),
    .Y(_04122_));
 NAND2x1_ASAP7_75t_R _31218_ (.A(_02067_),
    .B(_11499_),
    .Y(_11538_));
 OA21x2_ASAP7_75t_R _31219_ (.A1(_09605_),
    .A2(_11499_),
    .B(_11538_),
    .Y(_04123_));
 INVx1_ASAP7_75t_R _31220_ (.A(_00095_),
    .Y(_11539_));
 AND3x4_ASAP7_75t_R _31221_ (.A(_01714_),
    .B(_01715_),
    .C(_01716_),
    .Y(_11540_));
 NAND2x1_ASAP7_75t_R _31222_ (.A(_05632_),
    .B(_09353_),
    .Y(_11541_));
 NOR2x2_ASAP7_75t_R _31223_ (.A(_07150_),
    .B(_11541_),
    .Y(_11542_));
 NOR2x2_ASAP7_75t_R _31224_ (.A(_11540_),
    .B(_11542_),
    .Y(_11543_));
 TAPCELL_ASAP7_75t_R PHY_197 ();
 TAPCELL_ASAP7_75t_R PHY_196 ();
 TAPCELL_ASAP7_75t_R PHY_195 ();
 AO22x1_ASAP7_75t_R _31228_ (.A1(net23),
    .A2(_11540_),
    .B1(_09438_),
    .B2(_11542_),
    .Y(_11547_));
 AO21x1_ASAP7_75t_R _31229_ (.A1(_11539_),
    .A2(_11543_),
    .B(_11547_),
    .Y(_04124_));
 INVx1_ASAP7_75t_R _31230_ (.A(_00098_),
    .Y(_11548_));
 AO22x1_ASAP7_75t_R _31231_ (.A1(net24),
    .A2(_11540_),
    .B1(_09445_),
    .B2(_11542_),
    .Y(_11549_));
 AO21x1_ASAP7_75t_R _31232_ (.A1(_11548_),
    .A2(_11543_),
    .B(_11549_),
    .Y(_04125_));
 INVx1_ASAP7_75t_R _31233_ (.A(_00101_),
    .Y(_11550_));
 AO22x1_ASAP7_75t_R _31234_ (.A1(net1),
    .A2(_11540_),
    .B1(_09452_),
    .B2(_11542_),
    .Y(_11551_));
 AO21x1_ASAP7_75t_R _31235_ (.A1(_11550_),
    .A2(_11543_),
    .B(_11551_),
    .Y(_04126_));
 INVx1_ASAP7_75t_R _31236_ (.A(_00657_),
    .Y(_11552_));
 AO22x1_ASAP7_75t_R _31237_ (.A1(net2),
    .A2(_11540_),
    .B1(_09458_),
    .B2(_11542_),
    .Y(_11553_));
 AO21x1_ASAP7_75t_R _31238_ (.A1(_11552_),
    .A2(_11543_),
    .B(_11553_),
    .Y(_04127_));
 INVx1_ASAP7_75t_R _31239_ (.A(_00656_),
    .Y(_11554_));
 AO22x1_ASAP7_75t_R _31240_ (.A1(net3),
    .A2(_11540_),
    .B1(_09465_),
    .B2(_11542_),
    .Y(_11555_));
 AO21x1_ASAP7_75t_R _31241_ (.A1(_11554_),
    .A2(_11543_),
    .B(_11555_),
    .Y(_04128_));
 INVx1_ASAP7_75t_R _31242_ (.A(_00108_),
    .Y(_11556_));
 AO22x1_ASAP7_75t_R _31243_ (.A1(net4),
    .A2(_11540_),
    .B1(_09473_),
    .B2(_11542_),
    .Y(_11557_));
 AO21x1_ASAP7_75t_R _31244_ (.A1(_11556_),
    .A2(_11543_),
    .B(_11557_),
    .Y(_04129_));
 INVx1_ASAP7_75t_R _31245_ (.A(_00111_),
    .Y(_11558_));
 AO22x1_ASAP7_75t_R _31246_ (.A1(net5),
    .A2(_11540_),
    .B1(_09481_),
    .B2(_11542_),
    .Y(_11559_));
 AO21x1_ASAP7_75t_R _31247_ (.A1(_11558_),
    .A2(_11543_),
    .B(_11559_),
    .Y(_04130_));
 INVx1_ASAP7_75t_R _31248_ (.A(_00114_),
    .Y(_11560_));
 AO22x1_ASAP7_75t_R _31249_ (.A1(net6),
    .A2(_11540_),
    .B1(_09488_),
    .B2(_11542_),
    .Y(_11561_));
 AO21x1_ASAP7_75t_R _31250_ (.A1(_11560_),
    .A2(_11543_),
    .B(_11561_),
    .Y(_04131_));
 INVx1_ASAP7_75t_R _31251_ (.A(_00117_),
    .Y(_11562_));
 AO22x1_ASAP7_75t_R _31252_ (.A1(net7),
    .A2(_11540_),
    .B1(_09496_),
    .B2(_11542_),
    .Y(_11563_));
 AO21x1_ASAP7_75t_R _31253_ (.A1(_11562_),
    .A2(_11543_),
    .B(_11563_),
    .Y(_04132_));
 INVx1_ASAP7_75t_R _31254_ (.A(_00120_),
    .Y(_11564_));
 AO22x1_ASAP7_75t_R _31255_ (.A1(net8),
    .A2(_11540_),
    .B1(_09503_),
    .B2(_11542_),
    .Y(_11565_));
 AO21x1_ASAP7_75t_R _31256_ (.A1(_11564_),
    .A2(_11543_),
    .B(_11565_),
    .Y(_04133_));
 INVx1_ASAP7_75t_R _31257_ (.A(_00123_),
    .Y(_11566_));
 TAPCELL_ASAP7_75t_R PHY_194 ();
 TAPCELL_ASAP7_75t_R PHY_193 ();
 TAPCELL_ASAP7_75t_R PHY_192 ();
 AO22x1_ASAP7_75t_R _31261_ (.A1(net9),
    .A2(_11540_),
    .B1(_09512_),
    .B2(_11542_),
    .Y(_11570_));
 AO21x1_ASAP7_75t_R _31262_ (.A1(_11566_),
    .A2(_11543_),
    .B(_11570_),
    .Y(_04134_));
 INVx1_ASAP7_75t_R _31263_ (.A(_00126_),
    .Y(_11571_));
 AO22x1_ASAP7_75t_R _31264_ (.A1(net10),
    .A2(_11540_),
    .B1(_09519_),
    .B2(_11542_),
    .Y(_11572_));
 AO21x1_ASAP7_75t_R _31265_ (.A1(_11571_),
    .A2(_11543_),
    .B(_11572_),
    .Y(_04135_));
 INVx1_ASAP7_75t_R _31266_ (.A(_00129_),
    .Y(_11573_));
 AO22x1_ASAP7_75t_R _31267_ (.A1(net11),
    .A2(_11540_),
    .B1(_09526_),
    .B2(_11542_),
    .Y(_11574_));
 AO21x1_ASAP7_75t_R _31268_ (.A1(_11573_),
    .A2(_11543_),
    .B(_11574_),
    .Y(_04136_));
 INVx1_ASAP7_75t_R _31269_ (.A(_00132_),
    .Y(_11575_));
 AO22x1_ASAP7_75t_R _31270_ (.A1(net12),
    .A2(_11540_),
    .B1(_09532_),
    .B2(_11542_),
    .Y(_11576_));
 AO21x1_ASAP7_75t_R _31271_ (.A1(_11575_),
    .A2(_11543_),
    .B(_11576_),
    .Y(_04137_));
 INVx1_ASAP7_75t_R _31272_ (.A(_00135_),
    .Y(_11577_));
 AO22x1_ASAP7_75t_R _31273_ (.A1(net13),
    .A2(_11540_),
    .B1(_09539_),
    .B2(_11542_),
    .Y(_11578_));
 AO21x1_ASAP7_75t_R _31274_ (.A1(_11577_),
    .A2(_11543_),
    .B(_11578_),
    .Y(_04138_));
 INVx1_ASAP7_75t_R _31275_ (.A(_00138_),
    .Y(_11579_));
 AO22x1_ASAP7_75t_R _31276_ (.A1(net14),
    .A2(_11540_),
    .B1(_09545_),
    .B2(_11542_),
    .Y(_11580_));
 AO21x1_ASAP7_75t_R _31277_ (.A1(_11579_),
    .A2(_11543_),
    .B(_11580_),
    .Y(_04139_));
 INVx1_ASAP7_75t_R _31278_ (.A(_00141_),
    .Y(_11581_));
 AO22x1_ASAP7_75t_R _31279_ (.A1(net15),
    .A2(_11540_),
    .B1(_11192_),
    .B2(_11542_),
    .Y(_11582_));
 AO21x1_ASAP7_75t_R _31280_ (.A1(_11581_),
    .A2(_11543_),
    .B(_11582_),
    .Y(_04140_));
 INVx1_ASAP7_75t_R _31281_ (.A(_00144_),
    .Y(_11583_));
 AO22x1_ASAP7_75t_R _31282_ (.A1(net16),
    .A2(_11540_),
    .B1(_09565_),
    .B2(_11542_),
    .Y(_11584_));
 AO21x1_ASAP7_75t_R _31283_ (.A1(_11583_),
    .A2(_11543_),
    .B(_11584_),
    .Y(_04141_));
 INVx1_ASAP7_75t_R _31284_ (.A(_00147_),
    .Y(_11585_));
 AO22x1_ASAP7_75t_R _31285_ (.A1(net17),
    .A2(_11540_),
    .B1(_09572_),
    .B2(_11542_),
    .Y(_11586_));
 AO21x1_ASAP7_75t_R _31286_ (.A1(_11585_),
    .A2(_11543_),
    .B(_11586_),
    .Y(_04142_));
 INVx1_ASAP7_75t_R _31287_ (.A(_00150_),
    .Y(_11587_));
 AO22x1_ASAP7_75t_R _31288_ (.A1(net18),
    .A2(_11540_),
    .B1(_09578_),
    .B2(_11542_),
    .Y(_11588_));
 AO21x1_ASAP7_75t_R _31289_ (.A1(_11587_),
    .A2(_11543_),
    .B(_11588_),
    .Y(_04143_));
 INVx1_ASAP7_75t_R _31290_ (.A(_00153_),
    .Y(_11589_));
 AO22x1_ASAP7_75t_R _31291_ (.A1(net19),
    .A2(_11540_),
    .B1(_09585_),
    .B2(_11542_),
    .Y(_11590_));
 AO21x1_ASAP7_75t_R _31292_ (.A1(_11589_),
    .A2(_11543_),
    .B(_11590_),
    .Y(_04144_));
 INVx1_ASAP7_75t_R _31293_ (.A(_00156_),
    .Y(_11591_));
 AO22x1_ASAP7_75t_R _31294_ (.A1(net20),
    .A2(_11540_),
    .B1(_09591_),
    .B2(_11542_),
    .Y(_11592_));
 AO21x1_ASAP7_75t_R _31295_ (.A1(_11591_),
    .A2(_11543_),
    .B(_11592_),
    .Y(_04145_));
 INVx1_ASAP7_75t_R _31296_ (.A(_00159_),
    .Y(_11593_));
 AO22x1_ASAP7_75t_R _31297_ (.A1(net21),
    .A2(_11540_),
    .B1(_09598_),
    .B2(_11542_),
    .Y(_11594_));
 AO21x1_ASAP7_75t_R _31298_ (.A1(_11593_),
    .A2(_11543_),
    .B(_11594_),
    .Y(_04146_));
 INVx1_ASAP7_75t_R _31299_ (.A(_00161_),
    .Y(_11595_));
 AO22x1_ASAP7_75t_R _31300_ (.A1(net22),
    .A2(_11540_),
    .B1(_09605_),
    .B2(_11542_),
    .Y(_11596_));
 AO21x1_ASAP7_75t_R _31301_ (.A1(_11595_),
    .A2(_11543_),
    .B(_11596_),
    .Y(_04147_));
 AND3x1_ASAP7_75t_R _31302_ (.A(_14083_),
    .B(_07504_),
    .C(_09351_),
    .Y(_11597_));
 NAND2x1_ASAP7_75t_R _31303_ (.A(_06884_),
    .B(_11597_),
    .Y(_11598_));
 AND3x2_ASAP7_75t_R _31304_ (.A(_09364_),
    .B(_07504_),
    .C(_09351_),
    .Y(_11599_));
 AND3x1_ASAP7_75t_R _31305_ (.A(_07513_),
    .B(_10975_),
    .C(_11599_),
    .Y(_11600_));
 AOI21x1_ASAP7_75t_R _31306_ (.A1(_11095_),
    .A2(_11598_),
    .B(_11600_),
    .Y(_11601_));
 TAPCELL_ASAP7_75t_R PHY_191 ();
 AO21x2_ASAP7_75t_R _31308_ (.A1(_11095_),
    .A2(_11598_),
    .B(_11600_),
    .Y(_11603_));
 OA211x2_ASAP7_75t_R _31309_ (.A1(_02424_),
    .A2(_11112_),
    .B(_11100_),
    .C(_11603_),
    .Y(_11604_));
 AOI21x1_ASAP7_75t_R _31310_ (.A1(_02066_),
    .A2(net254),
    .B(_11604_),
    .Y(_04148_));
 TAPCELL_ASAP7_75t_R PHY_190 ();
 TAPCELL_ASAP7_75t_R PHY_189 ();
 INVx1_ASAP7_75t_R _31313_ (.A(_02423_),
    .Y(_11607_));
 AO32x1_ASAP7_75t_R _31314_ (.A1(_05991_),
    .A2(_11607_),
    .A3(_11108_),
    .B1(_11112_),
    .B2(_11107_),
    .Y(_11608_));
 TAPCELL_ASAP7_75t_R PHY_188 ();
 AO21x1_ASAP7_75t_R _31316_ (.A1(_02423_),
    .A2(_11108_),
    .B(net254),
    .Y(_11610_));
 AOI22x1_ASAP7_75t_R _31317_ (.A1(_11603_),
    .A2(_11608_),
    .B1(_11610_),
    .B2(_02065_),
    .Y(_04149_));
 OA211x2_ASAP7_75t_R _31318_ (.A1(_02426_),
    .A2(_11112_),
    .B(_11115_),
    .C(_11603_),
    .Y(_11611_));
 AOI21x1_ASAP7_75t_R _31319_ (.A1(_02064_),
    .A2(net254),
    .B(_11611_),
    .Y(_04150_));
 OR3x1_ASAP7_75t_R _31320_ (.A(_02063_),
    .B(_02425_),
    .C(_11112_),
    .Y(_11612_));
 OAI21x1_ASAP7_75t_R _31321_ (.A1(_09397_),
    .A2(_11108_),
    .B(_11612_),
    .Y(_11613_));
 AO21x1_ASAP7_75t_R _31322_ (.A1(_02425_),
    .A2(_11108_),
    .B(net254),
    .Y(_11614_));
 AOI22x1_ASAP7_75t_R _31323_ (.A1(_11603_),
    .A2(_11613_),
    .B1(_11614_),
    .B2(_02063_),
    .Y(_04151_));
 OA211x2_ASAP7_75t_R _31324_ (.A1(_02428_),
    .A2(_11112_),
    .B(_11125_),
    .C(_11603_),
    .Y(_11615_));
 AOI21x1_ASAP7_75t_R _31325_ (.A1(_02062_),
    .A2(_11601_),
    .B(_11615_),
    .Y(_04152_));
 INVx1_ASAP7_75t_R _31326_ (.A(_02427_),
    .Y(_11616_));
 TAPCELL_ASAP7_75t_R PHY_187 ();
 AO32x1_ASAP7_75t_R _31328_ (.A1(_05993_),
    .A2(_11616_),
    .A3(_11099_),
    .B1(_11174_),
    .B2(_11010_),
    .Y(_11618_));
 TAPCELL_ASAP7_75t_R PHY_186 ();
 AO21x1_ASAP7_75t_R _31330_ (.A1(_02427_),
    .A2(_11099_),
    .B(_11601_),
    .Y(_11620_));
 AOI22x1_ASAP7_75t_R _31331_ (.A1(_11603_),
    .A2(_11618_),
    .B1(_11620_),
    .B2(_02061_),
    .Y(_04153_));
 AO21x1_ASAP7_75t_R _31332_ (.A1(_02430_),
    .A2(_11099_),
    .B(_11133_),
    .Y(_11621_));
 TAPCELL_ASAP7_75t_R PHY_185 ();
 AND2x2_ASAP7_75t_R _31334_ (.A(_02060_),
    .B(_11601_),
    .Y(_11623_));
 AOI21x1_ASAP7_75t_R _31335_ (.A1(_11603_),
    .A2(_11621_),
    .B(_11623_),
    .Y(_04154_));
 AO21x1_ASAP7_75t_R _31336_ (.A1(_02429_),
    .A2(_11099_),
    .B(_11601_),
    .Y(_11624_));
 INVx1_ASAP7_75t_R _31337_ (.A(_02059_),
    .Y(_11625_));
 INVx1_ASAP7_75t_R _31338_ (.A(_02429_),
    .Y(_11626_));
 AO32x1_ASAP7_75t_R _31339_ (.A1(_11625_),
    .A2(_11626_),
    .A3(_11099_),
    .B1(_11174_),
    .B2(_11236_),
    .Y(_11627_));
 AOI22x1_ASAP7_75t_R _31340_ (.A1(_02059_),
    .A2(_11624_),
    .B1(_11627_),
    .B2(_11603_),
    .Y(_04155_));
 AO21x1_ASAP7_75t_R _31341_ (.A1(_02432_),
    .A2(_11099_),
    .B(_11140_),
    .Y(_11628_));
 AND2x2_ASAP7_75t_R _31342_ (.A(_02058_),
    .B(_11601_),
    .Y(_11629_));
 AOI21x1_ASAP7_75t_R _31343_ (.A1(_11603_),
    .A2(_11628_),
    .B(_11629_),
    .Y(_04156_));
 AO21x1_ASAP7_75t_R _31344_ (.A1(_02431_),
    .A2(_11099_),
    .B(_11601_),
    .Y(_11630_));
 OR3x1_ASAP7_75t_R _31345_ (.A(_02057_),
    .B(_02431_),
    .C(_11112_),
    .Y(_11631_));
 OA21x2_ASAP7_75t_R _31346_ (.A1(_09445_),
    .A2(_11108_),
    .B(_11631_),
    .Y(_11632_));
 NOR2x1_ASAP7_75t_R _31347_ (.A(_11601_),
    .B(_11632_),
    .Y(_11633_));
 AOI21x1_ASAP7_75t_R _31348_ (.A1(_02057_),
    .A2(_11630_),
    .B(_11633_),
    .Y(_04157_));
 AO21x1_ASAP7_75t_R _31349_ (.A1(_02434_),
    .A2(_11099_),
    .B(_11146_),
    .Y(_11634_));
 AND2x2_ASAP7_75t_R _31350_ (.A(_02056_),
    .B(_11601_),
    .Y(_11635_));
 AOI21x1_ASAP7_75t_R _31351_ (.A1(_11603_),
    .A2(_11634_),
    .B(_11635_),
    .Y(_04158_));
 AO21x1_ASAP7_75t_R _31352_ (.A1(_02433_),
    .A2(_11099_),
    .B(_11601_),
    .Y(_11636_));
 OR3x1_ASAP7_75t_R _31353_ (.A(_02055_),
    .B(_02433_),
    .C(_11112_),
    .Y(_11637_));
 OA21x2_ASAP7_75t_R _31354_ (.A1(_09458_),
    .A2(_11108_),
    .B(_11637_),
    .Y(_11638_));
 NOR2x1_ASAP7_75t_R _31355_ (.A(_11601_),
    .B(_11638_),
    .Y(_11639_));
 AOI21x1_ASAP7_75t_R _31356_ (.A1(_02055_),
    .A2(_11636_),
    .B(_11639_),
    .Y(_04159_));
 AO21x1_ASAP7_75t_R _31357_ (.A1(_02436_),
    .A2(_11099_),
    .B(_11152_),
    .Y(_11640_));
 AND2x2_ASAP7_75t_R _31358_ (.A(_02054_),
    .B(_11601_),
    .Y(_11641_));
 AOI21x1_ASAP7_75t_R _31359_ (.A1(_11603_),
    .A2(_11640_),
    .B(_11641_),
    .Y(_04160_));
 INVx1_ASAP7_75t_R _31360_ (.A(_02435_),
    .Y(_11642_));
 INVx1_ASAP7_75t_R _31361_ (.A(_09473_),
    .Y(_11643_));
 AO32x1_ASAP7_75t_R _31362_ (.A1(_05997_),
    .A2(_11642_),
    .A3(_11099_),
    .B1(_11174_),
    .B2(_11643_),
    .Y(_11644_));
 AO21x1_ASAP7_75t_R _31363_ (.A1(_02435_),
    .A2(_11099_),
    .B(_11601_),
    .Y(_11645_));
 AOI22x1_ASAP7_75t_R _31364_ (.A1(_11603_),
    .A2(_11644_),
    .B1(_11645_),
    .B2(_02053_),
    .Y(_04161_));
 AO21x1_ASAP7_75t_R _31365_ (.A1(_02438_),
    .A2(_11099_),
    .B(_11159_),
    .Y(_11646_));
 AND2x2_ASAP7_75t_R _31366_ (.A(_02052_),
    .B(_11601_),
    .Y(_11647_));
 AOI21x1_ASAP7_75t_R _31367_ (.A1(_11603_),
    .A2(_11646_),
    .B(_11647_),
    .Y(_04162_));
 INVx1_ASAP7_75t_R _31368_ (.A(_02051_),
    .Y(_11648_));
 AO21x1_ASAP7_75t_R _31369_ (.A1(_02437_),
    .A2(_11099_),
    .B(_11601_),
    .Y(_11649_));
 INVx1_ASAP7_75t_R _31370_ (.A(_02437_),
    .Y(_11650_));
 AO32x1_ASAP7_75t_R _31371_ (.A1(_02051_),
    .A2(_11650_),
    .A3(_11099_),
    .B1(_11174_),
    .B2(_09488_),
    .Y(_11651_));
 AO22x1_ASAP7_75t_R _31372_ (.A1(_11648_),
    .A2(_11649_),
    .B1(_11651_),
    .B2(_11603_),
    .Y(_04163_));
 OA211x2_ASAP7_75t_R _31373_ (.A1(_02440_),
    .A2(_11112_),
    .B(_11165_),
    .C(_11603_),
    .Y(_11652_));
 AOI21x1_ASAP7_75t_R _31374_ (.A1(_02050_),
    .A2(_11601_),
    .B(_11652_),
    .Y(_04164_));
 INVx1_ASAP7_75t_R _31375_ (.A(_02049_),
    .Y(_11653_));
 AO21x1_ASAP7_75t_R _31376_ (.A1(_02439_),
    .A2(_11099_),
    .B(_11601_),
    .Y(_11654_));
 INVx1_ASAP7_75t_R _31377_ (.A(_02439_),
    .Y(_11655_));
 AO32x1_ASAP7_75t_R _31378_ (.A1(_02049_),
    .A2(_11655_),
    .A3(_11099_),
    .B1(_11174_),
    .B2(_09503_),
    .Y(_11656_));
 AND2x2_ASAP7_75t_R _31379_ (.A(_11603_),
    .B(_11656_),
    .Y(_11657_));
 AO21x1_ASAP7_75t_R _31380_ (.A1(_11653_),
    .A2(_11654_),
    .B(_11657_),
    .Y(_04165_));
 OA211x2_ASAP7_75t_R _31381_ (.A1(_02442_),
    .A2(_11112_),
    .B(_11170_),
    .C(_11603_),
    .Y(_11658_));
 AOI21x1_ASAP7_75t_R _31382_ (.A1(_02048_),
    .A2(net254),
    .B(_11658_),
    .Y(_04166_));
 INVx1_ASAP7_75t_R _31383_ (.A(_02047_),
    .Y(_11659_));
 AO21x1_ASAP7_75t_R _31384_ (.A1(_02441_),
    .A2(_11099_),
    .B(net254),
    .Y(_11660_));
 INVx1_ASAP7_75t_R _31385_ (.A(_02441_),
    .Y(_11661_));
 AO32x1_ASAP7_75t_R _31386_ (.A1(_02047_),
    .A2(_11661_),
    .A3(_11099_),
    .B1(_11174_),
    .B2(_09519_),
    .Y(_11662_));
 AO22x1_ASAP7_75t_R _31387_ (.A1(_11659_),
    .A2(_11660_),
    .B1(_11662_),
    .B2(_11603_),
    .Y(_04167_));
 AO21x1_ASAP7_75t_R _31388_ (.A1(_02444_),
    .A2(_11099_),
    .B(_11179_),
    .Y(_11663_));
 AND2x2_ASAP7_75t_R _31389_ (.A(_02046_),
    .B(net254),
    .Y(_11664_));
 AOI21x1_ASAP7_75t_R _31390_ (.A1(_11603_),
    .A2(_11663_),
    .B(_11664_),
    .Y(_04168_));
 INVx1_ASAP7_75t_R _31391_ (.A(_02045_),
    .Y(_11665_));
 AO21x1_ASAP7_75t_R _31392_ (.A1(_02443_),
    .A2(_11099_),
    .B(net254),
    .Y(_11666_));
 INVx1_ASAP7_75t_R _31393_ (.A(_02443_),
    .Y(_11667_));
 AO32x1_ASAP7_75t_R _31394_ (.A1(_02045_),
    .A2(_11667_),
    .A3(_11099_),
    .B1(_11174_),
    .B2(_09532_),
    .Y(_11668_));
 AO22x1_ASAP7_75t_R _31395_ (.A1(_11665_),
    .A2(_11666_),
    .B1(_11668_),
    .B2(_11603_),
    .Y(_04169_));
 AOI21x1_ASAP7_75t_R _31396_ (.A1(_02446_),
    .A2(_11099_),
    .B(_11186_),
    .Y(_11669_));
 NAND2x1_ASAP7_75t_R _31397_ (.A(_02044_),
    .B(net254),
    .Y(_11670_));
 OA21x2_ASAP7_75t_R _31398_ (.A1(net254),
    .A2(_11669_),
    .B(_11670_),
    .Y(_04170_));
 INVx1_ASAP7_75t_R _31399_ (.A(_02043_),
    .Y(_11671_));
 INVx1_ASAP7_75t_R _31400_ (.A(_02445_),
    .Y(_11672_));
 INVx2_ASAP7_75t_R _31401_ (.A(_09545_),
    .Y(_11673_));
 AO32x1_ASAP7_75t_R _31402_ (.A1(_11671_),
    .A2(_11672_),
    .A3(_11099_),
    .B1(_11174_),
    .B2(_11673_),
    .Y(_11674_));
 AO21x1_ASAP7_75t_R _31403_ (.A1(_02445_),
    .A2(_11099_),
    .B(net254),
    .Y(_11675_));
 AOI22x1_ASAP7_75t_R _31404_ (.A1(_11603_),
    .A2(_11674_),
    .B1(_11675_),
    .B2(_02043_),
    .Y(_04171_));
 INVx1_ASAP7_75t_R _31405_ (.A(_02448_),
    .Y(_11676_));
 AO221x1_ASAP7_75t_R _31406_ (.A1(_11192_),
    .A2(_11174_),
    .B1(_11099_),
    .B2(_11676_),
    .C(net254),
    .Y(_11677_));
 OA21x2_ASAP7_75t_R _31407_ (.A1(\cs_registers_i.mhpmcounter[2][56] ),
    .A2(_11603_),
    .B(_11677_),
    .Y(_04172_));
 INVx1_ASAP7_75t_R _31408_ (.A(_02041_),
    .Y(_11678_));
 AO21x1_ASAP7_75t_R _31409_ (.A1(_02447_),
    .A2(_11099_),
    .B(net254),
    .Y(_11679_));
 INVx1_ASAP7_75t_R _31410_ (.A(_02447_),
    .Y(_11680_));
 AO32x1_ASAP7_75t_R _31411_ (.A1(_02041_),
    .A2(_11680_),
    .A3(_11099_),
    .B1(_11174_),
    .B2(_09565_),
    .Y(_11681_));
 AO22x1_ASAP7_75t_R _31412_ (.A1(_11678_),
    .A2(_11679_),
    .B1(_11681_),
    .B2(_11603_),
    .Y(_04173_));
 AO21x1_ASAP7_75t_R _31413_ (.A1(_02450_),
    .A2(_11099_),
    .B(_11198_),
    .Y(_11682_));
 AND2x2_ASAP7_75t_R _31414_ (.A(_02040_),
    .B(net254),
    .Y(_11683_));
 AOI21x1_ASAP7_75t_R _31415_ (.A1(_11603_),
    .A2(_11682_),
    .B(_11683_),
    .Y(_04174_));
 INVx1_ASAP7_75t_R _31416_ (.A(_02039_),
    .Y(_11684_));
 AO21x1_ASAP7_75t_R _31417_ (.A1(_02449_),
    .A2(_11099_),
    .B(net254),
    .Y(_11685_));
 INVx1_ASAP7_75t_R _31418_ (.A(_02449_),
    .Y(_11686_));
 AO32x1_ASAP7_75t_R _31419_ (.A1(_02039_),
    .A2(_11686_),
    .A3(_11099_),
    .B1(_11174_),
    .B2(_09578_),
    .Y(_11687_));
 AND2x2_ASAP7_75t_R _31420_ (.A(_11603_),
    .B(_11687_),
    .Y(_11688_));
 AO21x1_ASAP7_75t_R _31421_ (.A1(_11684_),
    .A2(_11685_),
    .B(_11688_),
    .Y(_04175_));
 OA211x2_ASAP7_75t_R _31422_ (.A1(_02452_),
    .A2(_11112_),
    .B(_11206_),
    .C(_11603_),
    .Y(_11689_));
 AOI21x1_ASAP7_75t_R _31423_ (.A1(_02038_),
    .A2(net254),
    .B(_11689_),
    .Y(_04176_));
 AO21x1_ASAP7_75t_R _31424_ (.A1(_02451_),
    .A2(_11099_),
    .B(net254),
    .Y(_11690_));
 OR3x1_ASAP7_75t_R _31425_ (.A(_02037_),
    .B(_02451_),
    .C(_11112_),
    .Y(_11691_));
 OA21x2_ASAP7_75t_R _31426_ (.A1(_09591_),
    .A2(_11108_),
    .B(_11691_),
    .Y(_11692_));
 NOR2x1_ASAP7_75t_R _31427_ (.A(net254),
    .B(_11692_),
    .Y(_11693_));
 AOI21x1_ASAP7_75t_R _31428_ (.A1(_02037_),
    .A2(_11690_),
    .B(_11693_),
    .Y(_04177_));
 OA211x2_ASAP7_75t_R _31429_ (.A1(_02454_),
    .A2(_11112_),
    .B(_11213_),
    .C(_11603_),
    .Y(_11694_));
 AOI21x1_ASAP7_75t_R _31430_ (.A1(_02036_),
    .A2(net254),
    .B(_11694_),
    .Y(_04178_));
 INVx1_ASAP7_75t_R _31431_ (.A(_02035_),
    .Y(_11695_));
 INVx1_ASAP7_75t_R _31432_ (.A(_02453_),
    .Y(_11696_));
 AO32x1_ASAP7_75t_R _31433_ (.A1(_11695_),
    .A2(_11696_),
    .A3(_11099_),
    .B1(_11174_),
    .B2(_11215_),
    .Y(_11697_));
 AO21x1_ASAP7_75t_R _31434_ (.A1(_02453_),
    .A2(_11108_),
    .B(net254),
    .Y(_11698_));
 AOI22x1_ASAP7_75t_R _31435_ (.A1(_11603_),
    .A2(_11697_),
    .B1(_11698_),
    .B2(_02035_),
    .Y(_04179_));
 NAND2x2_ASAP7_75t_R _31436_ (.A(_05582_),
    .B(_11497_),
    .Y(_11699_));
 TAPCELL_ASAP7_75t_R PHY_184 ();
 AO21x1_ASAP7_75t_R _31438_ (.A1(_05582_),
    .A2(_11497_),
    .B(_06870_),
    .Y(_11701_));
 OA21x2_ASAP7_75t_R _31439_ (.A1(_09390_),
    .A2(_11699_),
    .B(_11701_),
    .Y(_04180_));
 NAND2x1_ASAP7_75t_R _31440_ (.A(_02033_),
    .B(_11699_),
    .Y(_11702_));
 OA21x2_ASAP7_75t_R _31441_ (.A1(_09458_),
    .A2(_11699_),
    .B(_11702_),
    .Y(_04181_));
 NAND2x1_ASAP7_75t_R _31442_ (.A(_02032_),
    .B(_11699_),
    .Y(_11703_));
 OA21x2_ASAP7_75t_R _31443_ (.A1(_09465_),
    .A2(_11699_),
    .B(_11703_),
    .Y(_04182_));
 NAND2x1_ASAP7_75t_R _31444_ (.A(_02031_),
    .B(_11699_),
    .Y(_11704_));
 OA21x2_ASAP7_75t_R _31445_ (.A1(_09473_),
    .A2(_11699_),
    .B(_11704_),
    .Y(_04183_));
 NAND2x1_ASAP7_75t_R _31446_ (.A(_02030_),
    .B(_11699_),
    .Y(_11705_));
 OA21x2_ASAP7_75t_R _31447_ (.A1(_09488_),
    .A2(_11699_),
    .B(_11705_),
    .Y(_04184_));
 INVx1_ASAP7_75t_R _31448_ (.A(_05723_),
    .Y(_11706_));
 TAPCELL_ASAP7_75t_R PHY_183 ();
 AO221x2_ASAP7_75t_R _31450_ (.A1(_01719_),
    .A2(_01725_),
    .B1(_11706_),
    .B2(_13227_),
    .C(_06174_),
    .Y(_11708_));
 TAPCELL_ASAP7_75t_R PHY_182 ();
 TAPCELL_ASAP7_75t_R PHY_181 ();
 TAPCELL_ASAP7_75t_R PHY_180 ();
 TAPCELL_ASAP7_75t_R PHY_179 ();
 TAPCELL_ASAP7_75t_R PHY_178 ();
 AND2x2_ASAP7_75t_R _31456_ (.A(_00385_),
    .B(_01746_),
    .Y(_11714_));
 AO21x1_ASAP7_75t_R _31457_ (.A1(_05549_),
    .A2(_01723_),
    .B(_11714_),
    .Y(_11715_));
 OR4x1_ASAP7_75t_R _31458_ (.A(_01312_),
    .B(_06167_),
    .C(_06172_),
    .D(_11715_),
    .Y(_11716_));
 OAI21x1_ASAP7_75t_R _31459_ (.A1(_01641_),
    .A2(_11708_),
    .B(_11716_),
    .Y(_11717_));
 AND2x2_ASAP7_75t_R _31460_ (.A(_01311_),
    .B(_05527_),
    .Y(_11718_));
 INVx2_ASAP7_75t_R _31461_ (.A(_07523_),
    .Y(_11719_));
 AND3x4_ASAP7_75t_R _31462_ (.A(_07522_),
    .B(_11719_),
    .C(_09365_),
    .Y(_11720_));
 TAPCELL_ASAP7_75t_R PHY_177 ();
 TAPCELL_ASAP7_75t_R PHY_176 ();
 NOR3x1_ASAP7_75t_R _31465_ (.A(_02029_),
    .B(_11242_),
    .C(_11720_),
    .Y(_11723_));
 AO221x1_ASAP7_75t_R _31466_ (.A1(_11717_),
    .A2(_11718_),
    .B1(_11720_),
    .B2(_10974_),
    .C(_11723_),
    .Y(_04185_));
 AND3x4_ASAP7_75t_R _31467_ (.A(_05630_),
    .B(_07144_),
    .C(_09353_),
    .Y(_11724_));
 TAPCELL_ASAP7_75t_R PHY_175 ();
 NOR2x2_ASAP7_75t_R _31469_ (.A(_11242_),
    .B(_11724_),
    .Y(_11726_));
 TAPCELL_ASAP7_75t_R PHY_174 ();
 INVx1_ASAP7_75t_R _31471_ (.A(_02028_),
    .Y(_11728_));
 TAPCELL_ASAP7_75t_R PHY_173 ();
 TAPCELL_ASAP7_75t_R PHY_172 ();
 TAPCELL_ASAP7_75t_R PHY_171 ();
 TAPCELL_ASAP7_75t_R PHY_170 ();
 XOR2x1_ASAP7_75t_R _31476_ (.A(net421),
    .Y(_11733_),
    .B(_01720_));
 TAPCELL_ASAP7_75t_R PHY_169 ();
 AND2x2_ASAP7_75t_R _31478_ (.A(_00385_),
    .B(_00163_),
    .Y(_11735_));
 AO21x1_ASAP7_75t_R _31479_ (.A1(_05549_),
    .A2(_00164_),
    .B(_11735_),
    .Y(_11736_));
 OA222x2_ASAP7_75t_R _31480_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11708_),
    .B2(_01640_),
    .C1(_11736_),
    .C2(_01312_),
    .Y(_11737_));
 INVx1_ASAP7_75t_R _31481_ (.A(_11737_),
    .Y(_11738_));
 AND2x6_ASAP7_75t_R _31482_ (.A(_06340_),
    .B(_11242_),
    .Y(_11739_));
 TAPCELL_ASAP7_75t_R PHY_168 ();
 OA211x2_ASAP7_75t_R _31484_ (.A1(_06165_),
    .A2(_11733_),
    .B(_11738_),
    .C(_11739_),
    .Y(_11741_));
 AO221x1_ASAP7_75t_R _31485_ (.A1(_09363_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11728_),
    .C(_11741_),
    .Y(_04186_));
 TAPCELL_ASAP7_75t_R PHY_167 ();
 TAPCELL_ASAP7_75t_R PHY_166 ();
 TAPCELL_ASAP7_75t_R PHY_165 ();
 NOR2x1_ASAP7_75t_R _31489_ (.A(_00167_),
    .B(net421),
    .Y(_11745_));
 AO21x1_ASAP7_75t_R _31490_ (.A1(\cs_registers_i.pc_id_i[2] ),
    .A2(net421),
    .B(_11745_),
    .Y(_11746_));
 TAPCELL_ASAP7_75t_R PHY_164 ();
 AND2x2_ASAP7_75t_R _31492_ (.A(_00385_),
    .B(_00165_),
    .Y(_11748_));
 AO21x1_ASAP7_75t_R _31493_ (.A1(_05549_),
    .A2(_00166_),
    .B(_11748_),
    .Y(_11749_));
 OA222x2_ASAP7_75t_R _31494_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11708_),
    .B2(_01639_),
    .C1(_11749_),
    .C2(_01312_),
    .Y(_11750_));
 INVx1_ASAP7_75t_R _31495_ (.A(_11750_),
    .Y(_11751_));
 OA211x2_ASAP7_75t_R _31496_ (.A1(_06165_),
    .A2(_11746_),
    .B(_11751_),
    .C(_11739_),
    .Y(_11752_));
 AO221x1_ASAP7_75t_R _31497_ (.A1(_09390_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_07370_),
    .C(_11752_),
    .Y(_04187_));
 INVx1_ASAP7_75t_R _31498_ (.A(_02026_),
    .Y(_11753_));
 TAPCELL_ASAP7_75t_R PHY_163 ();
 TAPCELL_ASAP7_75t_R PHY_162 ();
 NOR2x1_ASAP7_75t_R _31501_ (.A(net421),
    .B(_00171_),
    .Y(_11756_));
 AO21x1_ASAP7_75t_R _31502_ (.A1(net421),
    .A2(\cs_registers_i.pc_id_i[3] ),
    .B(_11756_),
    .Y(_11757_));
 AND2x2_ASAP7_75t_R _31503_ (.A(_00385_),
    .B(_00168_),
    .Y(_11758_));
 AO21x1_ASAP7_75t_R _31504_ (.A1(_05549_),
    .A2(_00169_),
    .B(_11758_),
    .Y(_11759_));
 OA222x2_ASAP7_75t_R _31505_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11708_),
    .B2(_01638_),
    .C1(_11759_),
    .C2(_01312_),
    .Y(_11760_));
 INVx1_ASAP7_75t_R _31506_ (.A(_11760_),
    .Y(_11761_));
 OA211x2_ASAP7_75t_R _31507_ (.A1(_06165_),
    .A2(_11757_),
    .B(_11761_),
    .C(_11739_),
    .Y(_11762_));
 AO221x1_ASAP7_75t_R _31508_ (.A1(_09397_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11753_),
    .C(_11762_),
    .Y(_04188_));
 INVx1_ASAP7_75t_R _31509_ (.A(_02025_),
    .Y(_11763_));
 TAPCELL_ASAP7_75t_R PHY_161 ();
 TAPCELL_ASAP7_75t_R PHY_160 ();
 AND2x2_ASAP7_75t_R _31512_ (.A(_00385_),
    .B(_00172_),
    .Y(_11766_));
 AO21x1_ASAP7_75t_R _31513_ (.A1(_05549_),
    .A2(_00173_),
    .B(_11766_),
    .Y(_11767_));
 OAI22x1_ASAP7_75t_R _31514_ (.A1(_01637_),
    .A2(_11708_),
    .B1(_11767_),
    .B2(_01312_),
    .Y(_11768_));
 OAI21x1_ASAP7_75t_R _31515_ (.A1(net421),
    .A2(_02520_),
    .B(_00174_),
    .Y(_11769_));
 OR3x1_ASAP7_75t_R _31516_ (.A(net421),
    .B(_00174_),
    .C(_02520_),
    .Y(_11770_));
 TAPCELL_ASAP7_75t_R PHY_159 ();
 AO21x1_ASAP7_75t_R _31518_ (.A1(_11769_),
    .A2(_11770_),
    .B(_06165_),
    .Y(_11772_));
 OA211x2_ASAP7_75t_R _31519_ (.A1(_06172_),
    .A2(_11768_),
    .B(_11772_),
    .C(_11739_),
    .Y(_11773_));
 AO221x1_ASAP7_75t_R _31520_ (.A1(_09408_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11763_),
    .C(_11773_),
    .Y(_04189_));
 INVx1_ASAP7_75t_R _31521_ (.A(_02024_),
    .Y(_11774_));
 NOR2x1_ASAP7_75t_R _31522_ (.A(net421),
    .B(_00178_),
    .Y(_11775_));
 AO21x1_ASAP7_75t_R _31523_ (.A1(net421),
    .A2(\cs_registers_i.pc_id_i[5] ),
    .B(_11775_),
    .Y(_11776_));
 AND2x2_ASAP7_75t_R _31524_ (.A(_00385_),
    .B(_00175_),
    .Y(_11777_));
 AO21x1_ASAP7_75t_R _31525_ (.A1(_05549_),
    .A2(_00176_),
    .B(_11777_),
    .Y(_11778_));
 OA222x2_ASAP7_75t_R _31526_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11708_),
    .B2(_01636_),
    .C1(_11778_),
    .C2(_01312_),
    .Y(_11779_));
 INVx1_ASAP7_75t_R _31527_ (.A(_11779_),
    .Y(_11780_));
 OA211x2_ASAP7_75t_R _31528_ (.A1(_06165_),
    .A2(_11776_),
    .B(_11780_),
    .C(_11739_),
    .Y(_11781_));
 AO221x1_ASAP7_75t_R _31529_ (.A1(_09417_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11774_),
    .C(_11781_),
    .Y(_04190_));
 INVx1_ASAP7_75t_R _31530_ (.A(_02023_),
    .Y(_11782_));
 NAND2x1_ASAP7_75t_R _31531_ (.A(_00278_),
    .B(_00385_),
    .Y(_11783_));
 NAND2x1_ASAP7_75t_R _31532_ (.A(_05549_),
    .B(_00179_),
    .Y(_11784_));
 INVx3_ASAP7_75t_R _31533_ (.A(_11708_),
    .Y(_11785_));
 AO32x1_ASAP7_75t_R _31534_ (.A1(_06174_),
    .A2(_11783_),
    .A3(_11784_),
    .B1(_14885_),
    .B2(_11785_),
    .Y(_11786_));
 OAI21x1_ASAP7_75t_R _31535_ (.A1(net421),
    .A2(_02521_),
    .B(_00180_),
    .Y(_11787_));
 OR3x1_ASAP7_75t_R _31536_ (.A(net421),
    .B(_00180_),
    .C(_02521_),
    .Y(_11788_));
 AO21x1_ASAP7_75t_R _31537_ (.A1(_11787_),
    .A2(_11788_),
    .B(_06165_),
    .Y(_11789_));
 OA211x2_ASAP7_75t_R _31538_ (.A1(_06172_),
    .A2(_11786_),
    .B(_11789_),
    .C(_11739_),
    .Y(_11790_));
 AO221x1_ASAP7_75t_R _31539_ (.A1(_09426_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11782_),
    .C(_11790_),
    .Y(_04191_));
 INVx1_ASAP7_75t_R _31540_ (.A(_02022_),
    .Y(_11791_));
 NOR2x1_ASAP7_75t_R _31541_ (.A(net421),
    .B(_00183_),
    .Y(_11792_));
 AO21x1_ASAP7_75t_R _31542_ (.A1(net421),
    .A2(\cs_registers_i.pc_id_i[7] ),
    .B(_11792_),
    .Y(_11793_));
 AND2x2_ASAP7_75t_R _31543_ (.A(_00323_),
    .B(_00385_),
    .Y(_11794_));
 AO21x1_ASAP7_75t_R _31544_ (.A1(_05549_),
    .A2(_00181_),
    .B(_11794_),
    .Y(_11795_));
 OA222x2_ASAP7_75t_R _31545_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11708_),
    .B2(_01634_),
    .C1(_11795_),
    .C2(_01312_),
    .Y(_11796_));
 INVx1_ASAP7_75t_R _31546_ (.A(_11796_),
    .Y(_11797_));
 OA211x2_ASAP7_75t_R _31547_ (.A1(_06165_),
    .A2(_11793_),
    .B(_11797_),
    .C(_11739_),
    .Y(_11798_));
 AO221x1_ASAP7_75t_R _31548_ (.A1(_09432_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11791_),
    .C(_11798_),
    .Y(_04192_));
 INVx1_ASAP7_75t_R _31549_ (.A(_02021_),
    .Y(_11799_));
 NAND2x1_ASAP7_75t_R _31550_ (.A(_05549_),
    .B(_00185_),
    .Y(_11800_));
 NAND2x1_ASAP7_75t_R _31551_ (.A(_00385_),
    .B(_00184_),
    .Y(_11801_));
 AO32x1_ASAP7_75t_R _31552_ (.A1(_06174_),
    .A2(_11800_),
    .A3(_11801_),
    .B1(_14995_),
    .B2(_11785_),
    .Y(_11802_));
 OAI21x1_ASAP7_75t_R _31553_ (.A1(net421),
    .A2(_02522_),
    .B(_00186_),
    .Y(_11803_));
 OR3x1_ASAP7_75t_R _31554_ (.A(net421),
    .B(_00186_),
    .C(_02522_),
    .Y(_11804_));
 AO21x1_ASAP7_75t_R _31555_ (.A1(_11803_),
    .A2(_11804_),
    .B(_06165_),
    .Y(_11805_));
 OA211x2_ASAP7_75t_R _31556_ (.A1(_06172_),
    .A2(_11802_),
    .B(_11805_),
    .C(_11739_),
    .Y(_11806_));
 AO221x1_ASAP7_75t_R _31557_ (.A1(_09438_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11799_),
    .C(_11806_),
    .Y(_04193_));
 TAPCELL_ASAP7_75t_R PHY_158 ();
 INVx1_ASAP7_75t_R _31559_ (.A(_02020_),
    .Y(_11808_));
 NOR2x1_ASAP7_75t_R _31560_ (.A(_01722_),
    .B(_00190_),
    .Y(_11809_));
 AO21x1_ASAP7_75t_R _31561_ (.A1(_01722_),
    .A2(\cs_registers_i.pc_id_i[9] ),
    .B(_11809_),
    .Y(_11810_));
 AND2x2_ASAP7_75t_R _31562_ (.A(_00385_),
    .B(_00187_),
    .Y(_11811_));
 AO21x1_ASAP7_75t_R _31563_ (.A1(_05549_),
    .A2(_00188_),
    .B(_11811_),
    .Y(_11812_));
 OA222x2_ASAP7_75t_R _31564_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11708_),
    .B2(_01632_),
    .C1(_11812_),
    .C2(_01312_),
    .Y(_11813_));
 INVx1_ASAP7_75t_R _31565_ (.A(_11813_),
    .Y(_11814_));
 OA211x2_ASAP7_75t_R _31566_ (.A1(_06165_),
    .A2(_11810_),
    .B(_11814_),
    .C(_11739_),
    .Y(_11815_));
 AO221x1_ASAP7_75t_R _31567_ (.A1(_09445_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11808_),
    .C(_11815_),
    .Y(_04194_));
 INVx1_ASAP7_75t_R _31568_ (.A(_02019_),
    .Y(_11816_));
 NAND2x1_ASAP7_75t_R _31569_ (.A(_05549_),
    .B(_00192_),
    .Y(_11817_));
 NAND2x1_ASAP7_75t_R _31570_ (.A(_00385_),
    .B(_00191_),
    .Y(_11818_));
 AO32x1_ASAP7_75t_R _31571_ (.A1(_06174_),
    .A2(_11817_),
    .A3(_11818_),
    .B1(_15109_),
    .B2(_11785_),
    .Y(_11819_));
 OAI21x1_ASAP7_75t_R _31572_ (.A1(_01722_),
    .A2(_02523_),
    .B(_00193_),
    .Y(_11820_));
 TAPCELL_ASAP7_75t_R PHY_157 ();
 OR3x1_ASAP7_75t_R _31574_ (.A(_01722_),
    .B(_00193_),
    .C(_02523_),
    .Y(_11822_));
 AO21x1_ASAP7_75t_R _31575_ (.A1(_11820_),
    .A2(_11822_),
    .B(_06165_),
    .Y(_11823_));
 OA211x2_ASAP7_75t_R _31576_ (.A1(_06172_),
    .A2(_11819_),
    .B(_11823_),
    .C(_11739_),
    .Y(_11824_));
 AO221x1_ASAP7_75t_R _31577_ (.A1(_09452_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11816_),
    .C(_11824_),
    .Y(_04195_));
 INVx1_ASAP7_75t_R _31578_ (.A(_02018_),
    .Y(_11825_));
 NOR2x1_ASAP7_75t_R _31579_ (.A(_01722_),
    .B(_00197_),
    .Y(_11826_));
 AO21x1_ASAP7_75t_R _31580_ (.A1(_01722_),
    .A2(\cs_registers_i.pc_id_i[11] ),
    .B(_11826_),
    .Y(_11827_));
 AND2x2_ASAP7_75t_R _31581_ (.A(_00385_),
    .B(_00194_),
    .Y(_11828_));
 AO21x1_ASAP7_75t_R _31582_ (.A1(_05549_),
    .A2(_00195_),
    .B(_11828_),
    .Y(_11829_));
 OA222x2_ASAP7_75t_R _31583_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11708_),
    .B2(_01630_),
    .C1(_11829_),
    .C2(_01312_),
    .Y(_11830_));
 INVx1_ASAP7_75t_R _31584_ (.A(_11830_),
    .Y(_11831_));
 TAPCELL_ASAP7_75t_R PHY_156 ();
 OA211x2_ASAP7_75t_R _31586_ (.A1(_06165_),
    .A2(_11827_),
    .B(_11831_),
    .C(_11739_),
    .Y(_11833_));
 AO221x1_ASAP7_75t_R _31587_ (.A1(_09458_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11825_),
    .C(_11833_),
    .Y(_04196_));
 TAPCELL_ASAP7_75t_R PHY_155 ();
 INVx1_ASAP7_75t_R _31589_ (.A(_02017_),
    .Y(_11835_));
 AND2x2_ASAP7_75t_R _31590_ (.A(_00281_),
    .B(_00385_),
    .Y(_11836_));
 AO21x1_ASAP7_75t_R _31591_ (.A1(_05549_),
    .A2(_00198_),
    .B(_11836_),
    .Y(_11837_));
 OAI22x1_ASAP7_75t_R _31592_ (.A1(_01629_),
    .A2(_11708_),
    .B1(_11837_),
    .B2(_01312_),
    .Y(_11838_));
 OAI21x1_ASAP7_75t_R _31593_ (.A1(net421),
    .A2(_02524_),
    .B(_00199_),
    .Y(_11839_));
 OR3x1_ASAP7_75t_R _31594_ (.A(net421),
    .B(_00199_),
    .C(_02524_),
    .Y(_11840_));
 AO21x1_ASAP7_75t_R _31595_ (.A1(_11839_),
    .A2(_11840_),
    .B(_06165_),
    .Y(_11841_));
 OA211x2_ASAP7_75t_R _31596_ (.A1(_06172_),
    .A2(_11838_),
    .B(_11841_),
    .C(_11739_),
    .Y(_11842_));
 AO221x1_ASAP7_75t_R _31597_ (.A1(_09465_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11835_),
    .C(_11842_),
    .Y(_04197_));
 INVx1_ASAP7_75t_R _31598_ (.A(_02016_),
    .Y(_11843_));
 NOR2x1_ASAP7_75t_R _31599_ (.A(net421),
    .B(_00202_),
    .Y(_11844_));
 AO21x1_ASAP7_75t_R _31600_ (.A1(net421),
    .A2(\cs_registers_i.pc_id_i[13] ),
    .B(_11844_),
    .Y(_11845_));
 AND2x2_ASAP7_75t_R _31601_ (.A(_00282_),
    .B(_00385_),
    .Y(_11846_));
 AO21x1_ASAP7_75t_R _31602_ (.A1(_05549_),
    .A2(_00200_),
    .B(_11846_),
    .Y(_11847_));
 OA222x2_ASAP7_75t_R _31603_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11708_),
    .B2(_01628_),
    .C1(_11847_),
    .C2(_01312_),
    .Y(_11848_));
 INVx1_ASAP7_75t_R _31604_ (.A(_11848_),
    .Y(_11849_));
 OA211x2_ASAP7_75t_R _31605_ (.A1(_06165_),
    .A2(_11845_),
    .B(_11849_),
    .C(_11739_),
    .Y(_11850_));
 AO221x1_ASAP7_75t_R _31606_ (.A1(_09473_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11843_),
    .C(_11850_),
    .Y(_04198_));
 INVx1_ASAP7_75t_R _31607_ (.A(_02015_),
    .Y(_11851_));
 AND2x2_ASAP7_75t_R _31608_ (.A(_00279_),
    .B(_00385_),
    .Y(_11852_));
 AO21x1_ASAP7_75t_R _31609_ (.A1(_05549_),
    .A2(_00203_),
    .B(_11852_),
    .Y(_11853_));
 OAI22x1_ASAP7_75t_R _31610_ (.A1(_01627_),
    .A2(_11708_),
    .B1(_11853_),
    .B2(_01312_),
    .Y(_11854_));
 OAI21x1_ASAP7_75t_R _31611_ (.A1(net421),
    .A2(_02525_),
    .B(_00204_),
    .Y(_11855_));
 OR3x1_ASAP7_75t_R _31612_ (.A(net421),
    .B(_00204_),
    .C(_02525_),
    .Y(_11856_));
 AO21x1_ASAP7_75t_R _31613_ (.A1(_11855_),
    .A2(_11856_),
    .B(_06165_),
    .Y(_11857_));
 OA211x2_ASAP7_75t_R _31614_ (.A1(_06172_),
    .A2(_11854_),
    .B(_11857_),
    .C(_11739_),
    .Y(_11858_));
 AO221x1_ASAP7_75t_R _31615_ (.A1(_09481_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11851_),
    .C(_11858_),
    .Y(_04199_));
 INVx1_ASAP7_75t_R _31616_ (.A(_02014_),
    .Y(_11859_));
 NOR2x1_ASAP7_75t_R _31617_ (.A(_01722_),
    .B(_00207_),
    .Y(_11860_));
 AO21x1_ASAP7_75t_R _31618_ (.A1(_01722_),
    .A2(\cs_registers_i.pc_id_i[15] ),
    .B(_11860_),
    .Y(_11861_));
 AND2x2_ASAP7_75t_R _31619_ (.A(_00290_),
    .B(_00385_),
    .Y(_11862_));
 AO21x1_ASAP7_75t_R _31620_ (.A1(_05549_),
    .A2(_00205_),
    .B(_11862_),
    .Y(_11863_));
 OA222x2_ASAP7_75t_R _31621_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11708_),
    .B2(_01626_),
    .C1(_11863_),
    .C2(_01312_),
    .Y(_11864_));
 INVx1_ASAP7_75t_R _31622_ (.A(_11864_),
    .Y(_11865_));
 OA211x2_ASAP7_75t_R _31623_ (.A1(_06165_),
    .A2(_11861_),
    .B(_11865_),
    .C(_11739_),
    .Y(_11866_));
 AO221x1_ASAP7_75t_R _31624_ (.A1(_09488_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11859_),
    .C(_11866_),
    .Y(_04200_));
 INVx1_ASAP7_75t_R _31625_ (.A(_02013_),
    .Y(_11867_));
 AO32x1_ASAP7_75t_R _31626_ (.A1(_13433_),
    .A2(_00385_),
    .A3(_06174_),
    .B1(_15733_),
    .B2(_11785_),
    .Y(_11868_));
 OAI21x1_ASAP7_75t_R _31627_ (.A1(_01722_),
    .A2(_02526_),
    .B(_00208_),
    .Y(_11869_));
 OR3x1_ASAP7_75t_R _31628_ (.A(_01722_),
    .B(_00208_),
    .C(_02526_),
    .Y(_11870_));
 AO21x1_ASAP7_75t_R _31629_ (.A1(_11869_),
    .A2(_11870_),
    .B(_06165_),
    .Y(_11871_));
 TAPCELL_ASAP7_75t_R PHY_154 ();
 OA211x2_ASAP7_75t_R _31631_ (.A1(_06172_),
    .A2(_11868_),
    .B(_11871_),
    .C(_11739_),
    .Y(_11873_));
 AO21x1_ASAP7_75t_R _31632_ (.A1(_09496_),
    .A2(_11724_),
    .B(_11873_),
    .Y(_11874_));
 AO21x1_ASAP7_75t_R _31633_ (.A1(_11867_),
    .A2(_11726_),
    .B(_11874_),
    .Y(_04201_));
 INVx1_ASAP7_75t_R _31634_ (.A(_02012_),
    .Y(_11875_));
 NOR2x1_ASAP7_75t_R _31635_ (.A(net421),
    .B(_00210_),
    .Y(_11876_));
 AO21x1_ASAP7_75t_R _31636_ (.A1(net421),
    .A2(\cs_registers_i.pc_id_i[17] ),
    .B(_11876_),
    .Y(_11877_));
 NAND2x2_ASAP7_75t_R _31637_ (.A(_00385_),
    .B(_06174_),
    .Y(_11878_));
 TAPCELL_ASAP7_75t_R PHY_153 ();
 OA222x2_ASAP7_75t_R _31639_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11708_),
    .B2(_01624_),
    .C1(_11878_),
    .C2(net374),
    .Y(_11880_));
 INVx1_ASAP7_75t_R _31640_ (.A(_11880_),
    .Y(_11881_));
 OA211x2_ASAP7_75t_R _31641_ (.A1(_06165_),
    .A2(_11877_),
    .B(_11881_),
    .C(_11739_),
    .Y(_11882_));
 AO221x1_ASAP7_75t_R _31642_ (.A1(_09503_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11875_),
    .C(_11882_),
    .Y(_04202_));
 INVx1_ASAP7_75t_R _31643_ (.A(_02011_),
    .Y(_11883_));
 OAI22x1_ASAP7_75t_R _31644_ (.A1(_01623_),
    .A2(_11708_),
    .B1(_11878_),
    .B2(_00287_),
    .Y(_11884_));
 OAI21x1_ASAP7_75t_R _31645_ (.A1(net421),
    .A2(_02527_),
    .B(_00211_),
    .Y(_11885_));
 OR3x1_ASAP7_75t_R _31646_ (.A(net421),
    .B(_00211_),
    .C(_02527_),
    .Y(_11886_));
 AO21x1_ASAP7_75t_R _31647_ (.A1(_11885_),
    .A2(_11886_),
    .B(_06165_),
    .Y(_11887_));
 OA211x2_ASAP7_75t_R _31648_ (.A1(_06172_),
    .A2(_11884_),
    .B(_11887_),
    .C(_11739_),
    .Y(_11888_));
 AO21x1_ASAP7_75t_R _31649_ (.A1(_09512_),
    .A2(_11724_),
    .B(_11888_),
    .Y(_11889_));
 AO21x1_ASAP7_75t_R _31650_ (.A1(_11883_),
    .A2(_11726_),
    .B(_11889_),
    .Y(_04203_));
 INVx1_ASAP7_75t_R _31651_ (.A(_02010_),
    .Y(_11890_));
 NOR2x1_ASAP7_75t_R _31652_ (.A(_01722_),
    .B(_00213_),
    .Y(_11891_));
 AO21x1_ASAP7_75t_R _31653_ (.A1(_01722_),
    .A2(\cs_registers_i.pc_id_i[19] ),
    .B(_11891_),
    .Y(_11892_));
 OA222x2_ASAP7_75t_R _31654_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11708_),
    .B2(_01622_),
    .C1(_11878_),
    .C2(_00286_),
    .Y(_11893_));
 INVx1_ASAP7_75t_R _31655_ (.A(_11893_),
    .Y(_11894_));
 OA211x2_ASAP7_75t_R _31656_ (.A1(_06165_),
    .A2(_11892_),
    .B(_11894_),
    .C(_11739_),
    .Y(_11895_));
 AO221x1_ASAP7_75t_R _31657_ (.A1(_09519_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11890_),
    .C(_11895_),
    .Y(_04204_));
 INVx1_ASAP7_75t_R _31658_ (.A(_02009_),
    .Y(_11896_));
 OAI22x1_ASAP7_75t_R _31659_ (.A1(_01621_),
    .A2(_11708_),
    .B1(_11878_),
    .B2(net360),
    .Y(_11897_));
 OAI21x1_ASAP7_75t_R _31660_ (.A1(_01722_),
    .A2(_02528_),
    .B(_00214_),
    .Y(_11898_));
 OR3x1_ASAP7_75t_R _31661_ (.A(_01722_),
    .B(_00214_),
    .C(_02528_),
    .Y(_11899_));
 AO21x1_ASAP7_75t_R _31662_ (.A1(_11898_),
    .A2(_11899_),
    .B(_06165_),
    .Y(_11900_));
 OA211x2_ASAP7_75t_R _31663_ (.A1(_06172_),
    .A2(_11897_),
    .B(_11900_),
    .C(_11739_),
    .Y(_11901_));
 AO21x1_ASAP7_75t_R _31664_ (.A1(_09526_),
    .A2(_11724_),
    .B(_11901_),
    .Y(_11902_));
 AO21x1_ASAP7_75t_R _31665_ (.A1(_11896_),
    .A2(_11726_),
    .B(_11902_),
    .Y(_04205_));
 INVx1_ASAP7_75t_R _31666_ (.A(_02008_),
    .Y(_11903_));
 NOR2x1_ASAP7_75t_R _31667_ (.A(_01722_),
    .B(_00216_),
    .Y(_11904_));
 AO21x1_ASAP7_75t_R _31668_ (.A1(_01722_),
    .A2(\cs_registers_i.pc_id_i[21] ),
    .B(_11904_),
    .Y(_11905_));
 OA222x2_ASAP7_75t_R _31669_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11708_),
    .B2(_01620_),
    .C1(_11878_),
    .C2(_01745_),
    .Y(_11906_));
 INVx1_ASAP7_75t_R _31670_ (.A(_11906_),
    .Y(_11907_));
 OA211x2_ASAP7_75t_R _31671_ (.A1(_06165_),
    .A2(_11905_),
    .B(_11907_),
    .C(_11739_),
    .Y(_11908_));
 AO221x1_ASAP7_75t_R _31672_ (.A1(_09532_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11903_),
    .C(_11908_),
    .Y(_04206_));
 INVx1_ASAP7_75t_R _31673_ (.A(_02007_),
    .Y(_11909_));
 AO32x1_ASAP7_75t_R _31674_ (.A1(_13132_),
    .A2(_00385_),
    .A3(_06174_),
    .B1(_09225_),
    .B2(_11785_),
    .Y(_11910_));
 OAI21x1_ASAP7_75t_R _31675_ (.A1(_01722_),
    .A2(_02529_),
    .B(_00217_),
    .Y(_11911_));
 OR3x1_ASAP7_75t_R _31676_ (.A(_01722_),
    .B(_00217_),
    .C(_02529_),
    .Y(_11912_));
 AO21x1_ASAP7_75t_R _31677_ (.A1(_11911_),
    .A2(_11912_),
    .B(_06165_),
    .Y(_11913_));
 OA211x2_ASAP7_75t_R _31678_ (.A1(_06172_),
    .A2(_11910_),
    .B(_11913_),
    .C(_11739_),
    .Y(_11914_));
 AO21x1_ASAP7_75t_R _31679_ (.A1(_09539_),
    .A2(_11724_),
    .B(_11914_),
    .Y(_11915_));
 AO21x1_ASAP7_75t_R _31680_ (.A1(_11909_),
    .A2(_11726_),
    .B(_11915_),
    .Y(_04207_));
 INVx1_ASAP7_75t_R _31681_ (.A(_02006_),
    .Y(_11916_));
 NOR2x1_ASAP7_75t_R _31682_ (.A(net421),
    .B(_00219_),
    .Y(_11917_));
 AO21x1_ASAP7_75t_R _31683_ (.A1(net421),
    .A2(\cs_registers_i.pc_id_i[23] ),
    .B(_11917_),
    .Y(_11918_));
 OA222x2_ASAP7_75t_R _31684_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11708_),
    .B2(_01618_),
    .C1(_11878_),
    .C2(_00245_),
    .Y(_11919_));
 INVx1_ASAP7_75t_R _31685_ (.A(_11919_),
    .Y(_11920_));
 OA211x2_ASAP7_75t_R _31686_ (.A1(_06165_),
    .A2(_11918_),
    .B(_11920_),
    .C(_11739_),
    .Y(_11921_));
 AO21x1_ASAP7_75t_R _31687_ (.A1(_09545_),
    .A2(_11724_),
    .B(_11921_),
    .Y(_11922_));
 AO21x1_ASAP7_75t_R _31688_ (.A1(_11916_),
    .A2(_11726_),
    .B(_11922_),
    .Y(_04208_));
 INVx1_ASAP7_75t_R _31689_ (.A(_02005_),
    .Y(_11923_));
 OAI22x1_ASAP7_75t_R _31690_ (.A1(_01617_),
    .A2(_11708_),
    .B1(_11878_),
    .B2(net316),
    .Y(_11924_));
 OAI21x1_ASAP7_75t_R _31691_ (.A1(net421),
    .A2(_02530_),
    .B(_00220_),
    .Y(_11925_));
 OR3x1_ASAP7_75t_R _31692_ (.A(net421),
    .B(_00220_),
    .C(_02530_),
    .Y(_11926_));
 AO21x1_ASAP7_75t_R _31693_ (.A1(_11925_),
    .A2(_11926_),
    .B(_06165_),
    .Y(_11927_));
 OA211x2_ASAP7_75t_R _31694_ (.A1(_06172_),
    .A2(_11924_),
    .B(_11927_),
    .C(_11739_),
    .Y(_11928_));
 AO21x1_ASAP7_75t_R _31695_ (.A1(_11192_),
    .A2(_11724_),
    .B(_11928_),
    .Y(_11929_));
 AO21x1_ASAP7_75t_R _31696_ (.A1(_11923_),
    .A2(_11726_),
    .B(_11929_),
    .Y(_04209_));
 INVx1_ASAP7_75t_R _31697_ (.A(_02004_),
    .Y(_11930_));
 NOR2x1_ASAP7_75t_R _31698_ (.A(_01722_),
    .B(_00222_),
    .Y(_11931_));
 AO21x1_ASAP7_75t_R _31699_ (.A1(_01722_),
    .A2(\cs_registers_i.pc_id_i[25] ),
    .B(_11931_),
    .Y(_11932_));
 OA222x2_ASAP7_75t_R _31700_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_01743_),
    .B2(_11878_),
    .C1(_11708_),
    .C2(_01616_),
    .Y(_11933_));
 INVx1_ASAP7_75t_R _31701_ (.A(_11933_),
    .Y(_11934_));
 OA211x2_ASAP7_75t_R _31702_ (.A1(_06165_),
    .A2(_11932_),
    .B(_11934_),
    .C(_11739_),
    .Y(_11935_));
 AO221x1_ASAP7_75t_R _31703_ (.A1(_09565_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11930_),
    .C(_11935_),
    .Y(_04210_));
 INVx1_ASAP7_75t_R _31704_ (.A(_02003_),
    .Y(_11936_));
 AO32x1_ASAP7_75t_R _31705_ (.A1(_14141_),
    .A2(_00385_),
    .A3(_06174_),
    .B1(_09230_),
    .B2(_11785_),
    .Y(_11937_));
 OAI21x1_ASAP7_75t_R _31706_ (.A1(_01722_),
    .A2(_02531_),
    .B(_00223_),
    .Y(_11938_));
 OR3x1_ASAP7_75t_R _31707_ (.A(_01722_),
    .B(_00223_),
    .C(_02531_),
    .Y(_11939_));
 AO21x1_ASAP7_75t_R _31708_ (.A1(_11938_),
    .A2(_11939_),
    .B(_06165_),
    .Y(_11940_));
 OA211x2_ASAP7_75t_R _31709_ (.A1(_06172_),
    .A2(_11937_),
    .B(_11940_),
    .C(_11739_),
    .Y(_11941_));
 AO21x1_ASAP7_75t_R _31710_ (.A1(_09572_),
    .A2(_11724_),
    .B(_11941_),
    .Y(_11942_));
 AO21x1_ASAP7_75t_R _31711_ (.A1(_11936_),
    .A2(_11726_),
    .B(_11942_),
    .Y(_04211_));
 INVx1_ASAP7_75t_R _31712_ (.A(_02002_),
    .Y(_11943_));
 NOR2x1_ASAP7_75t_R _31713_ (.A(net421),
    .B(_00225_),
    .Y(_11944_));
 AO21x1_ASAP7_75t_R _31714_ (.A1(net421),
    .A2(\cs_registers_i.pc_id_i[27] ),
    .B(_11944_),
    .Y(_11945_));
 OA222x2_ASAP7_75t_R _31715_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_01742_),
    .B2(_11878_),
    .C1(_11708_),
    .C2(_01614_),
    .Y(_11946_));
 INVx1_ASAP7_75t_R _31716_ (.A(_11946_),
    .Y(_11947_));
 OA211x2_ASAP7_75t_R _31717_ (.A1(_06165_),
    .A2(_11945_),
    .B(_11947_),
    .C(_11739_),
    .Y(_11948_));
 AO221x1_ASAP7_75t_R _31718_ (.A1(_09578_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_11943_),
    .C(_11948_),
    .Y(_04212_));
 INVx1_ASAP7_75t_R _31719_ (.A(_02001_),
    .Y(_11949_));
 AO32x1_ASAP7_75t_R _31720_ (.A1(_00385_),
    .A2(_06174_),
    .A3(_14318_),
    .B1(_11785_),
    .B2(_09233_),
    .Y(_11950_));
 OAI21x1_ASAP7_75t_R _31721_ (.A1(_01722_),
    .A2(_02532_),
    .B(_00226_),
    .Y(_11951_));
 OR3x1_ASAP7_75t_R _31722_ (.A(_01722_),
    .B(_00226_),
    .C(_02532_),
    .Y(_11952_));
 AO21x1_ASAP7_75t_R _31723_ (.A1(_11951_),
    .A2(_11952_),
    .B(_06165_),
    .Y(_11953_));
 OA211x2_ASAP7_75t_R _31724_ (.A1(_06172_),
    .A2(_11950_),
    .B(_11953_),
    .C(_11739_),
    .Y(_11954_));
 AO21x1_ASAP7_75t_R _31725_ (.A1(_09585_),
    .A2(_11724_),
    .B(_11954_),
    .Y(_11955_));
 AO21x1_ASAP7_75t_R _31726_ (.A1(_11949_),
    .A2(_11726_),
    .B(_11955_),
    .Y(_04213_));
 NOR2x1_ASAP7_75t_R _31727_ (.A(_01722_),
    .B(_00228_),
    .Y(_11956_));
 AO21x1_ASAP7_75t_R _31728_ (.A1(_01722_),
    .A2(\cs_registers_i.pc_id_i[29] ),
    .B(_11956_),
    .Y(_11957_));
 OA222x2_ASAP7_75t_R _31729_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_01740_),
    .B2(_11878_),
    .C1(_11708_),
    .C2(_01612_),
    .Y(_11958_));
 INVx1_ASAP7_75t_R _31730_ (.A(_11958_),
    .Y(_11959_));
 OA211x2_ASAP7_75t_R _31731_ (.A1(_06165_),
    .A2(_11957_),
    .B(_11959_),
    .C(_11739_),
    .Y(_11960_));
 AO221x1_ASAP7_75t_R _31732_ (.A1(_09591_),
    .A2(_11720_),
    .B1(_11726_),
    .B2(_08501_),
    .C(_11960_),
    .Y(_04214_));
 INVx1_ASAP7_75t_R _31733_ (.A(_01999_),
    .Y(_11961_));
 AO32x1_ASAP7_75t_R _31734_ (.A1(_00385_),
    .A2(_06174_),
    .A3(_13369_),
    .B1(_11785_),
    .B2(_05326_),
    .Y(_11962_));
 OAI21x1_ASAP7_75t_R _31735_ (.A1(_01722_),
    .A2(_02533_),
    .B(_00229_),
    .Y(_11963_));
 OR3x1_ASAP7_75t_R _31736_ (.A(_01722_),
    .B(_00229_),
    .C(_02533_),
    .Y(_11964_));
 AO21x1_ASAP7_75t_R _31737_ (.A1(_11963_),
    .A2(_11964_),
    .B(_06165_),
    .Y(_11965_));
 OA211x2_ASAP7_75t_R _31738_ (.A1(_06172_),
    .A2(_11962_),
    .B(_11965_),
    .C(_11739_),
    .Y(_11966_));
 AO21x1_ASAP7_75t_R _31739_ (.A1(_11961_),
    .A2(_11726_),
    .B(_11966_),
    .Y(_11967_));
 AO21x1_ASAP7_75t_R _31740_ (.A1(_09598_),
    .A2(_11720_),
    .B(_11967_),
    .Y(_04215_));
 INVx1_ASAP7_75t_R _31741_ (.A(_01998_),
    .Y(_11968_));
 OR4x1_ASAP7_75t_R _31742_ (.A(_01722_),
    .B(_00227_),
    .C(_00229_),
    .D(_06053_),
    .Y(_11969_));
 XNOR2x1_ASAP7_75t_R _31743_ (.B(_11969_),
    .Y(_11970_),
    .A(_00230_));
 OA222x2_ASAP7_75t_R _31744_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11708_),
    .B2(_01610_),
    .C1(_11878_),
    .C2(_00280_),
    .Y(_11971_));
 AOI21x1_ASAP7_75t_R _31745_ (.A1(_06172_),
    .A2(_11970_),
    .B(_11971_),
    .Y(_11972_));
 AO32x1_ASAP7_75t_R _31746_ (.A1(_06340_),
    .A2(_11242_),
    .A3(_11972_),
    .B1(_11724_),
    .B2(_09605_),
    .Y(_11973_));
 AO21x1_ASAP7_75t_R _31747_ (.A1(_11968_),
    .A2(_11726_),
    .B(_11973_),
    .Y(_04216_));
 NAND2x1_ASAP7_75t_R _31748_ (.A(_01997_),
    .B(_11239_),
    .Y(_11974_));
 OA21x2_ASAP7_75t_R _31749_ (.A1(_09532_),
    .A2(_11239_),
    .B(_11974_),
    .Y(_04217_));
 NAND2x1_ASAP7_75t_R _31750_ (.A(_01996_),
    .B(_11239_),
    .Y(_11975_));
 OA21x2_ASAP7_75t_R _31751_ (.A1(_09503_),
    .A2(_11239_),
    .B(_11975_),
    .Y(_04218_));
 NAND2x2_ASAP7_75t_R _31752_ (.A(_11719_),
    .B(_11497_),
    .Y(_11976_));
 TAPCELL_ASAP7_75t_R PHY_152 ();
 TAPCELL_ASAP7_75t_R PHY_151 ();
 NAND2x1_ASAP7_75t_R _31755_ (.A(_01995_),
    .B(_11976_),
    .Y(_11979_));
 OA21x2_ASAP7_75t_R _31756_ (.A1(_10974_),
    .A2(_11976_),
    .B(_11979_),
    .Y(_04219_));
 NAND2x1_ASAP7_75t_R _31757_ (.A(_01994_),
    .B(_11976_),
    .Y(_11980_));
 OA21x2_ASAP7_75t_R _31758_ (.A1(_09363_),
    .A2(_11976_),
    .B(_11980_),
    .Y(_04220_));
 AO21x1_ASAP7_75t_R _31759_ (.A1(_11719_),
    .A2(_11497_),
    .B(_07369_),
    .Y(_11981_));
 OA21x2_ASAP7_75t_R _31760_ (.A1(_09390_),
    .A2(_11976_),
    .B(_11981_),
    .Y(_04221_));
 NAND2x1_ASAP7_75t_R _31761_ (.A(_01992_),
    .B(_11976_),
    .Y(_11982_));
 OA21x2_ASAP7_75t_R _31762_ (.A1(_09397_),
    .A2(_11976_),
    .B(_11982_),
    .Y(_04222_));
 NAND2x1_ASAP7_75t_R _31763_ (.A(_01991_),
    .B(_11976_),
    .Y(_11983_));
 OA21x2_ASAP7_75t_R _31764_ (.A1(_09408_),
    .A2(_11976_),
    .B(_11983_),
    .Y(_04223_));
 NAND2x1_ASAP7_75t_R _31765_ (.A(_01990_),
    .B(_11976_),
    .Y(_11984_));
 OA21x2_ASAP7_75t_R _31766_ (.A1(_09417_),
    .A2(_11976_),
    .B(_11984_),
    .Y(_04224_));
 NAND2x1_ASAP7_75t_R _31767_ (.A(_01989_),
    .B(_11976_),
    .Y(_11985_));
 OA21x2_ASAP7_75t_R _31768_ (.A1(_09426_),
    .A2(_11976_),
    .B(_11985_),
    .Y(_04225_));
 NAND2x1_ASAP7_75t_R _31769_ (.A(_01988_),
    .B(_11976_),
    .Y(_11986_));
 OA21x2_ASAP7_75t_R _31770_ (.A1(_09432_),
    .A2(_11976_),
    .B(_11986_),
    .Y(_04226_));
 NAND2x1_ASAP7_75t_R _31771_ (.A(_01987_),
    .B(_11976_),
    .Y(_11987_));
 OA21x2_ASAP7_75t_R _31772_ (.A1(_09438_),
    .A2(_11976_),
    .B(_11987_),
    .Y(_04227_));
 TAPCELL_ASAP7_75t_R PHY_150 ();
 NAND2x1_ASAP7_75t_R _31774_ (.A(_01986_),
    .B(_11976_),
    .Y(_11989_));
 OA21x2_ASAP7_75t_R _31775_ (.A1(_09445_),
    .A2(_11976_),
    .B(_11989_),
    .Y(_04228_));
 TAPCELL_ASAP7_75t_R PHY_149 ();
 NAND2x1_ASAP7_75t_R _31777_ (.A(_01985_),
    .B(_11976_),
    .Y(_11991_));
 OA21x2_ASAP7_75t_R _31778_ (.A1(_09452_),
    .A2(_11976_),
    .B(_11991_),
    .Y(_04229_));
 NAND2x1_ASAP7_75t_R _31779_ (.A(_01984_),
    .B(_11976_),
    .Y(_11992_));
 OA21x2_ASAP7_75t_R _31780_ (.A1(_09458_),
    .A2(_11976_),
    .B(_11992_),
    .Y(_04230_));
 NAND2x1_ASAP7_75t_R _31781_ (.A(_01983_),
    .B(_11976_),
    .Y(_11993_));
 OA21x2_ASAP7_75t_R _31782_ (.A1(_09465_),
    .A2(_11976_),
    .B(_11993_),
    .Y(_04231_));
 NAND2x1_ASAP7_75t_R _31783_ (.A(_01982_),
    .B(_11976_),
    .Y(_11994_));
 OA21x2_ASAP7_75t_R _31784_ (.A1(_09473_),
    .A2(_11976_),
    .B(_11994_),
    .Y(_04232_));
 NAND2x1_ASAP7_75t_R _31785_ (.A(_01981_),
    .B(_11976_),
    .Y(_11995_));
 OA21x2_ASAP7_75t_R _31786_ (.A1(_09481_),
    .A2(_11976_),
    .B(_11995_),
    .Y(_04233_));
 NAND2x1_ASAP7_75t_R _31787_ (.A(_01980_),
    .B(_11976_),
    .Y(_11996_));
 OA21x2_ASAP7_75t_R _31788_ (.A1(_09488_),
    .A2(_11976_),
    .B(_11996_),
    .Y(_04234_));
 NAND2x1_ASAP7_75t_R _31789_ (.A(_01979_),
    .B(_11976_),
    .Y(_11997_));
 OA21x2_ASAP7_75t_R _31790_ (.A1(_09496_),
    .A2(_11976_),
    .B(_11997_),
    .Y(_04235_));
 NAND2x1_ASAP7_75t_R _31791_ (.A(_01978_),
    .B(_11976_),
    .Y(_11998_));
 OA21x2_ASAP7_75t_R _31792_ (.A1(_09503_),
    .A2(_11976_),
    .B(_11998_),
    .Y(_04236_));
 NAND2x1_ASAP7_75t_R _31793_ (.A(_01977_),
    .B(_11976_),
    .Y(_11999_));
 OA21x2_ASAP7_75t_R _31794_ (.A1(_09512_),
    .A2(_11976_),
    .B(_11999_),
    .Y(_04237_));
 TAPCELL_ASAP7_75t_R PHY_148 ();
 NAND2x1_ASAP7_75t_R _31796_ (.A(_01976_),
    .B(_11976_),
    .Y(_12001_));
 OA21x2_ASAP7_75t_R _31797_ (.A1(_09519_),
    .A2(_11976_),
    .B(_12001_),
    .Y(_04238_));
 TAPCELL_ASAP7_75t_R PHY_147 ();
 NAND2x1_ASAP7_75t_R _31799_ (.A(_01975_),
    .B(_11976_),
    .Y(_12003_));
 OA21x2_ASAP7_75t_R _31800_ (.A1(_09526_),
    .A2(_11976_),
    .B(_12003_),
    .Y(_04239_));
 NAND2x1_ASAP7_75t_R _31801_ (.A(_01974_),
    .B(_11976_),
    .Y(_12004_));
 OA21x2_ASAP7_75t_R _31802_ (.A1(_09532_),
    .A2(_11976_),
    .B(_12004_),
    .Y(_04240_));
 NAND2x1_ASAP7_75t_R _31803_ (.A(_01973_),
    .B(_11976_),
    .Y(_12005_));
 OA21x2_ASAP7_75t_R _31804_ (.A1(_09539_),
    .A2(_11976_),
    .B(_12005_),
    .Y(_04241_));
 NAND2x1_ASAP7_75t_R _31805_ (.A(_01972_),
    .B(_11976_),
    .Y(_12006_));
 OA21x2_ASAP7_75t_R _31806_ (.A1(_09545_),
    .A2(_11976_),
    .B(_12006_),
    .Y(_04242_));
 NAND2x1_ASAP7_75t_R _31807_ (.A(_01971_),
    .B(_11976_),
    .Y(_12007_));
 OA21x2_ASAP7_75t_R _31808_ (.A1(_11192_),
    .A2(_11976_),
    .B(_12007_),
    .Y(_04243_));
 NAND2x1_ASAP7_75t_R _31809_ (.A(_01970_),
    .B(_11976_),
    .Y(_12008_));
 OA21x2_ASAP7_75t_R _31810_ (.A1(_09565_),
    .A2(_11976_),
    .B(_12008_),
    .Y(_04244_));
 NAND2x1_ASAP7_75t_R _31811_ (.A(_01969_),
    .B(_11976_),
    .Y(_12009_));
 OA21x2_ASAP7_75t_R _31812_ (.A1(_09572_),
    .A2(_11976_),
    .B(_12009_),
    .Y(_04245_));
 NAND2x1_ASAP7_75t_R _31813_ (.A(_01968_),
    .B(_11976_),
    .Y(_12010_));
 OA21x2_ASAP7_75t_R _31814_ (.A1(_09578_),
    .A2(_11976_),
    .B(_12010_),
    .Y(_04246_));
 NAND2x1_ASAP7_75t_R _31815_ (.A(_01967_),
    .B(_11976_),
    .Y(_12011_));
 OA21x2_ASAP7_75t_R _31816_ (.A1(_09585_),
    .A2(_11976_),
    .B(_12011_),
    .Y(_04247_));
 NAND2x1_ASAP7_75t_R _31817_ (.A(_01966_),
    .B(_11976_),
    .Y(_12012_));
 OA21x2_ASAP7_75t_R _31818_ (.A1(_09591_),
    .A2(_11976_),
    .B(_12012_),
    .Y(_04248_));
 NAND2x1_ASAP7_75t_R _31819_ (.A(_01965_),
    .B(_11976_),
    .Y(_12013_));
 OA21x2_ASAP7_75t_R _31820_ (.A1(_09598_),
    .A2(_11976_),
    .B(_12013_),
    .Y(_04249_));
 NAND2x1_ASAP7_75t_R _31821_ (.A(_01964_),
    .B(_11976_),
    .Y(_12014_));
 OA21x2_ASAP7_75t_R _31822_ (.A1(_09605_),
    .A2(_11976_),
    .B(_12014_),
    .Y(_04250_));
 TAPCELL_ASAP7_75t_R PHY_146 ();
 NAND2x2_ASAP7_75t_R _31824_ (.A(_06889_),
    .B(_11237_),
    .Y(_12016_));
 TAPCELL_ASAP7_75t_R PHY_145 ();
 TAPCELL_ASAP7_75t_R PHY_144 ();
 TAPCELL_ASAP7_75t_R PHY_143 ();
 AO21x1_ASAP7_75t_R _31828_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06197_),
    .Y(_12020_));
 OA21x2_ASAP7_75t_R _31829_ (.A1(_09496_),
    .A2(_12016_),
    .B(_12020_),
    .Y(_04251_));
 AO21x1_ASAP7_75t_R _31830_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06196_),
    .Y(_12021_));
 OA21x2_ASAP7_75t_R _31831_ (.A1(_09503_),
    .A2(_12016_),
    .B(_12021_),
    .Y(_04252_));
 AO21x1_ASAP7_75t_R _31832_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06194_),
    .Y(_12022_));
 OA21x2_ASAP7_75t_R _31833_ (.A1(_09512_),
    .A2(_12016_),
    .B(_12022_),
    .Y(_04253_));
 AO21x1_ASAP7_75t_R _31834_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06193_),
    .Y(_12023_));
 OA21x2_ASAP7_75t_R _31835_ (.A1(_09519_),
    .A2(_12016_),
    .B(_12023_),
    .Y(_04254_));
 AO21x1_ASAP7_75t_R _31836_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06203_),
    .Y(_12024_));
 OA21x2_ASAP7_75t_R _31837_ (.A1(_09526_),
    .A2(_12016_),
    .B(_12024_),
    .Y(_04255_));
 AO21x1_ASAP7_75t_R _31838_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06202_),
    .Y(_12025_));
 OA21x2_ASAP7_75t_R _31839_ (.A1(_09532_),
    .A2(_12016_),
    .B(_12025_),
    .Y(_04256_));
 AO21x1_ASAP7_75t_R _31840_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06200_),
    .Y(_12026_));
 OA21x2_ASAP7_75t_R _31841_ (.A1(_09539_),
    .A2(_12016_),
    .B(_12026_),
    .Y(_04257_));
 AO21x1_ASAP7_75t_R _31842_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06199_),
    .Y(_12027_));
 OA21x2_ASAP7_75t_R _31843_ (.A1(_09545_),
    .A2(_12016_),
    .B(_12027_),
    .Y(_04258_));
 AO21x1_ASAP7_75t_R _31844_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06217_),
    .Y(_12028_));
 OA21x2_ASAP7_75t_R _31845_ (.A1(_11192_),
    .A2(_12016_),
    .B(_12028_),
    .Y(_04259_));
 AO21x1_ASAP7_75t_R _31846_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06216_),
    .Y(_12029_));
 OA21x2_ASAP7_75t_R _31847_ (.A1(_09565_),
    .A2(_12016_),
    .B(_12029_),
    .Y(_04260_));
 AO21x1_ASAP7_75t_R _31848_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06220_),
    .Y(_12030_));
 OA21x2_ASAP7_75t_R _31849_ (.A1(_09572_),
    .A2(_12016_),
    .B(_12030_),
    .Y(_04261_));
 AO21x1_ASAP7_75t_R _31850_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06219_),
    .Y(_12031_));
 OA21x2_ASAP7_75t_R _31851_ (.A1(_09578_),
    .A2(_12016_),
    .B(_12031_),
    .Y(_04262_));
 AO21x1_ASAP7_75t_R _31852_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06207_),
    .Y(_12032_));
 OA21x2_ASAP7_75t_R _31853_ (.A1(_09585_),
    .A2(_12016_),
    .B(_12032_),
    .Y(_04263_));
 AO21x1_ASAP7_75t_R _31854_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06208_),
    .Y(_12033_));
 OA21x2_ASAP7_75t_R _31855_ (.A1(_09591_),
    .A2(_12016_),
    .B(_12033_),
    .Y(_04264_));
 AO21x1_ASAP7_75t_R _31856_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06206_),
    .Y(_12034_));
 OA21x2_ASAP7_75t_R _31857_ (.A1(_09598_),
    .A2(_12016_),
    .B(_12034_),
    .Y(_04265_));
 AO21x1_ASAP7_75t_R _31858_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06212_),
    .Y(_12035_));
 OA21x2_ASAP7_75t_R _31859_ (.A1(_09458_),
    .A2(_12016_),
    .B(_12035_),
    .Y(_04266_));
 AO21x1_ASAP7_75t_R _31860_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06214_),
    .Y(_12036_));
 OA21x2_ASAP7_75t_R _31861_ (.A1(_09432_),
    .A2(_12016_),
    .B(_12036_),
    .Y(_04267_));
 AO21x1_ASAP7_75t_R _31862_ (.A1(_06889_),
    .A2(_11237_),
    .B(_06211_),
    .Y(_12037_));
 OA21x2_ASAP7_75t_R _31863_ (.A1(_09397_),
    .A2(_12016_),
    .B(_12037_),
    .Y(_04268_));
 AND3x1_ASAP7_75t_R _31864_ (.A(_05629_),
    .B(_07515_),
    .C(_06903_),
    .Y(_12038_));
 AO21x2_ASAP7_75t_R _31865_ (.A1(_09365_),
    .A2(_12038_),
    .B(_11244_),
    .Y(_12039_));
 TAPCELL_ASAP7_75t_R PHY_142 ();
 OAI22x1_ASAP7_75t_R _31867_ (.A1(_01907_),
    .A2(_11231_),
    .B1(_12039_),
    .B2(_01945_),
    .Y(_04269_));
 AND4x1_ASAP7_75t_R _31868_ (.A(_01311_),
    .B(_06873_),
    .C(_09375_),
    .D(_11224_),
    .Y(_12041_));
 AOI21x1_ASAP7_75t_R _31869_ (.A1(_09365_),
    .A2(_12038_),
    .B(_11244_),
    .Y(_12042_));
 OA211x2_ASAP7_75t_R _31870_ (.A1(_01906_),
    .A2(_11231_),
    .B(_12039_),
    .C(_11225_),
    .Y(_12043_));
 OA21x2_ASAP7_75t_R _31871_ (.A1(_11107_),
    .A2(_11243_),
    .B(_12043_),
    .Y(_12044_));
 AO21x1_ASAP7_75t_R _31872_ (.A1(_01944_),
    .A2(_12042_),
    .B(_12044_),
    .Y(_12045_));
 NOR2x1_ASAP7_75t_R _31873_ (.A(_12041_),
    .B(_12045_),
    .Y(_04270_));
 TAPCELL_ASAP7_75t_R PHY_141 ();
 TAPCELL_ASAP7_75t_R PHY_140 ();
 AOI22x1_ASAP7_75t_R _31876_ (.A1(_09380_),
    .A2(_11242_),
    .B1(_11243_),
    .B2(_01905_),
    .Y(_12048_));
 OA211x2_ASAP7_75t_R _31877_ (.A1(_09390_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12048_),
    .Y(_12049_));
 AO21x1_ASAP7_75t_R _31878_ (.A1(_07377_),
    .A2(_12042_),
    .B(_12049_),
    .Y(_04271_));
 INVx1_ASAP7_75t_R _31879_ (.A(_01942_),
    .Y(_12050_));
 AOI22x1_ASAP7_75t_R _31880_ (.A1(_09400_),
    .A2(_11242_),
    .B1(_11243_),
    .B2(_01904_),
    .Y(_12051_));
 OA211x2_ASAP7_75t_R _31881_ (.A1(_09397_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12051_),
    .Y(_12052_));
 AO21x1_ASAP7_75t_R _31882_ (.A1(_12050_),
    .A2(_12042_),
    .B(_12052_),
    .Y(_04272_));
 INVx1_ASAP7_75t_R _31883_ (.A(_01941_),
    .Y(_12053_));
 AOI22x1_ASAP7_75t_R _31884_ (.A1(_09412_),
    .A2(_11242_),
    .B1(_11243_),
    .B2(_01903_),
    .Y(_12054_));
 OA211x2_ASAP7_75t_R _31885_ (.A1(_09408_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12054_),
    .Y(_12055_));
 AO21x1_ASAP7_75t_R _31886_ (.A1(_12053_),
    .A2(net271),
    .B(_12055_),
    .Y(_04273_));
 TAPCELL_ASAP7_75t_R PHY_139 ();
 TAPCELL_ASAP7_75t_R PHY_138 ();
 TAPCELL_ASAP7_75t_R PHY_137 ();
 OA22x2_ASAP7_75t_R _31890_ (.A1(_09421_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01902_),
    .Y(_12059_));
 OA211x2_ASAP7_75t_R _31891_ (.A1(_11010_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12059_),
    .Y(_12060_));
 AOI21x1_ASAP7_75t_R _31892_ (.A1(_01940_),
    .A2(net271),
    .B(_12060_),
    .Y(_04274_));
 TAPCELL_ASAP7_75t_R PHY_136 ();
 NOR2x2_ASAP7_75t_R _31894_ (.A(_11242_),
    .B(_11243_),
    .Y(_12062_));
 TAPCELL_ASAP7_75t_R PHY_135 ();
 TAPCELL_ASAP7_75t_R PHY_134 ();
 OAI22x1_ASAP7_75t_R _31897_ (.A1(_09428_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01901_),
    .Y(_12065_));
 AO21x1_ASAP7_75t_R _31898_ (.A1(_09426_),
    .A2(_12062_),
    .B(_12065_),
    .Y(_12066_));
 TAPCELL_ASAP7_75t_R PHY_133 ();
 NAND2x1_ASAP7_75t_R _31900_ (.A(_01939_),
    .B(_12042_),
    .Y(_12068_));
 OA21x2_ASAP7_75t_R _31901_ (.A1(_12042_),
    .A2(_12066_),
    .B(_12068_),
    .Y(_04275_));
 OA22x2_ASAP7_75t_R _31902_ (.A1(_09434_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01900_),
    .Y(_12069_));
 OA211x2_ASAP7_75t_R _31903_ (.A1(_11236_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12069_),
    .Y(_12070_));
 AOI21x1_ASAP7_75t_R _31904_ (.A1(_01938_),
    .A2(net271),
    .B(_12070_),
    .Y(_04276_));
 INVx1_ASAP7_75t_R _31905_ (.A(_09438_),
    .Y(_12071_));
 OA22x2_ASAP7_75t_R _31906_ (.A1(_09440_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01899_),
    .Y(_12072_));
 OA211x2_ASAP7_75t_R _31907_ (.A1(_12071_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12072_),
    .Y(_12073_));
 AOI21x1_ASAP7_75t_R _31908_ (.A1(_01937_),
    .A2(_12042_),
    .B(_12073_),
    .Y(_04277_));
 OAI22x1_ASAP7_75t_R _31909_ (.A1(_09447_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01898_),
    .Y(_12074_));
 AO21x1_ASAP7_75t_R _31910_ (.A1(_09445_),
    .A2(_12062_),
    .B(_12074_),
    .Y(_12075_));
 NAND2x1_ASAP7_75t_R _31911_ (.A(_01936_),
    .B(_12042_),
    .Y(_12076_));
 OA21x2_ASAP7_75t_R _31912_ (.A1(_12042_),
    .A2(_12075_),
    .B(_12076_),
    .Y(_04278_));
 OAI22x1_ASAP7_75t_R _31913_ (.A1(_09454_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01897_),
    .Y(_12077_));
 AO21x1_ASAP7_75t_R _31914_ (.A1(_09452_),
    .A2(_12062_),
    .B(_12077_),
    .Y(_12078_));
 NAND2x1_ASAP7_75t_R _31915_ (.A(_01935_),
    .B(_12042_),
    .Y(_12079_));
 OA21x2_ASAP7_75t_R _31916_ (.A1(_12042_),
    .A2(_12078_),
    .B(_12079_),
    .Y(_04279_));
 OAI22x1_ASAP7_75t_R _31917_ (.A1(_09461_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01896_),
    .Y(_12080_));
 AO21x1_ASAP7_75t_R _31918_ (.A1(_09458_),
    .A2(_12062_),
    .B(_12080_),
    .Y(_12081_));
 NAND2x1_ASAP7_75t_R _31919_ (.A(_01934_),
    .B(net272),
    .Y(_12082_));
 OA21x2_ASAP7_75t_R _31920_ (.A1(net272),
    .A2(_12081_),
    .B(_12082_),
    .Y(_04280_));
 OAI22x1_ASAP7_75t_R _31921_ (.A1(_09468_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01895_),
    .Y(_12083_));
 AO21x1_ASAP7_75t_R _31922_ (.A1(_09465_),
    .A2(_12062_),
    .B(_12083_),
    .Y(_12084_));
 NAND2x1_ASAP7_75t_R _31923_ (.A(_01933_),
    .B(_12042_),
    .Y(_12085_));
 OA21x2_ASAP7_75t_R _31924_ (.A1(_12042_),
    .A2(_12084_),
    .B(_12085_),
    .Y(_04281_));
 TAPCELL_ASAP7_75t_R PHY_132 ();
 OA22x2_ASAP7_75t_R _31926_ (.A1(_09476_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01894_),
    .Y(_12087_));
 OA211x2_ASAP7_75t_R _31927_ (.A1(_11643_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12087_),
    .Y(_12088_));
 AOI21x1_ASAP7_75t_R _31928_ (.A1(_01932_),
    .A2(net272),
    .B(_12088_),
    .Y(_04282_));
 OAI22x1_ASAP7_75t_R _31929_ (.A1(_09483_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01893_),
    .Y(_12089_));
 AO21x1_ASAP7_75t_R _31930_ (.A1(_09481_),
    .A2(_12062_),
    .B(_12089_),
    .Y(_12090_));
 NAND2x1_ASAP7_75t_R _31931_ (.A(_01931_),
    .B(net272),
    .Y(_12091_));
 OA21x2_ASAP7_75t_R _31932_ (.A1(net272),
    .A2(_12090_),
    .B(_12091_),
    .Y(_04283_));
 OAI22x1_ASAP7_75t_R _31933_ (.A1(_09491_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01892_),
    .Y(_12092_));
 AO21x1_ASAP7_75t_R _31934_ (.A1(_09488_),
    .A2(_12062_),
    .B(_12092_),
    .Y(_12093_));
 NAND2x1_ASAP7_75t_R _31935_ (.A(_01930_),
    .B(net272),
    .Y(_12094_));
 OA21x2_ASAP7_75t_R _31936_ (.A1(net272),
    .A2(_12093_),
    .B(_12094_),
    .Y(_04284_));
 INVx1_ASAP7_75t_R _31937_ (.A(_09496_),
    .Y(_12095_));
 OA22x2_ASAP7_75t_R _31938_ (.A1(_09499_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01891_),
    .Y(_12096_));
 OA211x2_ASAP7_75t_R _31939_ (.A1(_12095_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12096_),
    .Y(_12097_));
 AOI21x1_ASAP7_75t_R _31940_ (.A1(_01929_),
    .A2(net271),
    .B(_12097_),
    .Y(_04285_));
 TAPCELL_ASAP7_75t_R PHY_131 ();
 OAI22x1_ASAP7_75t_R _31942_ (.A1(_09506_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01890_),
    .Y(_12099_));
 AO21x1_ASAP7_75t_R _31943_ (.A1(_09503_),
    .A2(_12062_),
    .B(_12099_),
    .Y(_12100_));
 NAND2x1_ASAP7_75t_R _31944_ (.A(_01928_),
    .B(net272),
    .Y(_12101_));
 OA21x2_ASAP7_75t_R _31945_ (.A1(net272),
    .A2(_12100_),
    .B(_12101_),
    .Y(_04286_));
 AO21x2_ASAP7_75t_R _31946_ (.A1(_18196_),
    .A2(_08133_),
    .B(_09511_),
    .Y(_12102_));
 OA22x2_ASAP7_75t_R _31947_ (.A1(_09515_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01889_),
    .Y(_12103_));
 OA211x2_ASAP7_75t_R _31948_ (.A1(_12102_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12103_),
    .Y(_12104_));
 AOI21x1_ASAP7_75t_R _31949_ (.A1(_01927_),
    .A2(net271),
    .B(_12104_),
    .Y(_04287_));
 OAI22x1_ASAP7_75t_R _31950_ (.A1(_09522_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01888_),
    .Y(_12105_));
 AO21x1_ASAP7_75t_R _31951_ (.A1(_09519_),
    .A2(_12062_),
    .B(_12105_),
    .Y(_12106_));
 NAND2x1_ASAP7_75t_R _31952_ (.A(_01926_),
    .B(net272),
    .Y(_12107_));
 OA21x2_ASAP7_75t_R _31953_ (.A1(net272),
    .A2(_12106_),
    .B(_12107_),
    .Y(_04288_));
 OAI22x1_ASAP7_75t_R _31954_ (.A1(_09528_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01887_),
    .Y(_12108_));
 AO21x1_ASAP7_75t_R _31955_ (.A1(_09526_),
    .A2(_12062_),
    .B(_12108_),
    .Y(_12109_));
 NAND2x1_ASAP7_75t_R _31956_ (.A(_01925_),
    .B(net271),
    .Y(_12110_));
 OA21x2_ASAP7_75t_R _31957_ (.A1(net271),
    .A2(_12109_),
    .B(_12110_),
    .Y(_04289_));
 OAI22x1_ASAP7_75t_R _31958_ (.A1(_09535_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01886_),
    .Y(_12111_));
 AO21x1_ASAP7_75t_R _31959_ (.A1(_09532_),
    .A2(_12062_),
    .B(_12111_),
    .Y(_12112_));
 NAND2x1_ASAP7_75t_R _31960_ (.A(_01924_),
    .B(net272),
    .Y(_12113_));
 OA21x2_ASAP7_75t_R _31961_ (.A1(net272),
    .A2(_12112_),
    .B(_12113_),
    .Y(_04290_));
 OAI22x1_ASAP7_75t_R _31962_ (.A1(_09541_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01885_),
    .Y(_12114_));
 AO21x1_ASAP7_75t_R _31963_ (.A1(_09539_),
    .A2(_12062_),
    .B(_12114_),
    .Y(_12115_));
 NAND2x1_ASAP7_75t_R _31964_ (.A(_01923_),
    .B(net271),
    .Y(_12116_));
 OA21x2_ASAP7_75t_R _31965_ (.A1(net271),
    .A2(_12115_),
    .B(_12116_),
    .Y(_04291_));
 OA22x2_ASAP7_75t_R _31966_ (.A1(_09548_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01884_),
    .Y(_12117_));
 OA211x2_ASAP7_75t_R _31967_ (.A1(_11673_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12117_),
    .Y(_12118_));
 AOI21x1_ASAP7_75t_R _31968_ (.A1(_01922_),
    .A2(net272),
    .B(_12118_),
    .Y(_04292_));
 OA22x2_ASAP7_75t_R _31969_ (.A1(_09551_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01883_),
    .Y(_12119_));
 OA211x2_ASAP7_75t_R _31970_ (.A1(_09560_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12119_),
    .Y(_12120_));
 AOI21x1_ASAP7_75t_R _31971_ (.A1(_01921_),
    .A2(net272),
    .B(_12120_),
    .Y(_04293_));
 INVx1_ASAP7_75t_R _31972_ (.A(_09565_),
    .Y(_12121_));
 OA22x2_ASAP7_75t_R _31973_ (.A1(_09568_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01882_),
    .Y(_12122_));
 OA211x2_ASAP7_75t_R _31974_ (.A1(_12121_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12122_),
    .Y(_12123_));
 AOI21x1_ASAP7_75t_R _31975_ (.A1(_01920_),
    .A2(net272),
    .B(_12123_),
    .Y(_04294_));
 INVx1_ASAP7_75t_R _31976_ (.A(_09572_),
    .Y(_12124_));
 OA22x2_ASAP7_75t_R _31977_ (.A1(_09574_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01881_),
    .Y(_12125_));
 OA211x2_ASAP7_75t_R _31978_ (.A1(_12124_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12125_),
    .Y(_12126_));
 AOI21x1_ASAP7_75t_R _31979_ (.A1(_01919_),
    .A2(net272),
    .B(_12126_),
    .Y(_04295_));
 OA22x2_ASAP7_75t_R _31980_ (.A1(_09581_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01880_),
    .Y(_12127_));
 OA211x2_ASAP7_75t_R _31981_ (.A1(_11203_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12127_),
    .Y(_12128_));
 AOI21x1_ASAP7_75t_R _31982_ (.A1(_01918_),
    .A2(net272),
    .B(_12128_),
    .Y(_04296_));
 OAI22x1_ASAP7_75t_R _31983_ (.A1(_09587_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01879_),
    .Y(_12129_));
 AO21x1_ASAP7_75t_R _31984_ (.A1(_09585_),
    .A2(_12062_),
    .B(_12129_),
    .Y(_12130_));
 NAND2x1_ASAP7_75t_R _31985_ (.A(_01917_),
    .B(net271),
    .Y(_12131_));
 OA21x2_ASAP7_75t_R _31986_ (.A1(net271),
    .A2(_12130_),
    .B(_12131_),
    .Y(_04297_));
 OA22x2_ASAP7_75t_R _31987_ (.A1(_09594_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01878_),
    .Y(_12132_));
 OA211x2_ASAP7_75t_R _31988_ (.A1(_11209_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12132_),
    .Y(_12133_));
 AOI21x1_ASAP7_75t_R _31989_ (.A1(_01916_),
    .A2(net272),
    .B(_12133_),
    .Y(_04298_));
 OAI22x1_ASAP7_75t_R _31990_ (.A1(_09600_),
    .A2(_11226_),
    .B1(_11231_),
    .B2(_01877_),
    .Y(_12134_));
 AO21x1_ASAP7_75t_R _31991_ (.A1(_09598_),
    .A2(_12062_),
    .B(_12134_),
    .Y(_12135_));
 NAND2x1_ASAP7_75t_R _31992_ (.A(_01915_),
    .B(net271),
    .Y(_12136_));
 OA21x2_ASAP7_75t_R _31993_ (.A1(net271),
    .A2(_12135_),
    .B(_12136_),
    .Y(_04299_));
 INVx1_ASAP7_75t_R _31994_ (.A(_01914_),
    .Y(_12137_));
 AOI22x1_ASAP7_75t_R _31995_ (.A1(_09607_),
    .A2(_11242_),
    .B1(_11243_),
    .B2(_01876_),
    .Y(_12138_));
 OA211x2_ASAP7_75t_R _31996_ (.A1(_09605_),
    .A2(_11244_),
    .B(_12039_),
    .C(_12138_),
    .Y(_12139_));
 AO21x1_ASAP7_75t_R _31997_ (.A1(_12137_),
    .A2(net271),
    .B(_12139_),
    .Y(_04300_));
 AOI21x1_ASAP7_75t_R _31998_ (.A1(_05627_),
    .A2(_11599_),
    .B(_11244_),
    .Y(_12140_));
 AO21x2_ASAP7_75t_R _31999_ (.A1(_05627_),
    .A2(_11599_),
    .B(_11244_),
    .Y(_12141_));
 AND3x1_ASAP7_75t_R _32000_ (.A(net309),
    .B(_01311_),
    .C(_06170_),
    .Y(_12142_));
 AO21x1_ASAP7_75t_R _32001_ (.A1(net360),
    .A2(_05708_),
    .B(_12142_),
    .Y(_12143_));
 AND3x1_ASAP7_75t_R _32002_ (.A(_01745_),
    .B(_06832_),
    .C(_12143_),
    .Y(_12144_));
 OR3x1_ASAP7_75t_R _32003_ (.A(_06172_),
    .B(_11785_),
    .C(_12144_),
    .Y(_12145_));
 AOI21x1_ASAP7_75t_R _32004_ (.A1(_06340_),
    .A2(_12145_),
    .B(_06252_),
    .Y(_12146_));
 OA22x2_ASAP7_75t_R _32005_ (.A1(_02104_),
    .A2(_11231_),
    .B1(_12146_),
    .B2(_11226_),
    .Y(_12147_));
 OA211x2_ASAP7_75t_R _32006_ (.A1(_10973_),
    .A2(_11244_),
    .B(_12141_),
    .C(_12147_),
    .Y(_12148_));
 AOI21x1_ASAP7_75t_R _32007_ (.A1(_01913_),
    .A2(_12140_),
    .B(_12148_),
    .Y(_04301_));
 AO21x1_ASAP7_75t_R _32008_ (.A1(_01745_),
    .A2(_06831_),
    .B(_01725_),
    .Y(_12149_));
 NAND2x1_ASAP7_75t_R _32009_ (.A(_01312_),
    .B(_12149_),
    .Y(_12150_));
 OA211x2_ASAP7_75t_R _32010_ (.A1(_12144_),
    .A2(_12150_),
    .B(_06165_),
    .C(_06340_),
    .Y(_12151_));
 NOR2x1_ASAP7_75t_R _32011_ (.A(_06288_),
    .B(_12151_),
    .Y(_12152_));
 AND4x1_ASAP7_75t_R _32012_ (.A(_01311_),
    .B(_06873_),
    .C(_11224_),
    .D(_12152_),
    .Y(_12153_));
 OA211x2_ASAP7_75t_R _32013_ (.A1(_02103_),
    .A2(_11231_),
    .B(_12141_),
    .C(_11225_),
    .Y(_12154_));
 OA21x2_ASAP7_75t_R _32014_ (.A1(_11107_),
    .A2(_11243_),
    .B(_12154_),
    .Y(_12155_));
 AOI211x1_ASAP7_75t_R _32015_ (.A1(_01912_),
    .A2(_12140_),
    .B(_12153_),
    .C(_12155_),
    .Y(_04302_));
 OA211x2_ASAP7_75t_R _32016_ (.A1(_06846_),
    .A2(_11708_),
    .B(_11242_),
    .C(_06299_),
    .Y(_12156_));
 AO221x1_ASAP7_75t_R _32017_ (.A1(_02102_),
    .A2(_11243_),
    .B1(_12062_),
    .B2(_09391_),
    .C(_12156_),
    .Y(_12157_));
 OR2x2_ASAP7_75t_R _32018_ (.A(_01911_),
    .B(_12141_),
    .Y(_12158_));
 OAI21x1_ASAP7_75t_R _32019_ (.A1(_12140_),
    .A2(_12157_),
    .B(_12158_),
    .Y(_04303_));
 INVx1_ASAP7_75t_R _32020_ (.A(_01910_),
    .Y(_12159_));
 AND3x1_ASAP7_75t_R _32021_ (.A(_14155_),
    .B(_06340_),
    .C(_06832_),
    .Y(_12160_));
 OA33x2_ASAP7_75t_R _32022_ (.A1(_01718_),
    .A2(_11493_),
    .A3(_06262_),
    .B1(_06308_),
    .B2(_11226_),
    .B3(_12160_),
    .Y(_12161_));
 OA211x2_ASAP7_75t_R _32023_ (.A1(_09397_),
    .A2(_11244_),
    .B(_12141_),
    .C(_12161_),
    .Y(_12162_));
 AO21x1_ASAP7_75t_R _32024_ (.A1(_12159_),
    .A2(_12140_),
    .B(_12162_),
    .Y(_04304_));
 INVx1_ASAP7_75t_R _32025_ (.A(_09408_),
    .Y(_12163_));
 OA21x2_ASAP7_75t_R _32026_ (.A1(_02100_),
    .A2(_11231_),
    .B(_06318_),
    .Y(_12164_));
 OA211x2_ASAP7_75t_R _32027_ (.A1(_12163_),
    .A2(_11244_),
    .B(_12141_),
    .C(_12164_),
    .Y(_12165_));
 AOI21x1_ASAP7_75t_R _32028_ (.A1(_01909_),
    .A2(_12140_),
    .B(_12165_),
    .Y(_04305_));
 OA21x2_ASAP7_75t_R _32029_ (.A1(_02099_),
    .A2(_11231_),
    .B(_06224_),
    .Y(_12166_));
 OA211x2_ASAP7_75t_R _32030_ (.A1(_11215_),
    .A2(_11244_),
    .B(_12141_),
    .C(_12166_),
    .Y(_12167_));
 AOI21x1_ASAP7_75t_R _32031_ (.A1(_01908_),
    .A2(_12140_),
    .B(_12167_),
    .Y(_04306_));
 TAPCELL_ASAP7_75t_R PHY_130 ();
 AND2x2_ASAP7_75t_R _32033_ (.A(_01945_),
    .B(_11242_),
    .Y(_12169_));
 AOI21x1_ASAP7_75t_R _32034_ (.A1(_01907_),
    .A2(_11226_),
    .B(_12169_),
    .Y(_04307_));
 AND2x2_ASAP7_75t_R _32035_ (.A(_01944_),
    .B(_11242_),
    .Y(_12170_));
 AOI21x1_ASAP7_75t_R _32036_ (.A1(_01906_),
    .A2(_11226_),
    .B(_12170_),
    .Y(_04308_));
 TAPCELL_ASAP7_75t_R PHY_129 ();
 NAND2x1_ASAP7_75t_R _32038_ (.A(_01905_),
    .B(_11226_),
    .Y(_12172_));
 OA21x2_ASAP7_75t_R _32039_ (.A1(_07377_),
    .A2(_11226_),
    .B(_12172_),
    .Y(_04309_));
 NAND2x1_ASAP7_75t_R _32040_ (.A(_01904_),
    .B(_11226_),
    .Y(_12173_));
 OA21x2_ASAP7_75t_R _32041_ (.A1(_12050_),
    .A2(_11226_),
    .B(_12173_),
    .Y(_04310_));
 NAND2x1_ASAP7_75t_R _32042_ (.A(_01903_),
    .B(_11226_),
    .Y(_12174_));
 OA21x2_ASAP7_75t_R _32043_ (.A1(_12053_),
    .A2(_11226_),
    .B(_12174_),
    .Y(_04311_));
 TAPCELL_ASAP7_75t_R PHY_128 ();
 AND2x2_ASAP7_75t_R _32045_ (.A(_01940_),
    .B(_11242_),
    .Y(_12176_));
 AOI21x1_ASAP7_75t_R _32046_ (.A1(_01902_),
    .A2(_11226_),
    .B(_12176_),
    .Y(_04312_));
 AND2x2_ASAP7_75t_R _32047_ (.A(_01939_),
    .B(_11242_),
    .Y(_12177_));
 AOI21x1_ASAP7_75t_R _32048_ (.A1(_01901_),
    .A2(_11226_),
    .B(_12177_),
    .Y(_04313_));
 AND2x2_ASAP7_75t_R _32049_ (.A(_01938_),
    .B(_11242_),
    .Y(_12178_));
 AOI21x1_ASAP7_75t_R _32050_ (.A1(_01900_),
    .A2(_11226_),
    .B(_12178_),
    .Y(_04314_));
 AND2x2_ASAP7_75t_R _32051_ (.A(_01937_),
    .B(_11242_),
    .Y(_12179_));
 AOI21x1_ASAP7_75t_R _32052_ (.A1(_01899_),
    .A2(_11226_),
    .B(_12179_),
    .Y(_04315_));
 AND2x2_ASAP7_75t_R _32053_ (.A(_01936_),
    .B(_11242_),
    .Y(_12180_));
 AOI21x1_ASAP7_75t_R _32054_ (.A1(_01898_),
    .A2(_11226_),
    .B(_12180_),
    .Y(_04316_));
 AND2x2_ASAP7_75t_R _32055_ (.A(_01935_),
    .B(_11242_),
    .Y(_12181_));
 AOI21x1_ASAP7_75t_R _32056_ (.A1(_01897_),
    .A2(_11226_),
    .B(_12181_),
    .Y(_04317_));
 AND2x2_ASAP7_75t_R _32057_ (.A(_01934_),
    .B(_11242_),
    .Y(_12182_));
 AOI21x1_ASAP7_75t_R _32058_ (.A1(_01896_),
    .A2(_11226_),
    .B(_12182_),
    .Y(_04318_));
 AND2x2_ASAP7_75t_R _32059_ (.A(_01933_),
    .B(_11242_),
    .Y(_12183_));
 AOI21x1_ASAP7_75t_R _32060_ (.A1(_01895_),
    .A2(_11226_),
    .B(_12183_),
    .Y(_04319_));
 TAPCELL_ASAP7_75t_R PHY_127 ();
 AND2x2_ASAP7_75t_R _32062_ (.A(_01932_),
    .B(_11242_),
    .Y(_12185_));
 AOI21x1_ASAP7_75t_R _32063_ (.A1(_01894_),
    .A2(_11226_),
    .B(_12185_),
    .Y(_04320_));
 AND2x2_ASAP7_75t_R _32064_ (.A(_01931_),
    .B(_11242_),
    .Y(_12186_));
 AOI21x1_ASAP7_75t_R _32065_ (.A1(_01893_),
    .A2(_11226_),
    .B(_12186_),
    .Y(_04321_));
 TAPCELL_ASAP7_75t_R PHY_126 ();
 AND2x2_ASAP7_75t_R _32067_ (.A(_01930_),
    .B(_11242_),
    .Y(_12188_));
 AOI21x1_ASAP7_75t_R _32068_ (.A1(_01892_),
    .A2(_11226_),
    .B(_12188_),
    .Y(_04322_));
 AND2x2_ASAP7_75t_R _32069_ (.A(_01929_),
    .B(_11242_),
    .Y(_12189_));
 AOI21x1_ASAP7_75t_R _32070_ (.A1(_01891_),
    .A2(_11226_),
    .B(_12189_),
    .Y(_04323_));
 AND2x2_ASAP7_75t_R _32071_ (.A(_01928_),
    .B(_11242_),
    .Y(_12190_));
 AOI21x1_ASAP7_75t_R _32072_ (.A1(_01890_),
    .A2(_11226_),
    .B(_12190_),
    .Y(_04324_));
 AND2x2_ASAP7_75t_R _32073_ (.A(_01927_),
    .B(_11242_),
    .Y(_12191_));
 AOI21x1_ASAP7_75t_R _32074_ (.A1(_01889_),
    .A2(_11226_),
    .B(_12191_),
    .Y(_04325_));
 AND2x2_ASAP7_75t_R _32075_ (.A(_01926_),
    .B(_11242_),
    .Y(_12192_));
 AOI21x1_ASAP7_75t_R _32076_ (.A1(_01888_),
    .A2(_11226_),
    .B(_12192_),
    .Y(_04326_));
 AND2x2_ASAP7_75t_R _32077_ (.A(_01925_),
    .B(_11242_),
    .Y(_12193_));
 AOI21x1_ASAP7_75t_R _32078_ (.A1(_01887_),
    .A2(_11226_),
    .B(_12193_),
    .Y(_04327_));
 AND2x2_ASAP7_75t_R _32079_ (.A(_01924_),
    .B(_11242_),
    .Y(_12194_));
 AOI21x1_ASAP7_75t_R _32080_ (.A1(_01886_),
    .A2(_11226_),
    .B(_12194_),
    .Y(_04328_));
 AND2x2_ASAP7_75t_R _32081_ (.A(_01923_),
    .B(_11242_),
    .Y(_12195_));
 AOI21x1_ASAP7_75t_R _32082_ (.A1(_01885_),
    .A2(_11226_),
    .B(_12195_),
    .Y(_04329_));
 AND2x2_ASAP7_75t_R _32083_ (.A(_01922_),
    .B(_11242_),
    .Y(_12196_));
 AOI21x1_ASAP7_75t_R _32084_ (.A1(_01884_),
    .A2(_11226_),
    .B(_12196_),
    .Y(_04330_));
 AND2x2_ASAP7_75t_R _32085_ (.A(_01921_),
    .B(_11242_),
    .Y(_12197_));
 AOI21x1_ASAP7_75t_R _32086_ (.A1(_01883_),
    .A2(_11226_),
    .B(_12197_),
    .Y(_04331_));
 AND2x2_ASAP7_75t_R _32087_ (.A(_01920_),
    .B(_11242_),
    .Y(_12198_));
 AOI21x1_ASAP7_75t_R _32088_ (.A1(_01882_),
    .A2(_11226_),
    .B(_12198_),
    .Y(_04332_));
 AND2x2_ASAP7_75t_R _32089_ (.A(_01919_),
    .B(_11242_),
    .Y(_12199_));
 AOI21x1_ASAP7_75t_R _32090_ (.A1(_01881_),
    .A2(_11226_),
    .B(_12199_),
    .Y(_04333_));
 AND2x2_ASAP7_75t_R _32091_ (.A(_01918_),
    .B(_11242_),
    .Y(_12200_));
 AOI21x1_ASAP7_75t_R _32092_ (.A1(_01880_),
    .A2(_11226_),
    .B(_12200_),
    .Y(_04334_));
 AND2x2_ASAP7_75t_R _32093_ (.A(_01917_),
    .B(_11242_),
    .Y(_12201_));
 AOI21x1_ASAP7_75t_R _32094_ (.A1(_01879_),
    .A2(_11226_),
    .B(_12201_),
    .Y(_04335_));
 AND2x2_ASAP7_75t_R _32095_ (.A(_01916_),
    .B(_11242_),
    .Y(_12202_));
 AOI21x1_ASAP7_75t_R _32096_ (.A1(_01878_),
    .A2(_11226_),
    .B(_12202_),
    .Y(_04336_));
 AND2x2_ASAP7_75t_R _32097_ (.A(_01915_),
    .B(_11242_),
    .Y(_12203_));
 AOI21x1_ASAP7_75t_R _32098_ (.A1(_01877_),
    .A2(_11226_),
    .B(_12203_),
    .Y(_04337_));
 NAND2x1_ASAP7_75t_R _32099_ (.A(_01876_),
    .B(_11226_),
    .Y(_12204_));
 OA21x2_ASAP7_75t_R _32100_ (.A1(_12137_),
    .A2(_11226_),
    .B(_12204_),
    .Y(_04338_));
 AND3x2_ASAP7_75t_R _32101_ (.A(_05580_),
    .B(_05538_),
    .C(_05582_),
    .Y(_12205_));
 NAND2x2_ASAP7_75t_R _32102_ (.A(_09365_),
    .B(_12205_),
    .Y(_12206_));
 NAND2x1_ASAP7_75t_R _32103_ (.A(_00661_),
    .B(_12206_),
    .Y(_12207_));
 OA21x2_ASAP7_75t_R _32104_ (.A1(_10974_),
    .A2(_12206_),
    .B(_12207_),
    .Y(_04339_));
 AO21x1_ASAP7_75t_R _32105_ (.A1(_09365_),
    .A2(_12205_),
    .B(_07380_),
    .Y(_12208_));
 OA21x2_ASAP7_75t_R _32106_ (.A1(_09390_),
    .A2(_12206_),
    .B(_12208_),
    .Y(_04340_));
 NAND2x1_ASAP7_75t_R _32107_ (.A(_01727_),
    .B(_05757_),
    .Y(_12209_));
 OA21x2_ASAP7_75t_R _32108_ (.A1(_13530_),
    .A2(_05757_),
    .B(_12209_),
    .Y(_04343_));
 NAND2x1_ASAP7_75t_R _32109_ (.A(_01873_),
    .B(_05747_),
    .Y(_12210_));
 OA21x2_ASAP7_75t_R _32110_ (.A1(_06705_),
    .A2(_05747_),
    .B(_12210_),
    .Y(_04344_));
 NAND2x1_ASAP7_75t_R _32111_ (.A(_01728_),
    .B(_05757_),
    .Y(_12211_));
 OA21x2_ASAP7_75t_R _32112_ (.A1(_05778_),
    .A2(_05757_),
    .B(_12211_),
    .Y(_04345_));
 AND3x4_ASAP7_75t_R _32113_ (.A(net59),
    .B(_01609_),
    .C(_13645_),
    .Y(_12212_));
 NAND2x2_ASAP7_75t_R _32114_ (.A(_01316_),
    .B(_12212_),
    .Y(_12213_));
 TAPCELL_ASAP7_75t_R PHY_125 ();
 TAPCELL_ASAP7_75t_R PHY_124 ();
 NAND2x1_ASAP7_75t_R _32117_ (.A(_01871_),
    .B(_12213_),
    .Y(_12216_));
 OA21x2_ASAP7_75t_R _32118_ (.A1(net57),
    .A2(_12213_),
    .B(_12216_),
    .Y(_04346_));
 TAPCELL_ASAP7_75t_R PHY_123 ();
 TAPCELL_ASAP7_75t_R PHY_122 ();
 AO21x1_ASAP7_75t_R _32121_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07188_),
    .Y(_12219_));
 OA21x2_ASAP7_75t_R _32122_ (.A1(net58),
    .A2(_12213_),
    .B(_12219_),
    .Y(_04347_));
 NAND2x1_ASAP7_75t_R _32123_ (.A(_01869_),
    .B(_12213_),
    .Y(_12220_));
 OA21x2_ASAP7_75t_R _32124_ (.A1(net28),
    .A2(_12213_),
    .B(_12220_),
    .Y(_04348_));
 NAND2x1_ASAP7_75t_R _32125_ (.A(_01868_),
    .B(_12213_),
    .Y(_12221_));
 OA21x2_ASAP7_75t_R _32126_ (.A1(net29),
    .A2(_12213_),
    .B(_12221_),
    .Y(_04349_));
 AO21x1_ASAP7_75t_R _32127_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07474_),
    .Y(_12222_));
 OA21x2_ASAP7_75t_R _32128_ (.A1(net30),
    .A2(_12213_),
    .B(_12222_),
    .Y(_04350_));
 AO21x1_ASAP7_75t_R _32129_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07538_),
    .Y(_12223_));
 OA21x2_ASAP7_75t_R _32130_ (.A1(net31),
    .A2(_12213_),
    .B(_12223_),
    .Y(_04351_));
 AO21x1_ASAP7_75t_R _32131_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07614_),
    .Y(_12224_));
 OA21x2_ASAP7_75t_R _32132_ (.A1(net32),
    .A2(_12213_),
    .B(_12224_),
    .Y(_04352_));
 AO21x1_ASAP7_75t_R _32133_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07624_),
    .Y(_12225_));
 OA21x2_ASAP7_75t_R _32134_ (.A1(net33),
    .A2(_12213_),
    .B(_12225_),
    .Y(_04353_));
 AO21x1_ASAP7_75t_R _32135_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07116_),
    .Y(_12226_));
 OA21x2_ASAP7_75t_R _32136_ (.A1(net34),
    .A2(_12213_),
    .B(_12226_),
    .Y(_04354_));
 AO21x1_ASAP7_75t_R _32137_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07187_),
    .Y(_12227_));
 OA21x2_ASAP7_75t_R _32138_ (.A1(net35),
    .A2(_12213_),
    .B(_12227_),
    .Y(_04355_));
 TAPCELL_ASAP7_75t_R PHY_121 ();
 TAPCELL_ASAP7_75t_R PHY_120 ();
 AO21x1_ASAP7_75t_R _32141_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07813_),
    .Y(_12230_));
 OA21x2_ASAP7_75t_R _32142_ (.A1(net36),
    .A2(_12213_),
    .B(_12230_),
    .Y(_04356_));
 AO21x1_ASAP7_75t_R _32143_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07861_),
    .Y(_12231_));
 OA21x2_ASAP7_75t_R _32144_ (.A1(net37),
    .A2(_12213_),
    .B(_12231_),
    .Y(_04357_));
 AO21x1_ASAP7_75t_R _32145_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07473_),
    .Y(_12232_));
 OA21x2_ASAP7_75t_R _32146_ (.A1(net39),
    .A2(_12213_),
    .B(_12232_),
    .Y(_04358_));
 AO21x1_ASAP7_75t_R _32147_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07537_),
    .Y(_12233_));
 OA21x2_ASAP7_75t_R _32148_ (.A1(net40),
    .A2(_12213_),
    .B(_12233_),
    .Y(_04359_));
 AO21x1_ASAP7_75t_R _32149_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07613_),
    .Y(_12234_));
 OA21x2_ASAP7_75t_R _32150_ (.A1(net41),
    .A2(_12213_),
    .B(_12234_),
    .Y(_04360_));
 AO21x1_ASAP7_75t_R _32151_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07623_),
    .Y(_12235_));
 OA21x2_ASAP7_75t_R _32152_ (.A1(net42),
    .A2(_12213_),
    .B(_12235_),
    .Y(_04361_));
 AO21x1_ASAP7_75t_R _32153_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07718_),
    .Y(_12236_));
 OA21x2_ASAP7_75t_R _32154_ (.A1(net43),
    .A2(_12213_),
    .B(_12236_),
    .Y(_04362_));
 NAND2x1_ASAP7_75t_R _32155_ (.A(_01854_),
    .B(_12213_),
    .Y(_12237_));
 OA21x2_ASAP7_75t_R _32156_ (.A1(net44),
    .A2(_12213_),
    .B(_12237_),
    .Y(_04363_));
 AO21x1_ASAP7_75t_R _32157_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07811_),
    .Y(_12238_));
 OA21x2_ASAP7_75t_R _32158_ (.A1(net45),
    .A2(_12213_),
    .B(_12238_),
    .Y(_04364_));
 AO21x1_ASAP7_75t_R _32159_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07859_),
    .Y(_12239_));
 OA21x2_ASAP7_75t_R _32160_ (.A1(net46),
    .A2(_12213_),
    .B(_12239_),
    .Y(_04365_));
 AO21x1_ASAP7_75t_R _32161_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07903_),
    .Y(_12240_));
 OA21x2_ASAP7_75t_R _32162_ (.A1(net47),
    .A2(_12213_),
    .B(_12240_),
    .Y(_04366_));
 AO21x1_ASAP7_75t_R _32163_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07945_),
    .Y(_12241_));
 OA21x2_ASAP7_75t_R _32164_ (.A1(net48),
    .A2(_12213_),
    .B(_12241_),
    .Y(_04367_));
 AO21x1_ASAP7_75t_R _32165_ (.A1(_01316_),
    .A2(_12212_),
    .B(_07985_),
    .Y(_12242_));
 OA21x2_ASAP7_75t_R _32166_ (.A1(net50),
    .A2(_12213_),
    .B(_12242_),
    .Y(_04368_));
 NAND2x1_ASAP7_75t_R _32167_ (.A(_01733_),
    .B(_12213_),
    .Y(_12243_));
 OA21x2_ASAP7_75t_R _32168_ (.A1(net51),
    .A2(_12213_),
    .B(_12243_),
    .Y(_04369_));
 XNOR2x1_ASAP7_75t_R _32169_ (.B(_06666_),
    .Y(_12244_),
    .A(_06537_));
 OR3x2_ASAP7_75t_R _32170_ (.A(_06670_),
    .B(_06680_),
    .C(_12244_),
    .Y(_12245_));
 NAND2x1_ASAP7_75t_R _32171_ (.A(_01813_),
    .B(_06680_),
    .Y(_12246_));
 OR4x2_ASAP7_75t_R _32172_ (.A(_00239_),
    .B(_06655_),
    .C(_06656_),
    .D(_06665_),
    .Y(_12247_));
 TAPCELL_ASAP7_75t_R PHY_119 ();
 NAND2x1_ASAP7_75t_R _32174_ (.A(_01846_),
    .B(_12247_),
    .Y(_12249_));
 TAPCELL_ASAP7_75t_R PHY_118 ();
 TAPCELL_ASAP7_75t_R PHY_117 ();
 TAPCELL_ASAP7_75t_R PHY_116 ();
 NOR2x1_ASAP7_75t_R _32178_ (.A(_00239_),
    .B(_01813_),
    .Y(_12253_));
 AO31x2_ASAP7_75t_R _32179_ (.A1(net96),
    .A2(_00239_),
    .A3(_06666_),
    .B(_12253_),
    .Y(_12254_));
 INVx1_ASAP7_75t_R _32180_ (.A(_06665_),
    .Y(_12255_));
 AND4x2_ASAP7_75t_R _32181_ (.A(_06537_),
    .B(_00239_),
    .C(_06607_),
    .D(_12255_),
    .Y(_12256_));
 AO22x1_ASAP7_75t_R _32182_ (.A1(_00240_),
    .A2(_12254_),
    .B1(_12256_),
    .B2(net96),
    .Y(_12257_));
 AO32x1_ASAP7_75t_R _32183_ (.A1(_12245_),
    .A2(_12246_),
    .A3(_12249_),
    .B1(_12257_),
    .B2(_06617_),
    .Y(_04371_));
 XNOR2x1_ASAP7_75t_R _32184_ (.B(_06666_),
    .Y(_12258_),
    .A(_00240_));
 AND3x4_ASAP7_75t_R _32185_ (.A(_00239_),
    .B(_06617_),
    .C(_12258_),
    .Y(_12259_));
 TAPCELL_ASAP7_75t_R PHY_115 ();
 TAPCELL_ASAP7_75t_R PHY_114 ();
 OA21x2_ASAP7_75t_R _32188_ (.A1(_06537_),
    .A2(_06670_),
    .B(_06666_),
    .Y(_12262_));
 NOR2x2_ASAP7_75t_R _32189_ (.A(_00239_),
    .B(_12262_),
    .Y(_12263_));
 TAPCELL_ASAP7_75t_R PHY_113 ();
 INVx1_ASAP7_75t_R _32191_ (.A(_01812_),
    .Y(_12265_));
 INVx1_ASAP7_75t_R _32192_ (.A(_01845_),
    .Y(_12266_));
 OA21x2_ASAP7_75t_R _32193_ (.A1(_06670_),
    .A2(_12244_),
    .B(_12247_),
    .Y(_12267_));
 TAPCELL_ASAP7_75t_R PHY_112 ();
 AO222x2_ASAP7_75t_R _32195_ (.A1(net107),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12265_),
    .C1(_12266_),
    .C2(_12267_),
    .Y(_04372_));
 INVx1_ASAP7_75t_R _32196_ (.A(_01811_),
    .Y(_12269_));
 INVx1_ASAP7_75t_R _32197_ (.A(_01844_),
    .Y(_12270_));
 AO222x2_ASAP7_75t_R _32198_ (.A1(net118),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12269_),
    .C1(_12270_),
    .C2(_12267_),
    .Y(_04373_));
 NAND2x1_ASAP7_75t_R _32199_ (.A(_01810_),
    .B(_06680_),
    .Y(_12271_));
 NAND2x1_ASAP7_75t_R _32200_ (.A(_01843_),
    .B(_12247_),
    .Y(_12272_));
 NOR2x1_ASAP7_75t_R _32201_ (.A(_00239_),
    .B(_01810_),
    .Y(_12273_));
 AO31x2_ASAP7_75t_R _32202_ (.A1(net121),
    .A2(_00239_),
    .A3(_06666_),
    .B(_12273_),
    .Y(_12274_));
 AO22x1_ASAP7_75t_R _32203_ (.A1(net121),
    .A2(_12256_),
    .B1(_12274_),
    .B2(_00240_),
    .Y(_12275_));
 AO32x1_ASAP7_75t_R _32204_ (.A1(_12245_),
    .A2(_12271_),
    .A3(_12272_),
    .B1(_12275_),
    .B2(_06617_),
    .Y(_04374_));
 INVx1_ASAP7_75t_R _32205_ (.A(_01809_),
    .Y(_12276_));
 INVx1_ASAP7_75t_R _32206_ (.A(_01842_),
    .Y(_12277_));
 AO222x2_ASAP7_75t_R _32207_ (.A1(net122),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12276_),
    .C1(_12277_),
    .C2(_12267_),
    .Y(_04375_));
 INVx1_ASAP7_75t_R _32208_ (.A(_01808_),
    .Y(_12278_));
 INVx1_ASAP7_75t_R _32209_ (.A(_01841_),
    .Y(_12279_));
 AO222x2_ASAP7_75t_R _32210_ (.A1(net123),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12278_),
    .C1(_12279_),
    .C2(_12267_),
    .Y(_04376_));
 NAND2x1_ASAP7_75t_R _32211_ (.A(_01807_),
    .B(_06680_),
    .Y(_12280_));
 NAND2x1_ASAP7_75t_R _32212_ (.A(_01840_),
    .B(_12247_),
    .Y(_12281_));
 NOR2x1_ASAP7_75t_R _32213_ (.A(_00239_),
    .B(_01807_),
    .Y(_12282_));
 AO31x2_ASAP7_75t_R _32214_ (.A1(net124),
    .A2(_00239_),
    .A3(_06666_),
    .B(_12282_),
    .Y(_12283_));
 AO22x1_ASAP7_75t_R _32215_ (.A1(net124),
    .A2(_12256_),
    .B1(_12283_),
    .B2(_00240_),
    .Y(_12284_));
 AO32x1_ASAP7_75t_R _32216_ (.A1(_12245_),
    .A2(_12280_),
    .A3(_12281_),
    .B1(_12284_),
    .B2(_06617_),
    .Y(_04377_));
 INVx1_ASAP7_75t_R _32217_ (.A(_01806_),
    .Y(_12285_));
 INVx1_ASAP7_75t_R _32218_ (.A(_01839_),
    .Y(_12286_));
 AO222x2_ASAP7_75t_R _32219_ (.A1(net125),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12285_),
    .C1(_12286_),
    .C2(_12267_),
    .Y(_04378_));
 INVx1_ASAP7_75t_R _32220_ (.A(_01805_),
    .Y(_12287_));
 INVx1_ASAP7_75t_R _32221_ (.A(_01838_),
    .Y(_12288_));
 AO222x2_ASAP7_75t_R _32222_ (.A1(net126),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12287_),
    .C1(_12288_),
    .C2(_12267_),
    .Y(_04379_));
 INVx1_ASAP7_75t_R _32223_ (.A(_01804_),
    .Y(_12289_));
 INVx1_ASAP7_75t_R _32224_ (.A(_01837_),
    .Y(_12290_));
 AO222x2_ASAP7_75t_R _32225_ (.A1(net127),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12289_),
    .C1(_12290_),
    .C2(_12267_),
    .Y(_04380_));
 NAND2x1_ASAP7_75t_R _32226_ (.A(_01803_),
    .B(_06680_),
    .Y(_12291_));
 NAND2x1_ASAP7_75t_R _32227_ (.A(_01836_),
    .B(_12247_),
    .Y(_12292_));
 NOR2x1_ASAP7_75t_R _32228_ (.A(_00239_),
    .B(_01803_),
    .Y(_12293_));
 AO31x2_ASAP7_75t_R _32229_ (.A1(net97),
    .A2(_00239_),
    .A3(_06666_),
    .B(_12293_),
    .Y(_12294_));
 AO22x1_ASAP7_75t_R _32230_ (.A1(net97),
    .A2(_12256_),
    .B1(_12294_),
    .B2(_00240_),
    .Y(_12295_));
 AO32x1_ASAP7_75t_R _32231_ (.A1(_12245_),
    .A2(_12291_),
    .A3(_12292_),
    .B1(_12295_),
    .B2(_06617_),
    .Y(_04381_));
 INVx1_ASAP7_75t_R _32232_ (.A(_01802_),
    .Y(_12296_));
 INVx1_ASAP7_75t_R _32233_ (.A(_01835_),
    .Y(_12297_));
 AO222x2_ASAP7_75t_R _32234_ (.A1(net98),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12296_),
    .C1(_12297_),
    .C2(_12267_),
    .Y(_04382_));
 INVx1_ASAP7_75t_R _32235_ (.A(_01801_),
    .Y(_12298_));
 INVx1_ASAP7_75t_R _32236_ (.A(_01834_),
    .Y(_12299_));
 AO222x2_ASAP7_75t_R _32237_ (.A1(net99),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12298_),
    .C1(_12299_),
    .C2(_12267_),
    .Y(_04383_));
 TAPCELL_ASAP7_75t_R PHY_111 ();
 INVx1_ASAP7_75t_R _32239_ (.A(_01800_),
    .Y(_12301_));
 INVx1_ASAP7_75t_R _32240_ (.A(_01833_),
    .Y(_12302_));
 TAPCELL_ASAP7_75t_R PHY_110 ();
 TAPCELL_ASAP7_75t_R PHY_109 ();
 AO222x2_ASAP7_75t_R _32243_ (.A1(net100),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12301_),
    .C1(_12302_),
    .C2(_12267_),
    .Y(_04384_));
 TAPCELL_ASAP7_75t_R PHY_108 ();
 INVx1_ASAP7_75t_R _32245_ (.A(_01799_),
    .Y(_12306_));
 INVx1_ASAP7_75t_R _32246_ (.A(_01832_),
    .Y(_12307_));
 AO222x2_ASAP7_75t_R _32247_ (.A1(net101),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12306_),
    .C1(_12307_),
    .C2(_12267_),
    .Y(_04385_));
 INVx1_ASAP7_75t_R _32248_ (.A(_01798_),
    .Y(_12308_));
 INVx1_ASAP7_75t_R _32249_ (.A(_01831_),
    .Y(_12309_));
 AO222x2_ASAP7_75t_R _32250_ (.A1(net102),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12308_),
    .C1(_12309_),
    .C2(_12267_),
    .Y(_04386_));
 INVx1_ASAP7_75t_R _32251_ (.A(_01797_),
    .Y(_12310_));
 INVx1_ASAP7_75t_R _32252_ (.A(_01830_),
    .Y(_12311_));
 AO222x2_ASAP7_75t_R _32253_ (.A1(net103),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12310_),
    .C1(_12311_),
    .C2(_12267_),
    .Y(_04387_));
 INVx1_ASAP7_75t_R _32254_ (.A(_01796_),
    .Y(_12312_));
 INVx1_ASAP7_75t_R _32255_ (.A(_01829_),
    .Y(_12313_));
 AO222x2_ASAP7_75t_R _32256_ (.A1(net104),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12312_),
    .C1(_12313_),
    .C2(_12267_),
    .Y(_04388_));
 INVx1_ASAP7_75t_R _32257_ (.A(_01795_),
    .Y(_12314_));
 INVx1_ASAP7_75t_R _32258_ (.A(_01828_),
    .Y(_12315_));
 AO222x2_ASAP7_75t_R _32259_ (.A1(net105),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12314_),
    .C1(_12315_),
    .C2(_12267_),
    .Y(_04389_));
 INVx1_ASAP7_75t_R _32260_ (.A(_01794_),
    .Y(_12316_));
 INVx1_ASAP7_75t_R _32261_ (.A(_01827_),
    .Y(_12317_));
 AO222x2_ASAP7_75t_R _32262_ (.A1(net106),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12316_),
    .C1(_12317_),
    .C2(_12267_),
    .Y(_04390_));
 INVx1_ASAP7_75t_R _32263_ (.A(_01793_),
    .Y(_12318_));
 INVx1_ASAP7_75t_R _32264_ (.A(_01826_),
    .Y(_12319_));
 AO222x2_ASAP7_75t_R _32265_ (.A1(net108),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12318_),
    .C1(_12319_),
    .C2(_12267_),
    .Y(_04391_));
 INVx1_ASAP7_75t_R _32266_ (.A(_01792_),
    .Y(_12320_));
 INVx1_ASAP7_75t_R _32267_ (.A(_01825_),
    .Y(_12321_));
 AO222x2_ASAP7_75t_R _32268_ (.A1(net109),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12320_),
    .C1(_12321_),
    .C2(_12267_),
    .Y(_04392_));
 INVx1_ASAP7_75t_R _32269_ (.A(_01791_),
    .Y(_12322_));
 INVx1_ASAP7_75t_R _32270_ (.A(_01824_),
    .Y(_12323_));
 AO222x2_ASAP7_75t_R _32271_ (.A1(net110),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12322_),
    .C1(_12323_),
    .C2(_12267_),
    .Y(_04393_));
 INVx1_ASAP7_75t_R _32272_ (.A(_01790_),
    .Y(_12324_));
 INVx1_ASAP7_75t_R _32273_ (.A(_01823_),
    .Y(_12325_));
 AO222x2_ASAP7_75t_R _32274_ (.A1(net111),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12324_),
    .C1(_12325_),
    .C2(_12267_),
    .Y(_04394_));
 INVx1_ASAP7_75t_R _32275_ (.A(_01789_),
    .Y(_12326_));
 INVx1_ASAP7_75t_R _32276_ (.A(_01822_),
    .Y(_12327_));
 AO222x2_ASAP7_75t_R _32277_ (.A1(net112),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12326_),
    .C1(_12327_),
    .C2(_12267_),
    .Y(_04395_));
 INVx1_ASAP7_75t_R _32278_ (.A(_01788_),
    .Y(_12328_));
 INVx1_ASAP7_75t_R _32279_ (.A(_01821_),
    .Y(_12329_));
 AO222x2_ASAP7_75t_R _32280_ (.A1(net113),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12328_),
    .C1(_12329_),
    .C2(_12267_),
    .Y(_04396_));
 INVx1_ASAP7_75t_R _32281_ (.A(_01787_),
    .Y(_12330_));
 INVx1_ASAP7_75t_R _32282_ (.A(_01820_),
    .Y(_12331_));
 AO222x2_ASAP7_75t_R _32283_ (.A1(net114),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12330_),
    .C1(_12331_),
    .C2(_12267_),
    .Y(_04397_));
 INVx1_ASAP7_75t_R _32284_ (.A(_01786_),
    .Y(_12332_));
 INVx1_ASAP7_75t_R _32285_ (.A(_01819_),
    .Y(_12333_));
 AO222x2_ASAP7_75t_R _32286_ (.A1(net115),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12332_),
    .C1(_12333_),
    .C2(_12267_),
    .Y(_04398_));
 INVx1_ASAP7_75t_R _32287_ (.A(_01785_),
    .Y(_12334_));
 INVx1_ASAP7_75t_R _32288_ (.A(_01818_),
    .Y(_12335_));
 AO222x2_ASAP7_75t_R _32289_ (.A1(net116),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12334_),
    .C1(_12335_),
    .C2(_12267_),
    .Y(_04399_));
 INVx1_ASAP7_75t_R _32290_ (.A(_01784_),
    .Y(_12336_));
 INVx1_ASAP7_75t_R _32291_ (.A(_01817_),
    .Y(_12337_));
 AO222x2_ASAP7_75t_R _32292_ (.A1(net117),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12336_),
    .C1(_12337_),
    .C2(_12267_),
    .Y(_04400_));
 INVx1_ASAP7_75t_R _32293_ (.A(_01783_),
    .Y(_12338_));
 INVx1_ASAP7_75t_R _32294_ (.A(_01816_),
    .Y(_12339_));
 AO222x2_ASAP7_75t_R _32295_ (.A1(net119),
    .A2(_12259_),
    .B1(_12263_),
    .B2(_12338_),
    .C1(_12339_),
    .C2(_12267_),
    .Y(_04401_));
 INVx1_ASAP7_75t_R _32296_ (.A(_01738_),
    .Y(_12340_));
 INVx1_ASAP7_75t_R _32297_ (.A(_01782_),
    .Y(_12341_));
 AO222x2_ASAP7_75t_R _32298_ (.A1(_12340_),
    .A2(_12267_),
    .B1(_12263_),
    .B2(_12341_),
    .C1(_12259_),
    .C2(net120),
    .Y(_04402_));
 AND2x2_ASAP7_75t_R _32299_ (.A(_00239_),
    .B(_06538_),
    .Y(_12342_));
 AO21x1_ASAP7_75t_R _32300_ (.A1(_06511_),
    .A2(_01781_),
    .B(_12342_),
    .Y(_12343_));
 AO211x2_ASAP7_75t_R _32301_ (.A1(_06617_),
    .A2(_12258_),
    .B(_06680_),
    .C(_01814_),
    .Y(_12344_));
 OAI21x1_ASAP7_75t_R _32302_ (.A1(_12267_),
    .A2(_12343_),
    .B(_12344_),
    .Y(_04403_));
 NAND2x1_ASAP7_75t_R _32303_ (.A(_06537_),
    .B(_00239_),
    .Y(_12345_));
 AO31x2_ASAP7_75t_R _32304_ (.A1(_06558_),
    .A2(_06606_),
    .A3(_12255_),
    .B(_12345_),
    .Y(_12346_));
 AO21x2_ASAP7_75t_R _32305_ (.A1(_12247_),
    .A2(_12346_),
    .B(_06670_),
    .Y(_12347_));
 NAND2x2_ASAP7_75t_R _32306_ (.A(_06674_),
    .B(_12347_),
    .Y(_12348_));
 TAPCELL_ASAP7_75t_R PHY_107 ();
 TAPCELL_ASAP7_75t_R PHY_106 ();
 TAPCELL_ASAP7_75t_R PHY_105 ();
 TAPCELL_ASAP7_75t_R PHY_104 ();
 TAPCELL_ASAP7_75t_R PHY_103 ();
 NAND2x1_ASAP7_75t_R _32312_ (.A(net96),
    .B(net413),
    .Y(_12354_));
 OA21x2_ASAP7_75t_R _32313_ (.A1(net413),
    .A2(_01780_),
    .B(_12354_),
    .Y(_12355_));
 AO21x1_ASAP7_75t_R _32314_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12355_),
    .Y(_12356_));
 OAI21x1_ASAP7_75t_R _32315_ (.A1(_01813_),
    .A2(_12348_),
    .B(_12356_),
    .Y(_04404_));
 NAND2x1_ASAP7_75t_R _32316_ (.A(net107),
    .B(_01815_),
    .Y(_12357_));
 OA21x2_ASAP7_75t_R _32317_ (.A1(_01815_),
    .A2(_01779_),
    .B(_12357_),
    .Y(_12358_));
 AO21x1_ASAP7_75t_R _32318_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12358_),
    .Y(_12359_));
 OAI21x1_ASAP7_75t_R _32319_ (.A1(_01812_),
    .A2(_12348_),
    .B(_12359_),
    .Y(_04405_));
 NAND2x1_ASAP7_75t_R _32320_ (.A(net118),
    .B(_01815_),
    .Y(_12360_));
 OA21x2_ASAP7_75t_R _32321_ (.A1(_01815_),
    .A2(_01778_),
    .B(_12360_),
    .Y(_12361_));
 AO21x1_ASAP7_75t_R _32322_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12361_),
    .Y(_12362_));
 OAI21x1_ASAP7_75t_R _32323_ (.A1(_01811_),
    .A2(_12348_),
    .B(_12362_),
    .Y(_04406_));
 NAND2x1_ASAP7_75t_R _32324_ (.A(net121),
    .B(net413),
    .Y(_12363_));
 OA21x2_ASAP7_75t_R _32325_ (.A1(net413),
    .A2(_01777_),
    .B(_12363_),
    .Y(_12364_));
 AO21x1_ASAP7_75t_R _32326_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12364_),
    .Y(_12365_));
 OAI21x1_ASAP7_75t_R _32327_ (.A1(_01810_),
    .A2(_12348_),
    .B(_12365_),
    .Y(_04407_));
 NAND2x1_ASAP7_75t_R _32328_ (.A(net122),
    .B(net413),
    .Y(_12366_));
 OA21x2_ASAP7_75t_R _32329_ (.A1(net413),
    .A2(_01776_),
    .B(_12366_),
    .Y(_12367_));
 AO21x1_ASAP7_75t_R _32330_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12367_),
    .Y(_12368_));
 OAI21x1_ASAP7_75t_R _32331_ (.A1(_01809_),
    .A2(_12348_),
    .B(_12368_),
    .Y(_04408_));
 NAND2x1_ASAP7_75t_R _32332_ (.A(net123),
    .B(_01815_),
    .Y(_12369_));
 OA21x2_ASAP7_75t_R _32333_ (.A1(_01815_),
    .A2(_01775_),
    .B(_12369_),
    .Y(_12370_));
 AO21x1_ASAP7_75t_R _32334_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12370_),
    .Y(_12371_));
 OAI21x1_ASAP7_75t_R _32335_ (.A1(_01808_),
    .A2(_12348_),
    .B(_12371_),
    .Y(_04409_));
 TAPCELL_ASAP7_75t_R PHY_102 ();
 NAND2x1_ASAP7_75t_R _32337_ (.A(net124),
    .B(net413),
    .Y(_12373_));
 OA21x2_ASAP7_75t_R _32338_ (.A1(net413),
    .A2(_01774_),
    .B(_12373_),
    .Y(_12374_));
 AO21x1_ASAP7_75t_R _32339_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12374_),
    .Y(_12375_));
 OAI21x1_ASAP7_75t_R _32340_ (.A1(_01807_),
    .A2(_12348_),
    .B(_12375_),
    .Y(_04410_));
 NOR2x1_ASAP7_75t_R _32341_ (.A(net413),
    .B(_01773_),
    .Y(_12376_));
 AO21x1_ASAP7_75t_R _32342_ (.A1(net125),
    .A2(net413),
    .B(_12376_),
    .Y(_12377_));
 AND3x1_ASAP7_75t_R _32343_ (.A(_12285_),
    .B(_06674_),
    .C(_12347_),
    .Y(_12378_));
 AO21x1_ASAP7_75t_R _32344_ (.A1(_12348_),
    .A2(_12377_),
    .B(_12378_),
    .Y(_04411_));
 NAND2x1_ASAP7_75t_R _32345_ (.A(net126),
    .B(_01815_),
    .Y(_12379_));
 OA21x2_ASAP7_75t_R _32346_ (.A1(_01815_),
    .A2(_01772_),
    .B(_12379_),
    .Y(_12380_));
 AO21x1_ASAP7_75t_R _32347_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12380_),
    .Y(_12381_));
 OAI21x1_ASAP7_75t_R _32348_ (.A1(_01805_),
    .A2(_12348_),
    .B(_12381_),
    .Y(_04412_));
 NAND2x1_ASAP7_75t_R _32349_ (.A(net127),
    .B(net413),
    .Y(_12382_));
 OA21x2_ASAP7_75t_R _32350_ (.A1(net413),
    .A2(_01771_),
    .B(_12382_),
    .Y(_12383_));
 AO21x1_ASAP7_75t_R _32351_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12383_),
    .Y(_12384_));
 OAI21x1_ASAP7_75t_R _32352_ (.A1(_01804_),
    .A2(_12348_),
    .B(_12384_),
    .Y(_04413_));
 TAPCELL_ASAP7_75t_R PHY_101 ();
 TAPCELL_ASAP7_75t_R PHY_100 ();
 NAND2x1_ASAP7_75t_R _32355_ (.A(net97),
    .B(net413),
    .Y(_12387_));
 OA21x2_ASAP7_75t_R _32356_ (.A1(net413),
    .A2(_01770_),
    .B(_12387_),
    .Y(_12388_));
 AO21x1_ASAP7_75t_R _32357_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12388_),
    .Y(_12389_));
 OAI21x1_ASAP7_75t_R _32358_ (.A1(_01803_),
    .A2(_12348_),
    .B(_12389_),
    .Y(_04414_));
 TAPCELL_ASAP7_75t_R PHY_99 ();
 TAPCELL_ASAP7_75t_R PHY_98 ();
 NAND2x1_ASAP7_75t_R _32361_ (.A(net98),
    .B(net413),
    .Y(_12392_));
 OA21x2_ASAP7_75t_R _32362_ (.A1(net413),
    .A2(_01769_),
    .B(_12392_),
    .Y(_12393_));
 AO21x1_ASAP7_75t_R _32363_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12393_),
    .Y(_12394_));
 OAI21x1_ASAP7_75t_R _32364_ (.A1(_01802_),
    .A2(_12348_),
    .B(_12394_),
    .Y(_04415_));
 NAND2x1_ASAP7_75t_R _32365_ (.A(net99),
    .B(_01815_),
    .Y(_12395_));
 OA21x2_ASAP7_75t_R _32366_ (.A1(_01815_),
    .A2(_01768_),
    .B(_12395_),
    .Y(_12396_));
 AO21x1_ASAP7_75t_R _32367_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12396_),
    .Y(_12397_));
 OAI21x1_ASAP7_75t_R _32368_ (.A1(_01801_),
    .A2(_12348_),
    .B(_12397_),
    .Y(_04416_));
 NAND2x1_ASAP7_75t_R _32369_ (.A(net100),
    .B(_01815_),
    .Y(_12398_));
 OA21x2_ASAP7_75t_R _32370_ (.A1(_01815_),
    .A2(_01767_),
    .B(_12398_),
    .Y(_12399_));
 AO21x1_ASAP7_75t_R _32371_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12399_),
    .Y(_12400_));
 OAI21x1_ASAP7_75t_R _32372_ (.A1(_01800_),
    .A2(_12348_),
    .B(_12400_),
    .Y(_04417_));
 NAND2x1_ASAP7_75t_R _32373_ (.A(net101),
    .B(net413),
    .Y(_12401_));
 OA21x2_ASAP7_75t_R _32374_ (.A1(net413),
    .A2(_01766_),
    .B(_12401_),
    .Y(_12402_));
 AO21x1_ASAP7_75t_R _32375_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12402_),
    .Y(_12403_));
 OAI21x1_ASAP7_75t_R _32376_ (.A1(_01799_),
    .A2(_12348_),
    .B(_12403_),
    .Y(_04418_));
 NAND2x1_ASAP7_75t_R _32377_ (.A(net102),
    .B(_01815_),
    .Y(_12404_));
 OA21x2_ASAP7_75t_R _32378_ (.A1(_01815_),
    .A2(_01765_),
    .B(_12404_),
    .Y(_12405_));
 AO21x1_ASAP7_75t_R _32379_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12405_),
    .Y(_12406_));
 OAI21x1_ASAP7_75t_R _32380_ (.A1(_01798_),
    .A2(_12348_),
    .B(_12406_),
    .Y(_04419_));
 AND2x2_ASAP7_75t_R _32381_ (.A(_06532_),
    .B(_01815_),
    .Y(_12407_));
 AO221x1_ASAP7_75t_R _32382_ (.A1(_06509_),
    .A2(_01764_),
    .B1(_06674_),
    .B2(_12347_),
    .C(_12407_),
    .Y(_12408_));
 OAI21x1_ASAP7_75t_R _32383_ (.A1(_01797_),
    .A2(_12348_),
    .B(_12408_),
    .Y(_04420_));
 NAND2x1_ASAP7_75t_R _32384_ (.A(net104),
    .B(_01815_),
    .Y(_12409_));
 OA21x2_ASAP7_75t_R _32385_ (.A1(_01815_),
    .A2(_01763_),
    .B(_12409_),
    .Y(_12410_));
 AO21x1_ASAP7_75t_R _32386_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12410_),
    .Y(_12411_));
 OAI21x1_ASAP7_75t_R _32387_ (.A1(_01796_),
    .A2(_12348_),
    .B(_12411_),
    .Y(_04421_));
 TAPCELL_ASAP7_75t_R PHY_97 ();
 NAND2x1_ASAP7_75t_R _32389_ (.A(net105),
    .B(_01815_),
    .Y(_12413_));
 OA21x2_ASAP7_75t_R _32390_ (.A1(_01815_),
    .A2(_01762_),
    .B(_12413_),
    .Y(_12414_));
 AO21x1_ASAP7_75t_R _32391_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12414_),
    .Y(_12415_));
 OAI21x1_ASAP7_75t_R _32392_ (.A1(_01795_),
    .A2(_12348_),
    .B(_12415_),
    .Y(_04422_));
 NAND2x1_ASAP7_75t_R _32393_ (.A(net106),
    .B(net413),
    .Y(_12416_));
 OA21x2_ASAP7_75t_R _32394_ (.A1(net413),
    .A2(_01761_),
    .B(_12416_),
    .Y(_12417_));
 AO21x1_ASAP7_75t_R _32395_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12417_),
    .Y(_12418_));
 OAI21x1_ASAP7_75t_R _32396_ (.A1(_01794_),
    .A2(_12348_),
    .B(_12418_),
    .Y(_04423_));
 NAND2x1_ASAP7_75t_R _32397_ (.A(net108),
    .B(net413),
    .Y(_12419_));
 OA21x2_ASAP7_75t_R _32398_ (.A1(net413),
    .A2(_01760_),
    .B(_12419_),
    .Y(_12420_));
 AO21x1_ASAP7_75t_R _32399_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12420_),
    .Y(_12421_));
 OAI21x1_ASAP7_75t_R _32400_ (.A1(_01793_),
    .A2(_12348_),
    .B(_12421_),
    .Y(_04424_));
 TAPCELL_ASAP7_75t_R PHY_96 ();
 TAPCELL_ASAP7_75t_R PHY_95 ();
 TAPCELL_ASAP7_75t_R PHY_94 ();
 NAND2x1_ASAP7_75t_R _32404_ (.A(net109),
    .B(_01815_),
    .Y(_12425_));
 OA21x2_ASAP7_75t_R _32405_ (.A1(_01815_),
    .A2(_01759_),
    .B(_12425_),
    .Y(_12426_));
 AO21x1_ASAP7_75t_R _32406_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12426_),
    .Y(_12427_));
 OAI21x1_ASAP7_75t_R _32407_ (.A1(_01792_),
    .A2(_12348_),
    .B(_12427_),
    .Y(_04425_));
 TAPCELL_ASAP7_75t_R PHY_93 ();
 NAND2x1_ASAP7_75t_R _32409_ (.A(net110),
    .B(net413),
    .Y(_12429_));
 OA21x2_ASAP7_75t_R _32410_ (.A1(net413),
    .A2(_01758_),
    .B(_12429_),
    .Y(_12430_));
 AO21x1_ASAP7_75t_R _32411_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12430_),
    .Y(_12431_));
 OAI21x1_ASAP7_75t_R _32412_ (.A1(_01791_),
    .A2(_12348_),
    .B(_12431_),
    .Y(_04426_));
 NAND2x1_ASAP7_75t_R _32413_ (.A(net111),
    .B(net413),
    .Y(_12432_));
 OA21x2_ASAP7_75t_R _32414_ (.A1(net413),
    .A2(_01757_),
    .B(_12432_),
    .Y(_12433_));
 AO21x1_ASAP7_75t_R _32415_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12433_),
    .Y(_12434_));
 OAI21x1_ASAP7_75t_R _32416_ (.A1(_01790_),
    .A2(_12348_),
    .B(_12434_),
    .Y(_04427_));
 NAND2x1_ASAP7_75t_R _32417_ (.A(net112),
    .B(net413),
    .Y(_12435_));
 OA21x2_ASAP7_75t_R _32418_ (.A1(net413),
    .A2(_01756_),
    .B(_12435_),
    .Y(_12436_));
 AO21x1_ASAP7_75t_R _32419_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12436_),
    .Y(_12437_));
 OAI21x1_ASAP7_75t_R _32420_ (.A1(_01789_),
    .A2(_12348_),
    .B(_12437_),
    .Y(_04428_));
 NAND2x1_ASAP7_75t_R _32421_ (.A(net113),
    .B(net413),
    .Y(_12438_));
 OA21x2_ASAP7_75t_R _32422_ (.A1(net413),
    .A2(_01755_),
    .B(_12438_),
    .Y(_12439_));
 AO21x1_ASAP7_75t_R _32423_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12439_),
    .Y(_12440_));
 OAI21x1_ASAP7_75t_R _32424_ (.A1(_01788_),
    .A2(_12348_),
    .B(_12440_),
    .Y(_04429_));
 NAND2x1_ASAP7_75t_R _32425_ (.A(net114),
    .B(net413),
    .Y(_12441_));
 OA21x2_ASAP7_75t_R _32426_ (.A1(net413),
    .A2(_01754_),
    .B(_12441_),
    .Y(_12442_));
 AO21x1_ASAP7_75t_R _32427_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12442_),
    .Y(_12443_));
 OAI21x1_ASAP7_75t_R _32428_ (.A1(_01787_),
    .A2(_12348_),
    .B(_12443_),
    .Y(_04430_));
 NAND2x1_ASAP7_75t_R _32429_ (.A(net115),
    .B(net413),
    .Y(_12444_));
 OA21x2_ASAP7_75t_R _32430_ (.A1(net413),
    .A2(_01753_),
    .B(_12444_),
    .Y(_12445_));
 AO21x1_ASAP7_75t_R _32431_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12445_),
    .Y(_12446_));
 OAI21x1_ASAP7_75t_R _32432_ (.A1(_01786_),
    .A2(_12348_),
    .B(_12446_),
    .Y(_04431_));
 NAND2x1_ASAP7_75t_R _32433_ (.A(net116),
    .B(_01815_),
    .Y(_12447_));
 OA21x2_ASAP7_75t_R _32434_ (.A1(_01815_),
    .A2(_01752_),
    .B(_12447_),
    .Y(_12448_));
 AO21x1_ASAP7_75t_R _32435_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12448_),
    .Y(_12449_));
 OAI21x1_ASAP7_75t_R _32436_ (.A1(_01785_),
    .A2(_12348_),
    .B(_12449_),
    .Y(_04432_));
 NAND2x1_ASAP7_75t_R _32437_ (.A(net117),
    .B(_01815_),
    .Y(_12450_));
 OA21x2_ASAP7_75t_R _32438_ (.A1(_01815_),
    .A2(_01751_),
    .B(_12450_),
    .Y(_12451_));
 AO21x1_ASAP7_75t_R _32439_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12451_),
    .Y(_12452_));
 OAI21x1_ASAP7_75t_R _32440_ (.A1(_01784_),
    .A2(_12348_),
    .B(_12452_),
    .Y(_04433_));
 NAND2x1_ASAP7_75t_R _32441_ (.A(net119),
    .B(net413),
    .Y(_12453_));
 OA21x2_ASAP7_75t_R _32442_ (.A1(net413),
    .A2(_01750_),
    .B(_12453_),
    .Y(_12454_));
 AO21x1_ASAP7_75t_R _32443_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12454_),
    .Y(_12455_));
 OAI21x1_ASAP7_75t_R _32444_ (.A1(_01783_),
    .A2(_12348_),
    .B(_12455_),
    .Y(_04434_));
 NAND2x1_ASAP7_75t_R _32445_ (.A(net120),
    .B(_01815_),
    .Y(_12456_));
 OA21x2_ASAP7_75t_R _32446_ (.A1(_01815_),
    .A2(_01749_),
    .B(_12456_),
    .Y(_12457_));
 AO21x1_ASAP7_75t_R _32447_ (.A1(_06674_),
    .A2(_12347_),
    .B(_12457_),
    .Y(_12458_));
 OAI21x1_ASAP7_75t_R _32448_ (.A1(_01782_),
    .A2(_12348_),
    .B(_12458_),
    .Y(_04435_));
 AND2x2_ASAP7_75t_R _32449_ (.A(_06538_),
    .B(_01815_),
    .Y(_12459_));
 AO221x1_ASAP7_75t_R _32450_ (.A1(_06509_),
    .A2(_01748_),
    .B1(_06674_),
    .B2(_12347_),
    .C(_12459_),
    .Y(_12460_));
 OAI21x1_ASAP7_75t_R _32451_ (.A1(_01781_),
    .A2(_12348_),
    .B(_12460_),
    .Y(_04436_));
 OR3x4_ASAP7_75t_R _32452_ (.A(_00239_),
    .B(_06509_),
    .C(_06670_),
    .Y(_12461_));
 TAPCELL_ASAP7_75t_R PHY_92 ();
 TAPCELL_ASAP7_75t_R PHY_91 ();
 TAPCELL_ASAP7_75t_R PHY_90 ();
 NAND2x1_ASAP7_75t_R _32456_ (.A(_01780_),
    .B(_12461_),
    .Y(_12465_));
 OA21x2_ASAP7_75t_R _32457_ (.A1(net96),
    .A2(_12461_),
    .B(_12465_),
    .Y(_04437_));
 NAND2x1_ASAP7_75t_R _32458_ (.A(_01779_),
    .B(_12461_),
    .Y(_12466_));
 OA21x2_ASAP7_75t_R _32459_ (.A1(net107),
    .A2(_12461_),
    .B(_12466_),
    .Y(_04438_));
 NAND2x1_ASAP7_75t_R _32460_ (.A(_01778_),
    .B(_12461_),
    .Y(_12467_));
 OA21x2_ASAP7_75t_R _32461_ (.A1(net118),
    .A2(_12461_),
    .B(_12467_),
    .Y(_04439_));
 NAND2x1_ASAP7_75t_R _32462_ (.A(_01777_),
    .B(_12461_),
    .Y(_12468_));
 OA21x2_ASAP7_75t_R _32463_ (.A1(net121),
    .A2(_12461_),
    .B(_12468_),
    .Y(_04440_));
 NAND2x1_ASAP7_75t_R _32464_ (.A(_01776_),
    .B(_12461_),
    .Y(_12469_));
 OA21x2_ASAP7_75t_R _32465_ (.A1(net122),
    .A2(_12461_),
    .B(_12469_),
    .Y(_04441_));
 NAND2x1_ASAP7_75t_R _32466_ (.A(_01775_),
    .B(_12461_),
    .Y(_12470_));
 OA21x2_ASAP7_75t_R _32467_ (.A1(net123),
    .A2(_12461_),
    .B(_12470_),
    .Y(_04442_));
 NAND2x1_ASAP7_75t_R _32468_ (.A(_01774_),
    .B(_12461_),
    .Y(_12471_));
 OA21x2_ASAP7_75t_R _32469_ (.A1(net124),
    .A2(_12461_),
    .B(_12471_),
    .Y(_04443_));
 TAPCELL_ASAP7_75t_R PHY_89 ();
 NAND2x1_ASAP7_75t_R _32471_ (.A(_01773_),
    .B(_12461_),
    .Y(_12473_));
 OA21x2_ASAP7_75t_R _32472_ (.A1(net125),
    .A2(_12461_),
    .B(_12473_),
    .Y(_04444_));
 NAND2x1_ASAP7_75t_R _32473_ (.A(_01772_),
    .B(_12461_),
    .Y(_12474_));
 OA21x2_ASAP7_75t_R _32474_ (.A1(net126),
    .A2(_12461_),
    .B(_12474_),
    .Y(_04445_));
 NAND2x1_ASAP7_75t_R _32475_ (.A(_01771_),
    .B(_12461_),
    .Y(_12475_));
 OA21x2_ASAP7_75t_R _32476_ (.A1(net127),
    .A2(_12461_),
    .B(_12475_),
    .Y(_04446_));
 TAPCELL_ASAP7_75t_R PHY_88 ();
 NAND2x1_ASAP7_75t_R _32478_ (.A(_01770_),
    .B(_12461_),
    .Y(_12477_));
 OA21x2_ASAP7_75t_R _32479_ (.A1(net97),
    .A2(_12461_),
    .B(_12477_),
    .Y(_04447_));
 NAND2x1_ASAP7_75t_R _32480_ (.A(_01769_),
    .B(_12461_),
    .Y(_12478_));
 OA21x2_ASAP7_75t_R _32481_ (.A1(net98),
    .A2(_12461_),
    .B(_12478_),
    .Y(_04448_));
 NAND2x1_ASAP7_75t_R _32482_ (.A(_01768_),
    .B(_12461_),
    .Y(_12479_));
 OA21x2_ASAP7_75t_R _32483_ (.A1(net99),
    .A2(_12461_),
    .B(_12479_),
    .Y(_04449_));
 NAND2x1_ASAP7_75t_R _32484_ (.A(_01767_),
    .B(_12461_),
    .Y(_12480_));
 OA21x2_ASAP7_75t_R _32485_ (.A1(net100),
    .A2(_12461_),
    .B(_12480_),
    .Y(_04450_));
 NAND2x1_ASAP7_75t_R _32486_ (.A(_01766_),
    .B(_12461_),
    .Y(_12481_));
 OA21x2_ASAP7_75t_R _32487_ (.A1(net101),
    .A2(_12461_),
    .B(_12481_),
    .Y(_04451_));
 NAND2x1_ASAP7_75t_R _32488_ (.A(_01765_),
    .B(_12461_),
    .Y(_12482_));
 OA21x2_ASAP7_75t_R _32489_ (.A1(net102),
    .A2(_12461_),
    .B(_12482_),
    .Y(_04452_));
 NAND2x1_ASAP7_75t_R _32490_ (.A(_01764_),
    .B(_12461_),
    .Y(_12483_));
 OA21x2_ASAP7_75t_R _32491_ (.A1(net103),
    .A2(_12461_),
    .B(_12483_),
    .Y(_04453_));
 TAPCELL_ASAP7_75t_R PHY_87 ();
 NAND2x1_ASAP7_75t_R _32493_ (.A(_01763_),
    .B(_12461_),
    .Y(_12485_));
 OA21x2_ASAP7_75t_R _32494_ (.A1(net104),
    .A2(_12461_),
    .B(_12485_),
    .Y(_04454_));
 NAND2x1_ASAP7_75t_R _32495_ (.A(_01762_),
    .B(_12461_),
    .Y(_12486_));
 OA21x2_ASAP7_75t_R _32496_ (.A1(net105),
    .A2(_12461_),
    .B(_12486_),
    .Y(_04455_));
 NAND2x1_ASAP7_75t_R _32497_ (.A(_01761_),
    .B(_12461_),
    .Y(_12487_));
 OA21x2_ASAP7_75t_R _32498_ (.A1(net106),
    .A2(_12461_),
    .B(_12487_),
    .Y(_04456_));
 TAPCELL_ASAP7_75t_R PHY_86 ();
 NAND2x1_ASAP7_75t_R _32500_ (.A(_01760_),
    .B(_12461_),
    .Y(_12489_));
 OA21x2_ASAP7_75t_R _32501_ (.A1(net108),
    .A2(_12461_),
    .B(_12489_),
    .Y(_04457_));
 NAND2x1_ASAP7_75t_R _32502_ (.A(_01759_),
    .B(_12461_),
    .Y(_12490_));
 OA21x2_ASAP7_75t_R _32503_ (.A1(net109),
    .A2(_12461_),
    .B(_12490_),
    .Y(_04458_));
 NAND2x1_ASAP7_75t_R _32504_ (.A(_01758_),
    .B(_12461_),
    .Y(_12491_));
 OA21x2_ASAP7_75t_R _32505_ (.A1(net110),
    .A2(_12461_),
    .B(_12491_),
    .Y(_04459_));
 NAND2x1_ASAP7_75t_R _32506_ (.A(_01757_),
    .B(_12461_),
    .Y(_12492_));
 OA21x2_ASAP7_75t_R _32507_ (.A1(net111),
    .A2(_12461_),
    .B(_12492_),
    .Y(_04460_));
 NAND2x1_ASAP7_75t_R _32508_ (.A(_01756_),
    .B(_12461_),
    .Y(_12493_));
 OA21x2_ASAP7_75t_R _32509_ (.A1(net112),
    .A2(_12461_),
    .B(_12493_),
    .Y(_04461_));
 NAND2x1_ASAP7_75t_R _32510_ (.A(_01755_),
    .B(_12461_),
    .Y(_12494_));
 OA21x2_ASAP7_75t_R _32511_ (.A1(net113),
    .A2(_12461_),
    .B(_12494_),
    .Y(_04462_));
 NAND2x1_ASAP7_75t_R _32512_ (.A(_01754_),
    .B(_12461_),
    .Y(_12495_));
 OA21x2_ASAP7_75t_R _32513_ (.A1(net114),
    .A2(_12461_),
    .B(_12495_),
    .Y(_04463_));
 NAND2x1_ASAP7_75t_R _32514_ (.A(_01753_),
    .B(_12461_),
    .Y(_12496_));
 OA21x2_ASAP7_75t_R _32515_ (.A1(net115),
    .A2(_12461_),
    .B(_12496_),
    .Y(_04464_));
 NAND2x1_ASAP7_75t_R _32516_ (.A(_01752_),
    .B(_12461_),
    .Y(_12497_));
 OA21x2_ASAP7_75t_R _32517_ (.A1(net116),
    .A2(_12461_),
    .B(_12497_),
    .Y(_04465_));
 NAND2x1_ASAP7_75t_R _32518_ (.A(_01751_),
    .B(_12461_),
    .Y(_12498_));
 OA21x2_ASAP7_75t_R _32519_ (.A1(net117),
    .A2(_12461_),
    .B(_12498_),
    .Y(_04466_));
 NAND2x1_ASAP7_75t_R _32520_ (.A(_01750_),
    .B(_12461_),
    .Y(_12499_));
 OA21x2_ASAP7_75t_R _32521_ (.A1(net119),
    .A2(_12461_),
    .B(_12499_),
    .Y(_04467_));
 NAND2x1_ASAP7_75t_R _32522_ (.A(_01749_),
    .B(_12461_),
    .Y(_12500_));
 OA21x2_ASAP7_75t_R _32523_ (.A1(net120),
    .A2(_12461_),
    .B(_12500_),
    .Y(_04468_));
 NAND2x1_ASAP7_75t_R _32524_ (.A(_01748_),
    .B(_12461_),
    .Y(_12501_));
 OA21x2_ASAP7_75t_R _32525_ (.A1(net94),
    .A2(_12461_),
    .B(_12501_),
    .Y(_04469_));
 INVx1_ASAP7_75t_R _32526_ (.A(net61),
    .Y(_12502_));
 NAND2x1_ASAP7_75t_R _32527_ (.A(_01747_),
    .B(_12502_),
    .Y(_04470_));
 NAND2x1_ASAP7_75t_R _32528_ (.A(_05677_),
    .B(_06258_),
    .Y(_12503_));
 NAND2x1_ASAP7_75t_R _32529_ (.A(_06186_),
    .B(_12503_),
    .Y(_04503_));
 TAPCELL_ASAP7_75t_R PHY_85 ();
 TAPCELL_ASAP7_75t_R PHY_84 ();
 AND2x2_ASAP7_75t_R _32532_ (.A(net417),
    .B(net96),
    .Y(_12506_));
 AO21x1_ASAP7_75t_R _32533_ (.A1(_06528_),
    .A2(net103),
    .B(_12506_),
    .Y(_12507_));
 NAND2x1_ASAP7_75t_R _32534_ (.A(net417),
    .B(_01846_),
    .Y(_12508_));
 OA211x2_ASAP7_75t_R _32535_ (.A1(net417),
    .A2(_12311_),
    .B(_12508_),
    .C(_06537_),
    .Y(_12509_));
 AO21x2_ASAP7_75t_R _32536_ (.A1(_00240_),
    .A2(_12507_),
    .B(_12509_),
    .Y(_12510_));
 TAPCELL_ASAP7_75t_R PHY_83 ();
 TAPCELL_ASAP7_75t_R PHY_82 ();
 TAPCELL_ASAP7_75t_R PHY_81 ();
 NAND2x1_ASAP7_75t_R _32540_ (.A(_01723_),
    .B(_09270_),
    .Y(_12514_));
 OA21x2_ASAP7_75t_R _32541_ (.A1(_09270_),
    .A2(_12510_),
    .B(_12514_),
    .Y(_02597_));
 AND2x2_ASAP7_75t_R _32542_ (.A(net417),
    .B(net107),
    .Y(_12515_));
 AO21x1_ASAP7_75t_R _32543_ (.A1(_06528_),
    .A2(net104),
    .B(_12515_),
    .Y(_12516_));
 NAND2x1_ASAP7_75t_R _32544_ (.A(net416),
    .B(_01845_),
    .Y(_12517_));
 OA211x2_ASAP7_75t_R _32545_ (.A1(net416),
    .A2(_12313_),
    .B(_12517_),
    .C(_06537_),
    .Y(_12518_));
 AO21x2_ASAP7_75t_R _32546_ (.A1(_00240_),
    .A2(_12516_),
    .B(_12518_),
    .Y(_12519_));
 TAPCELL_ASAP7_75t_R PHY_80 ();
 TAPCELL_ASAP7_75t_R PHY_79 ();
 NAND2x1_ASAP7_75t_R _32549_ (.A(_00164_),
    .B(_09270_),
    .Y(_12522_));
 OA21x2_ASAP7_75t_R _32550_ (.A1(_09270_),
    .A2(_12519_),
    .B(_12522_),
    .Y(_02598_));
 AND2x2_ASAP7_75t_R _32551_ (.A(net416),
    .B(net118),
    .Y(_12523_));
 AO21x1_ASAP7_75t_R _32552_ (.A1(_06528_),
    .A2(net105),
    .B(_12523_),
    .Y(_12524_));
 NAND2x1_ASAP7_75t_R _32553_ (.A(net416),
    .B(_01844_),
    .Y(_12525_));
 OA211x2_ASAP7_75t_R _32554_ (.A1(net416),
    .A2(_12315_),
    .B(_12525_),
    .C(_06537_),
    .Y(_12526_));
 AO21x2_ASAP7_75t_R _32555_ (.A1(net414),
    .A2(_12524_),
    .B(_12526_),
    .Y(_12527_));
 TAPCELL_ASAP7_75t_R PHY_78 ();
 NAND2x1_ASAP7_75t_R _32557_ (.A(_00166_),
    .B(_09270_),
    .Y(_12529_));
 OA21x2_ASAP7_75t_R _32558_ (.A1(_09270_),
    .A2(_12527_),
    .B(_12529_),
    .Y(_02599_));
 AND2x2_ASAP7_75t_R _32559_ (.A(net417),
    .B(net121),
    .Y(_12530_));
 AO21x1_ASAP7_75t_R _32560_ (.A1(_06528_),
    .A2(net106),
    .B(_12530_),
    .Y(_12531_));
 NAND2x1_ASAP7_75t_R _32561_ (.A(net417),
    .B(_01843_),
    .Y(_12532_));
 OA211x2_ASAP7_75t_R _32562_ (.A1(net417),
    .A2(_12317_),
    .B(_12532_),
    .C(_06537_),
    .Y(_12533_));
 AO21x2_ASAP7_75t_R _32563_ (.A1(_00240_),
    .A2(_12531_),
    .B(_12533_),
    .Y(_12534_));
 TAPCELL_ASAP7_75t_R PHY_77 ();
 NAND2x1_ASAP7_75t_R _32565_ (.A(_00169_),
    .B(_09270_),
    .Y(_12536_));
 OA21x2_ASAP7_75t_R _32566_ (.A1(_09270_),
    .A2(_12534_),
    .B(_12536_),
    .Y(_02600_));
 AND2x2_ASAP7_75t_R _32567_ (.A(net417),
    .B(net122),
    .Y(_12537_));
 AO21x1_ASAP7_75t_R _32568_ (.A1(_06528_),
    .A2(net108),
    .B(_12537_),
    .Y(_12538_));
 NAND2x1_ASAP7_75t_R _32569_ (.A(net417),
    .B(_01842_),
    .Y(_12539_));
 OA211x2_ASAP7_75t_R _32570_ (.A1(net417),
    .A2(_12319_),
    .B(_12539_),
    .C(_06537_),
    .Y(_12540_));
 AO21x2_ASAP7_75t_R _32571_ (.A1(_00240_),
    .A2(_12538_),
    .B(_12540_),
    .Y(_12541_));
 TAPCELL_ASAP7_75t_R PHY_76 ();
 NAND2x1_ASAP7_75t_R _32573_ (.A(_00173_),
    .B(_09270_),
    .Y(_12543_));
 OA21x2_ASAP7_75t_R _32574_ (.A1(_09270_),
    .A2(_12541_),
    .B(_12543_),
    .Y(_02601_));
 AND2x2_ASAP7_75t_R _32575_ (.A(net416),
    .B(net123),
    .Y(_12544_));
 AO21x1_ASAP7_75t_R _32576_ (.A1(_06528_),
    .A2(net109),
    .B(_12544_),
    .Y(_12545_));
 NAND2x1_ASAP7_75t_R _32577_ (.A(net416),
    .B(_01841_),
    .Y(_12546_));
 OA211x2_ASAP7_75t_R _32578_ (.A1(net416),
    .A2(_12321_),
    .B(_12546_),
    .C(_06537_),
    .Y(_12547_));
 AO21x2_ASAP7_75t_R _32579_ (.A1(_00240_),
    .A2(_12545_),
    .B(_12547_),
    .Y(_12548_));
 TAPCELL_ASAP7_75t_R PHY_75 ();
 NAND2x1_ASAP7_75t_R _32581_ (.A(_00176_),
    .B(_09270_),
    .Y(_12550_));
 OA21x2_ASAP7_75t_R _32582_ (.A1(_09270_),
    .A2(_12548_),
    .B(_12550_),
    .Y(_02602_));
 AND2x2_ASAP7_75t_R _32583_ (.A(_00662_),
    .B(net124),
    .Y(_12551_));
 AO21x1_ASAP7_75t_R _32584_ (.A1(_06528_),
    .A2(net110),
    .B(_12551_),
    .Y(_12552_));
 NAND2x1_ASAP7_75t_R _32585_ (.A(_00662_),
    .B(_01840_),
    .Y(_12553_));
 OA211x2_ASAP7_75t_R _32586_ (.A1(_00662_),
    .A2(_12323_),
    .B(_12553_),
    .C(_06537_),
    .Y(_12554_));
 AO21x2_ASAP7_75t_R _32587_ (.A1(_00240_),
    .A2(_12552_),
    .B(_12554_),
    .Y(_12555_));
 TAPCELL_ASAP7_75t_R PHY_74 ();
 NAND2x1_ASAP7_75t_R _32589_ (.A(_00179_),
    .B(_09270_),
    .Y(_12557_));
 OA21x2_ASAP7_75t_R _32590_ (.A1(_09270_),
    .A2(_12555_),
    .B(_12557_),
    .Y(_02603_));
 AND2x2_ASAP7_75t_R _32591_ (.A(net417),
    .B(net125),
    .Y(_12558_));
 AO21x1_ASAP7_75t_R _32592_ (.A1(_06528_),
    .A2(net111),
    .B(_12558_),
    .Y(_12559_));
 NAND2x1_ASAP7_75t_R _32593_ (.A(net417),
    .B(_01839_),
    .Y(_12560_));
 OA211x2_ASAP7_75t_R _32594_ (.A1(net417),
    .A2(_12325_),
    .B(_12560_),
    .C(_06537_),
    .Y(_12561_));
 AO21x2_ASAP7_75t_R _32595_ (.A1(_00240_),
    .A2(_12559_),
    .B(_12561_),
    .Y(_12562_));
 TAPCELL_ASAP7_75t_R PHY_73 ();
 NAND2x1_ASAP7_75t_R _32597_ (.A(_00181_),
    .B(_09270_),
    .Y(_12564_));
 OA21x2_ASAP7_75t_R _32598_ (.A1(_09270_),
    .A2(_12562_),
    .B(_12564_),
    .Y(_02604_));
 TAPCELL_ASAP7_75t_R PHY_72 ();
 TAPCELL_ASAP7_75t_R PHY_71 ();
 AND2x2_ASAP7_75t_R _32601_ (.A(net416),
    .B(net126),
    .Y(_12567_));
 AO21x1_ASAP7_75t_R _32602_ (.A1(_06528_),
    .A2(net112),
    .B(_12567_),
    .Y(_12568_));
 NAND2x1_ASAP7_75t_R _32603_ (.A(net416),
    .B(_01838_),
    .Y(_12569_));
 OA211x2_ASAP7_75t_R _32604_ (.A1(net416),
    .A2(_12327_),
    .B(_12569_),
    .C(_06537_),
    .Y(_12570_));
 AO21x2_ASAP7_75t_R _32605_ (.A1(_00240_),
    .A2(_12568_),
    .B(_12570_),
    .Y(_12571_));
 TAPCELL_ASAP7_75t_R PHY_70 ();
 TAPCELL_ASAP7_75t_R PHY_69 ();
 NAND2x1_ASAP7_75t_R _32608_ (.A(_00185_),
    .B(_09270_),
    .Y(_12574_));
 OA21x2_ASAP7_75t_R _32609_ (.A1(_09270_),
    .A2(_12571_),
    .B(_12574_),
    .Y(_02605_));
 AND2x2_ASAP7_75t_R _32610_ (.A(net417),
    .B(net127),
    .Y(_12575_));
 AO21x1_ASAP7_75t_R _32611_ (.A1(_06528_),
    .A2(net113),
    .B(_12575_),
    .Y(_12576_));
 NAND2x1_ASAP7_75t_R _32612_ (.A(net417),
    .B(_01837_),
    .Y(_12577_));
 OA211x2_ASAP7_75t_R _32613_ (.A1(net417),
    .A2(_12329_),
    .B(_12577_),
    .C(_06537_),
    .Y(_12578_));
 AO21x2_ASAP7_75t_R _32614_ (.A1(_00240_),
    .A2(_12576_),
    .B(_12578_),
    .Y(_12579_));
 NAND2x1_ASAP7_75t_R _32615_ (.A(_00188_),
    .B(_09270_),
    .Y(_12580_));
 OA21x2_ASAP7_75t_R _32616_ (.A1(_09270_),
    .A2(_12579_),
    .B(_12580_),
    .Y(_02606_));
 AND2x2_ASAP7_75t_R _32617_ (.A(net417),
    .B(net97),
    .Y(_12581_));
 AO21x1_ASAP7_75t_R _32618_ (.A1(_06528_),
    .A2(net114),
    .B(_12581_),
    .Y(_12582_));
 NAND2x1_ASAP7_75t_R _32619_ (.A(net417),
    .B(_01836_),
    .Y(_12583_));
 OA211x2_ASAP7_75t_R _32620_ (.A1(net417),
    .A2(_12331_),
    .B(_12583_),
    .C(_06537_),
    .Y(_12584_));
 AO21x2_ASAP7_75t_R _32621_ (.A1(_00240_),
    .A2(_12582_),
    .B(_12584_),
    .Y(_12585_));
 TAPCELL_ASAP7_75t_R PHY_68 ();
 NAND2x1_ASAP7_75t_R _32623_ (.A(_00192_),
    .B(_09270_),
    .Y(_12587_));
 OA21x2_ASAP7_75t_R _32624_ (.A1(_09270_),
    .A2(_12585_),
    .B(_12587_),
    .Y(_02607_));
 AND2x2_ASAP7_75t_R _32625_ (.A(net417),
    .B(net98),
    .Y(_12588_));
 AO21x1_ASAP7_75t_R _32626_ (.A1(_06528_),
    .A2(net115),
    .B(_12588_),
    .Y(_12589_));
 NAND2x1_ASAP7_75t_R _32627_ (.A(net417),
    .B(_01835_),
    .Y(_12590_));
 OA211x2_ASAP7_75t_R _32628_ (.A1(net417),
    .A2(_12333_),
    .B(_12590_),
    .C(_06537_),
    .Y(_12591_));
 AO21x2_ASAP7_75t_R _32629_ (.A1(_00240_),
    .A2(_12589_),
    .B(_12591_),
    .Y(_12592_));
 TAPCELL_ASAP7_75t_R PHY_67 ();
 TAPCELL_ASAP7_75t_R PHY_66 ();
 NAND2x1_ASAP7_75t_R _32632_ (.A(_00195_),
    .B(_09270_),
    .Y(_12595_));
 OA21x2_ASAP7_75t_R _32633_ (.A1(_09270_),
    .A2(_12592_),
    .B(_12595_),
    .Y(_02608_));
 AND2x2_ASAP7_75t_R _32634_ (.A(net416),
    .B(net99),
    .Y(_12596_));
 AO21x1_ASAP7_75t_R _32635_ (.A1(_06528_),
    .A2(net116),
    .B(_12596_),
    .Y(_12597_));
 NAND2x1_ASAP7_75t_R _32636_ (.A(net416),
    .B(_01834_),
    .Y(_12598_));
 OA211x2_ASAP7_75t_R _32637_ (.A1(net416),
    .A2(_12335_),
    .B(_12598_),
    .C(_06537_),
    .Y(_12599_));
 AO21x2_ASAP7_75t_R _32638_ (.A1(net414),
    .A2(_12597_),
    .B(_12599_),
    .Y(_12600_));
 TAPCELL_ASAP7_75t_R PHY_65 ();
 TAPCELL_ASAP7_75t_R PHY_64 ();
 TAPCELL_ASAP7_75t_R PHY_63 ();
 NAND2x1_ASAP7_75t_R _32642_ (.A(_00198_),
    .B(_09270_),
    .Y(_12604_));
 OA21x2_ASAP7_75t_R _32643_ (.A1(_09270_),
    .A2(_12600_),
    .B(_12604_),
    .Y(_02609_));
 AND2x2_ASAP7_75t_R _32644_ (.A(net416),
    .B(net100),
    .Y(_12605_));
 AO21x1_ASAP7_75t_R _32645_ (.A1(_06528_),
    .A2(net117),
    .B(_12605_),
    .Y(_12606_));
 NAND2x1_ASAP7_75t_R _32646_ (.A(net416),
    .B(_01833_),
    .Y(_12607_));
 OA211x2_ASAP7_75t_R _32647_ (.A1(net416),
    .A2(_12337_),
    .B(_12607_),
    .C(_06537_),
    .Y(_12608_));
 AO21x2_ASAP7_75t_R _32648_ (.A1(net414),
    .A2(_12606_),
    .B(_12608_),
    .Y(_12609_));
 TAPCELL_ASAP7_75t_R PHY_62 ();
 TAPCELL_ASAP7_75t_R PHY_61 ();
 TAPCELL_ASAP7_75t_R PHY_60 ();
 NAND2x1_ASAP7_75t_R _32652_ (.A(_00200_),
    .B(_09270_),
    .Y(_12613_));
 OA21x2_ASAP7_75t_R _32653_ (.A1(_09270_),
    .A2(_12609_),
    .B(_12613_),
    .Y(_02610_));
 AND2x2_ASAP7_75t_R _32654_ (.A(net417),
    .B(net101),
    .Y(_12614_));
 AO21x1_ASAP7_75t_R _32655_ (.A1(_06528_),
    .A2(net119),
    .B(_12614_),
    .Y(_12615_));
 NAND2x1_ASAP7_75t_R _32656_ (.A(net417),
    .B(_01832_),
    .Y(_12616_));
 OA211x2_ASAP7_75t_R _32657_ (.A1(net417),
    .A2(_12339_),
    .B(_12616_),
    .C(_06537_),
    .Y(_12617_));
 AO21x2_ASAP7_75t_R _32658_ (.A1(_00240_),
    .A2(_12615_),
    .B(_12617_),
    .Y(_12618_));
 TAPCELL_ASAP7_75t_R PHY_59 ();
 TAPCELL_ASAP7_75t_R PHY_58 ();
 NAND2x1_ASAP7_75t_R _32661_ (.A(_00203_),
    .B(_09270_),
    .Y(_12621_));
 OA21x2_ASAP7_75t_R _32662_ (.A1(_09270_),
    .A2(_12618_),
    .B(_12621_),
    .Y(_02611_));
 AND2x2_ASAP7_75t_R _32663_ (.A(net102),
    .B(net416),
    .Y(_12622_));
 AO21x1_ASAP7_75t_R _32664_ (.A1(net120),
    .A2(_06528_),
    .B(_12622_),
    .Y(_12623_));
 NAND2x1_ASAP7_75t_R _32665_ (.A(net416),
    .B(_01831_),
    .Y(_12624_));
 OA211x2_ASAP7_75t_R _32666_ (.A1(net416),
    .A2(_12340_),
    .B(_12624_),
    .C(_06537_),
    .Y(_12625_));
 AO21x2_ASAP7_75t_R _32667_ (.A1(net414),
    .A2(_12623_),
    .B(_12625_),
    .Y(_12626_));
 TAPCELL_ASAP7_75t_R PHY_57 ();
 TAPCELL_ASAP7_75t_R PHY_56 ();
 NAND2x1_ASAP7_75t_R _32670_ (.A(_00205_),
    .B(_09270_),
    .Y(_12629_));
 OA21x2_ASAP7_75t_R _32671_ (.A1(_09270_),
    .A2(_12626_),
    .B(_12629_),
    .Y(_02612_));
 TAPCELL_ASAP7_75t_R PHY_55 ();
 AND2x4_ASAP7_75t_R _32673_ (.A(_12510_),
    .B(_12519_),
    .Y(_12631_));
 NAND2x1_ASAP7_75t_R _32674_ (.A(_09257_),
    .B(_12631_),
    .Y(_12632_));
 OA21x2_ASAP7_75t_R _32675_ (.A1(_05549_),
    .A2(_09257_),
    .B(_12632_),
    .Y(_02613_));
 INVx1_ASAP7_75t_R _32676_ (.A(_01814_),
    .Y(_12633_));
 OA22x2_ASAP7_75t_R _32677_ (.A1(_00239_),
    .A2(_01781_),
    .B1(_12345_),
    .B2(_06538_),
    .Y(_12634_));
 OR4x1_ASAP7_75t_R _32678_ (.A(_00662_),
    .B(_12633_),
    .C(_09270_),
    .D(_12634_),
    .Y(_12635_));
 OAI21x1_ASAP7_75t_R _32679_ (.A1(_01722_),
    .A2(_09257_),
    .B(_12635_),
    .Y(_02614_));
 OA21x2_ASAP7_75t_R _32680_ (.A1(_06538_),
    .A2(_06536_),
    .B(_00239_),
    .Y(_12636_));
 OAI21x1_ASAP7_75t_R _32681_ (.A1(_00662_),
    .A2(_12636_),
    .B(_06540_),
    .Y(_12637_));
 NOR2x1_ASAP7_75t_R _32682_ (.A(_01781_),
    .B(_09256_),
    .Y(_12638_));
 OR4x1_ASAP7_75t_R _32683_ (.A(_00662_),
    .B(_00239_),
    .C(_12633_),
    .D(_12638_),
    .Y(_12639_));
 AND3x1_ASAP7_75t_R _32684_ (.A(_09257_),
    .B(_12637_),
    .C(_12639_),
    .Y(_12640_));
 AO21x1_ASAP7_75t_R _32685_ (.A1(_05719_),
    .A2(_09270_),
    .B(_12640_),
    .Y(_02615_));
 NAND2x1_ASAP7_75t_R _32686_ (.A(_00662_),
    .B(_09257_),
    .Y(_12641_));
 OA21x2_ASAP7_75t_R _32687_ (.A1(\cs_registers_i.pc_id_i[1] ),
    .A2(_09257_),
    .B(_12641_),
    .Y(_02616_));
 NAND2x1_ASAP7_75t_R _32688_ (.A(_17536_),
    .B(_09257_),
    .Y(_12642_));
 OA21x2_ASAP7_75t_R _32689_ (.A1(\cs_registers_i.pc_id_i[2] ),
    .A2(_09257_),
    .B(_12642_),
    .Y(_02617_));
 NAND2x1_ASAP7_75t_R _32690_ (.A(_01606_),
    .B(_09257_),
    .Y(_12643_));
 OA21x2_ASAP7_75t_R _32691_ (.A1(\cs_registers_i.pc_id_i[3] ),
    .A2(_09257_),
    .B(_12643_),
    .Y(_02618_));
 NAND2x1_ASAP7_75t_R _32692_ (.A(_01605_),
    .B(_09257_),
    .Y(_12644_));
 OA21x2_ASAP7_75t_R _32693_ (.A1(_14764_),
    .A2(_09257_),
    .B(_12644_),
    .Y(_02619_));
 NAND2x1_ASAP7_75t_R _32694_ (.A(_01604_),
    .B(_09257_),
    .Y(_12645_));
 OA21x2_ASAP7_75t_R _32695_ (.A1(\cs_registers_i.pc_id_i[5] ),
    .A2(_09257_),
    .B(_12645_),
    .Y(_02620_));
 NAND2x1_ASAP7_75t_R _32696_ (.A(_01603_),
    .B(_09257_),
    .Y(_12646_));
 OA21x2_ASAP7_75t_R _32697_ (.A1(_14937_),
    .A2(_09257_),
    .B(_12646_),
    .Y(_02621_));
 NAND2x1_ASAP7_75t_R _32698_ (.A(_01602_),
    .B(_09257_),
    .Y(_12647_));
 OA21x2_ASAP7_75t_R _32699_ (.A1(\cs_registers_i.pc_id_i[7] ),
    .A2(_09257_),
    .B(_12647_),
    .Y(_02622_));
 TAPCELL_ASAP7_75t_R PHY_54 ();
 AND2x2_ASAP7_75t_R _32701_ (.A(_01601_),
    .B(_09257_),
    .Y(_12649_));
 AOI21x1_ASAP7_75t_R _32702_ (.A1(_00186_),
    .A2(_09270_),
    .B(_12649_),
    .Y(_02623_));
 TAPCELL_ASAP7_75t_R PHY_53 ();
 NAND2x1_ASAP7_75t_R _32704_ (.A(_01600_),
    .B(_09257_),
    .Y(_12651_));
 OA21x2_ASAP7_75t_R _32705_ (.A1(\cs_registers_i.pc_id_i[9] ),
    .A2(_09257_),
    .B(_12651_),
    .Y(_02624_));
 TAPCELL_ASAP7_75t_R PHY_52 ();
 NAND2x1_ASAP7_75t_R _32707_ (.A(_01599_),
    .B(_09257_),
    .Y(_12653_));
 OA21x2_ASAP7_75t_R _32708_ (.A1(_15158_),
    .A2(_09257_),
    .B(_12653_),
    .Y(_02625_));
 NAND2x1_ASAP7_75t_R _32709_ (.A(_01598_),
    .B(_09257_),
    .Y(_12654_));
 OA21x2_ASAP7_75t_R _32710_ (.A1(\cs_registers_i.pc_id_i[11] ),
    .A2(_09257_),
    .B(_12654_),
    .Y(_02626_));
 AND2x2_ASAP7_75t_R _32711_ (.A(_01597_),
    .B(_09257_),
    .Y(_12655_));
 AOI21x1_ASAP7_75t_R _32712_ (.A1(_00199_),
    .A2(_09270_),
    .B(_12655_),
    .Y(_02627_));
 NAND2x1_ASAP7_75t_R _32713_ (.A(_01596_),
    .B(_09257_),
    .Y(_12656_));
 OA21x2_ASAP7_75t_R _32714_ (.A1(\cs_registers_i.pc_id_i[13] ),
    .A2(_09257_),
    .B(_12656_),
    .Y(_02628_));
 AND2x2_ASAP7_75t_R _32715_ (.A(_01595_),
    .B(_09257_),
    .Y(_12657_));
 AOI21x1_ASAP7_75t_R _32716_ (.A1(_00204_),
    .A2(_09270_),
    .B(_12657_),
    .Y(_02629_));
 NAND2x1_ASAP7_75t_R _32717_ (.A(_01594_),
    .B(_09257_),
    .Y(_12658_));
 OA21x2_ASAP7_75t_R _32718_ (.A1(\cs_registers_i.pc_id_i[15] ),
    .A2(_09257_),
    .B(_12658_),
    .Y(_02630_));
 AND2x2_ASAP7_75t_R _32719_ (.A(_01593_),
    .B(_09257_),
    .Y(_12659_));
 AOI21x1_ASAP7_75t_R _32720_ (.A1(_00208_),
    .A2(_09270_),
    .B(_12659_),
    .Y(_02631_));
 NAND2x1_ASAP7_75t_R _32721_ (.A(_01592_),
    .B(_09257_),
    .Y(_12660_));
 OA21x2_ASAP7_75t_R _32722_ (.A1(\cs_registers_i.pc_id_i[17] ),
    .A2(_09257_),
    .B(_12660_),
    .Y(_02632_));
 AND2x2_ASAP7_75t_R _32723_ (.A(_01591_),
    .B(_09257_),
    .Y(_12661_));
 AOI21x1_ASAP7_75t_R _32724_ (.A1(_00211_),
    .A2(_09270_),
    .B(_12661_),
    .Y(_02633_));
 NAND2x1_ASAP7_75t_R _32725_ (.A(_01590_),
    .B(_09257_),
    .Y(_12662_));
 OA21x2_ASAP7_75t_R _32726_ (.A1(\cs_registers_i.pc_id_i[19] ),
    .A2(_09257_),
    .B(_12662_),
    .Y(_02634_));
 AND2x2_ASAP7_75t_R _32727_ (.A(_01589_),
    .B(_09257_),
    .Y(_12663_));
 AOI21x1_ASAP7_75t_R _32728_ (.A1(_00214_),
    .A2(_09270_),
    .B(_12663_),
    .Y(_02635_));
 NAND2x1_ASAP7_75t_R _32729_ (.A(_01588_),
    .B(_09257_),
    .Y(_12664_));
 OA21x2_ASAP7_75t_R _32730_ (.A1(\cs_registers_i.pc_id_i[21] ),
    .A2(_09257_),
    .B(_12664_),
    .Y(_02636_));
 AND2x2_ASAP7_75t_R _32731_ (.A(_01587_),
    .B(_09257_),
    .Y(_12665_));
 AOI21x1_ASAP7_75t_R _32732_ (.A1(_00217_),
    .A2(_09270_),
    .B(_12665_),
    .Y(_02637_));
 NAND2x1_ASAP7_75t_R _32733_ (.A(_01586_),
    .B(_09257_),
    .Y(_12666_));
 OA21x2_ASAP7_75t_R _32734_ (.A1(\cs_registers_i.pc_id_i[23] ),
    .A2(_09257_),
    .B(_12666_),
    .Y(_02638_));
 AND2x2_ASAP7_75t_R _32735_ (.A(_01585_),
    .B(_09257_),
    .Y(_12667_));
 AOI21x1_ASAP7_75t_R _32736_ (.A1(_00220_),
    .A2(_09270_),
    .B(_12667_),
    .Y(_02639_));
 NAND2x1_ASAP7_75t_R _32737_ (.A(_01584_),
    .B(_09257_),
    .Y(_12668_));
 OA21x2_ASAP7_75t_R _32738_ (.A1(\cs_registers_i.pc_id_i[25] ),
    .A2(_09257_),
    .B(_12668_),
    .Y(_02640_));
 AND2x2_ASAP7_75t_R _32739_ (.A(_01583_),
    .B(_09257_),
    .Y(_12669_));
 AOI21x1_ASAP7_75t_R _32740_ (.A1(_00223_),
    .A2(_09270_),
    .B(_12669_),
    .Y(_02641_));
 TAPCELL_ASAP7_75t_R PHY_51 ();
 NAND2x1_ASAP7_75t_R _32742_ (.A(_01582_),
    .B(_09257_),
    .Y(_12671_));
 OA21x2_ASAP7_75t_R _32743_ (.A1(\cs_registers_i.pc_id_i[27] ),
    .A2(_09257_),
    .B(_12671_),
    .Y(_02642_));
 AND2x2_ASAP7_75t_R _32744_ (.A(_01581_),
    .B(_09257_),
    .Y(_12672_));
 AOI21x1_ASAP7_75t_R _32745_ (.A1(_00226_),
    .A2(_09270_),
    .B(_12672_),
    .Y(_02643_));
 NAND2x1_ASAP7_75t_R _32746_ (.A(_01580_),
    .B(_09257_),
    .Y(_12673_));
 OA21x2_ASAP7_75t_R _32747_ (.A1(\cs_registers_i.pc_id_i[29] ),
    .A2(_09257_),
    .B(_12673_),
    .Y(_02644_));
 NAND2x1_ASAP7_75t_R _32748_ (.A(_01579_),
    .B(_09257_),
    .Y(_12674_));
 OA21x2_ASAP7_75t_R _32749_ (.A1(_05370_),
    .A2(_09257_),
    .B(_12674_),
    .Y(_02645_));
 AND2x2_ASAP7_75t_R _32750_ (.A(_01578_),
    .B(_09257_),
    .Y(_12675_));
 AOI21x1_ASAP7_75t_R _32751_ (.A1(_00230_),
    .A2(_09270_),
    .B(_12675_),
    .Y(_02646_));
 AND4x2_ASAP7_75t_R _32752_ (.A(_05582_),
    .B(_11107_),
    .C(_10973_),
    .D(_11497_),
    .Y(_12676_));
 AO21x1_ASAP7_75t_R _32753_ (.A1(_01577_),
    .A2(_11699_),
    .B(_06880_),
    .Y(_12677_));
 OAI22x1_ASAP7_75t_R _32754_ (.A1(_02140_),
    .A2(_06873_),
    .B1(_12676_),
    .B2(_12677_),
    .Y(_02863_));
 AO21x1_ASAP7_75t_R _32755_ (.A1(_01576_),
    .A2(_11699_),
    .B(_06880_),
    .Y(_12678_));
 OAI22x1_ASAP7_75t_R _32756_ (.A1(_17592_),
    .A2(_06873_),
    .B1(_12676_),
    .B2(_12678_),
    .Y(_02864_));
 NAND2x1_ASAP7_75t_R _32757_ (.A(_01875_),
    .B(_14628_),
    .Y(_12679_));
 OA21x2_ASAP7_75t_R _32758_ (.A1(_14577_),
    .A2(_14628_),
    .B(_12679_),
    .Y(_04341_));
 AND3x1_ASAP7_75t_R _32759_ (.A(_00279_),
    .B(_01875_),
    .C(_14626_),
    .Y(_12680_));
 AOI21x1_ASAP7_75t_R _32760_ (.A1(_01874_),
    .A2(_14628_),
    .B(_12680_),
    .Y(_04342_));
 INVx1_ASAP7_75t_R _32761_ (.A(_01847_),
    .Y(_12681_));
 AOI21x1_ASAP7_75t_R _32762_ (.A1(_00240_),
    .A2(_12516_),
    .B(_12518_),
    .Y(_12682_));
 AND2x6_ASAP7_75t_R _32763_ (.A(_12510_),
    .B(_12682_),
    .Y(_12683_));
 TAPCELL_ASAP7_75t_R PHY_50 ();
 AOI21x1_ASAP7_75t_R _32765_ (.A1(net414),
    .A2(_12623_),
    .B(_12625_),
    .Y(_12685_));
 OR3x4_ASAP7_75t_R _32766_ (.A(_12609_),
    .B(_12618_),
    .C(_12685_),
    .Y(_12686_));
 AOI21x1_ASAP7_75t_R _32767_ (.A1(_00240_),
    .A2(_12582_),
    .B(_12584_),
    .Y(_12687_));
 AOI21x1_ASAP7_75t_R _32768_ (.A1(net414),
    .A2(_12597_),
    .B(_12599_),
    .Y(_12688_));
 AO21x1_ASAP7_75t_R _32769_ (.A1(_12687_),
    .A2(_12592_),
    .B(_12688_),
    .Y(_12689_));
 OR2x2_ASAP7_75t_R _32770_ (.A(_12548_),
    .B(_12555_),
    .Y(_12690_));
 OR3x4_ASAP7_75t_R _32771_ (.A(_12527_),
    .B(_12534_),
    .C(_12690_),
    .Y(_12691_));
 OR2x2_ASAP7_75t_R _32772_ (.A(_12541_),
    .B(_12691_),
    .Y(_12692_));
 AND3x4_ASAP7_75t_R _32773_ (.A(_12609_),
    .B(_12618_),
    .C(_12685_),
    .Y(_12693_));
 NAND2x1_ASAP7_75t_R _32774_ (.A(_12688_),
    .B(_12693_),
    .Y(_12694_));
 OAI22x1_ASAP7_75t_R _32775_ (.A1(_12686_),
    .A2(_12689_),
    .B1(_12692_),
    .B2(_12694_),
    .Y(_12695_));
 AOI21x1_ASAP7_75t_R _32776_ (.A1(_00240_),
    .A2(_12507_),
    .B(_12509_),
    .Y(_12696_));
 AND2x6_ASAP7_75t_R _32777_ (.A(_12696_),
    .B(_12682_),
    .Y(_12697_));
 TAPCELL_ASAP7_75t_R PHY_49 ();
 AOI21x1_ASAP7_75t_R _32779_ (.A1(_00240_),
    .A2(_12615_),
    .B(_12617_),
    .Y(_12699_));
 AND2x2_ASAP7_75t_R _32780_ (.A(net297),
    .B(_12626_),
    .Y(_12700_));
 NOR2x2_ASAP7_75t_R _32781_ (.A(_12609_),
    .B(_12700_),
    .Y(_12701_));
 OR4x1_ASAP7_75t_R _32782_ (.A(_12562_),
    .B(_12579_),
    .C(_12585_),
    .D(_12592_),
    .Y(_12702_));
 OR2x4_ASAP7_75t_R _32783_ (.A(_12571_),
    .B(_12702_),
    .Y(_12703_));
 OR4x1_ASAP7_75t_R _32784_ (.A(_12600_),
    .B(_12618_),
    .C(_12690_),
    .D(_12703_),
    .Y(_12704_));
 NAND2x1_ASAP7_75t_R _32785_ (.A(_12701_),
    .B(_12704_),
    .Y(_12705_));
 AO22x1_ASAP7_75t_R _32786_ (.A1(_12683_),
    .A2(_12695_),
    .B1(_12697_),
    .B2(_12705_),
    .Y(_12706_));
 OR3x4_ASAP7_75t_R _32787_ (.A(_12609_),
    .B(_12618_),
    .C(_12626_),
    .Y(_12707_));
 TAPCELL_ASAP7_75t_R PHY_48 ();
 AND2x6_ASAP7_75t_R _32789_ (.A(_12696_),
    .B(_12519_),
    .Y(_12709_));
 TAPCELL_ASAP7_75t_R PHY_47 ();
 OR3x1_ASAP7_75t_R _32791_ (.A(_12600_),
    .B(_12618_),
    .C(_12692_),
    .Y(_12711_));
 AOI21x1_ASAP7_75t_R _32792_ (.A1(_12626_),
    .A2(_12711_),
    .B(_12703_),
    .Y(_12712_));
 TAPCELL_ASAP7_75t_R PHY_46 ();
 AND2x2_ASAP7_75t_R _32794_ (.A(net297),
    .B(_12685_),
    .Y(_12714_));
 OR3x1_ASAP7_75t_R _32795_ (.A(_12609_),
    .B(_12712_),
    .C(_12714_),
    .Y(_12715_));
 OA211x2_ASAP7_75t_R _32796_ (.A1(_12600_),
    .A2(_12707_),
    .B(_12709_),
    .C(_12715_),
    .Y(_12716_));
 OR3x1_ASAP7_75t_R _32797_ (.A(_09270_),
    .B(_12706_),
    .C(_12716_),
    .Y(_12717_));
 OA21x2_ASAP7_75t_R _32798_ (.A1(_12681_),
    .A2(_09257_),
    .B(_12717_),
    .Y(_04370_));
 TAPCELL_ASAP7_75t_R PHY_45 ();
 TAPCELL_ASAP7_75t_R PHY_44 ();
 AND3x1_ASAP7_75t_R _32801_ (.A(_12682_),
    .B(net297),
    .C(_12626_),
    .Y(_12720_));
 TAPCELL_ASAP7_75t_R PHY_43 ();
 OA211x2_ASAP7_75t_R _32803_ (.A1(_12609_),
    .A2(_12720_),
    .B(_09257_),
    .C(_12696_),
    .Y(_12722_));
 AOI21x1_ASAP7_75t_R _32804_ (.A1(_01746_),
    .A2(_09270_),
    .B(_12722_),
    .Y(_04471_));
 AOI21x1_ASAP7_75t_R _32805_ (.A1(net414),
    .A2(_12606_),
    .B(_12608_),
    .Y(_12723_));
 AND3x4_ASAP7_75t_R _32806_ (.A(_12723_),
    .B(_12699_),
    .C(_12626_),
    .Y(_12724_));
 TAPCELL_ASAP7_75t_R PHY_42 ();
 AND3x2_ASAP7_75t_R _32808_ (.A(_12585_),
    .B(_12592_),
    .C(_12600_),
    .Y(_12726_));
 AND2x4_ASAP7_75t_R _32809_ (.A(_12724_),
    .B(_12726_),
    .Y(_12727_));
 NAND2x1_ASAP7_75t_R _32810_ (.A(_12510_),
    .B(_12727_),
    .Y(_12728_));
 OA21x2_ASAP7_75t_R _32811_ (.A1(_12510_),
    .A2(_12701_),
    .B(_12728_),
    .Y(_12729_));
 OR3x1_ASAP7_75t_R _32812_ (.A(_09270_),
    .B(_12519_),
    .C(_12729_),
    .Y(_12730_));
 OA21x2_ASAP7_75t_R _32813_ (.A1(_13272_),
    .A2(_09257_),
    .B(_12730_),
    .Y(_04472_));
 INVx1_ASAP7_75t_R _32814_ (.A(_12702_),
    .Y(_12731_));
 NAND2x2_ASAP7_75t_R _32815_ (.A(_12571_),
    .B(_12731_),
    .Y(_12732_));
 AND2x4_ASAP7_75t_R _32816_ (.A(_12609_),
    .B(net297),
    .Y(_12733_));
 AO221x1_ASAP7_75t_R _32817_ (.A1(_12527_),
    .A2(_12727_),
    .B1(_12732_),
    .B2(_12693_),
    .C(_12733_),
    .Y(_12734_));
 TAPCELL_ASAP7_75t_R PHY_41 ();
 NOR2x2_ASAP7_75t_R _32819_ (.A(_12541_),
    .B(_12691_),
    .Y(_12736_));
 AND2x2_ASAP7_75t_R _32820_ (.A(_12724_),
    .B(_12736_),
    .Y(_12737_));
 NOR2x2_ASAP7_75t_R _32821_ (.A(_12688_),
    .B(_12703_),
    .Y(_12738_));
 INVx1_ASAP7_75t_R _32822_ (.A(_12738_),
    .Y(_12739_));
 AO21x2_ASAP7_75t_R _32823_ (.A1(net297),
    .A2(_12626_),
    .B(_12609_),
    .Y(_12740_));
 NAND2x2_ASAP7_75t_R _32824_ (.A(_12696_),
    .B(net296),
    .Y(_12741_));
 AND2x2_ASAP7_75t_R _32825_ (.A(_12519_),
    .B(_12741_),
    .Y(_12742_));
 AO21x2_ASAP7_75t_R _32826_ (.A1(_12697_),
    .A2(_12740_),
    .B(_12742_),
    .Y(_12743_));
 AO32x1_ASAP7_75t_R _32827_ (.A1(_12709_),
    .A2(_12737_),
    .A3(_12739_),
    .B1(_12743_),
    .B2(_12527_),
    .Y(_12744_));
 AO21x1_ASAP7_75t_R _32828_ (.A1(_12683_),
    .A2(_12734_),
    .B(_12744_),
    .Y(_12745_));
 OR2x2_ASAP7_75t_R _32829_ (.A(_09270_),
    .B(_12745_),
    .Y(_12746_));
 OA21x2_ASAP7_75t_R _32830_ (.A1(_13271_),
    .A2(_09257_),
    .B(_12746_),
    .Y(_04473_));
 AND3x1_ASAP7_75t_R _32831_ (.A(_12683_),
    .B(_12700_),
    .C(_12726_),
    .Y(_12747_));
 OR2x2_ASAP7_75t_R _32832_ (.A(_12743_),
    .B(_12747_),
    .Y(_12748_));
 AO221x1_ASAP7_75t_R _32833_ (.A1(_12683_),
    .A2(_12733_),
    .B1(_12748_),
    .B2(_12534_),
    .C(_09270_),
    .Y(_12749_));
 OA21x2_ASAP7_75t_R _32834_ (.A1(_13256_),
    .A2(_09257_),
    .B(_12749_),
    .Y(_04474_));
 NAND2x1_ASAP7_75t_R _32835_ (.A(_12626_),
    .B(_12726_),
    .Y(_12750_));
 AND2x6_ASAP7_75t_R _32836_ (.A(_12618_),
    .B(_12626_),
    .Y(_12751_));
 OR2x2_ASAP7_75t_R _32837_ (.A(_12733_),
    .B(_12751_),
    .Y(_12752_));
 INVx1_ASAP7_75t_R _32838_ (.A(_12752_),
    .Y(_12753_));
 TAPCELL_ASAP7_75t_R PHY_40 ();
 OA211x2_ASAP7_75t_R _32840_ (.A1(_12541_),
    .A2(_12750_),
    .B(_12753_),
    .C(_12683_),
    .Y(_12755_));
 AND2x2_ASAP7_75t_R _32841_ (.A(net296),
    .B(_12685_),
    .Y(_12756_));
 TAPCELL_ASAP7_75t_R PHY_39 ();
 NAND2x2_ASAP7_75t_R _32843_ (.A(net296),
    .B(_12618_),
    .Y(_12758_));
 AND3x1_ASAP7_75t_R _32844_ (.A(_12697_),
    .B(_12756_),
    .C(_12758_),
    .Y(_12759_));
 AO21x1_ASAP7_75t_R _32845_ (.A1(_12697_),
    .A2(_12758_),
    .B(_12631_),
    .Y(_12760_));
 OA21x2_ASAP7_75t_R _32846_ (.A1(_12541_),
    .A2(_12759_),
    .B(_12760_),
    .Y(_12761_));
 TAPCELL_ASAP7_75t_R PHY_38 ();
 OR3x1_ASAP7_75t_R _32848_ (.A(_12685_),
    .B(_12691_),
    .C(_12738_),
    .Y(_12763_));
 AO21x1_ASAP7_75t_R _32849_ (.A1(net296),
    .A2(_12763_),
    .B(_12541_),
    .Y(_12764_));
 AND3x1_ASAP7_75t_R _32850_ (.A(_12709_),
    .B(_12758_),
    .C(_12764_),
    .Y(_12765_));
 OR4x1_ASAP7_75t_R _32851_ (.A(_09270_),
    .B(_12755_),
    .C(_12761_),
    .D(_12765_),
    .Y(_12766_));
 OA21x2_ASAP7_75t_R _32852_ (.A1(_13273_),
    .A2(_09257_),
    .B(_12766_),
    .Y(_04475_));
 AND2x4_ASAP7_75t_R _32853_ (.A(_12693_),
    .B(_12732_),
    .Y(_12767_));
 AND2x4_ASAP7_75t_R _32854_ (.A(_12585_),
    .B(_12592_),
    .Y(_12768_));
 OA211x2_ASAP7_75t_R _32855_ (.A1(_12548_),
    .A2(_12688_),
    .B(_12724_),
    .C(_12768_),
    .Y(_12769_));
 OR3x1_ASAP7_75t_R _32856_ (.A(_12767_),
    .B(_12752_),
    .C(_12769_),
    .Y(_12770_));
 NAND2x2_ASAP7_75t_R _32857_ (.A(net296),
    .B(_12685_),
    .Y(_12771_));
 AO22x1_ASAP7_75t_R _32858_ (.A1(_12548_),
    .A2(_12631_),
    .B1(_12771_),
    .B2(_12696_),
    .Y(_12772_));
 TAPCELL_ASAP7_75t_R PHY_37 ();
 NAND2x1_ASAP7_75t_R _32860_ (.A(_12682_),
    .B(net297),
    .Y(_12774_));
 AO21x1_ASAP7_75t_R _32861_ (.A1(net296),
    .A2(_12774_),
    .B(_12548_),
    .Y(_12775_));
 AO221x1_ASAP7_75t_R _32862_ (.A1(_12683_),
    .A2(_12770_),
    .B1(_12772_),
    .B2(_12775_),
    .C(_09270_),
    .Y(_12776_));
 OA21x2_ASAP7_75t_R _32863_ (.A1(_13238_),
    .A2(_09257_),
    .B(_12776_),
    .Y(_04476_));
 NAND2x1_ASAP7_75t_R _32864_ (.A(_12510_),
    .B(_12682_),
    .Y(_12777_));
 TAPCELL_ASAP7_75t_R PHY_36 ();
 AO21x1_ASAP7_75t_R _32866_ (.A1(_12682_),
    .A2(_12740_),
    .B(_12510_),
    .Y(_12779_));
 OA211x2_ASAP7_75t_R _32867_ (.A1(_12777_),
    .A2(_12727_),
    .B(_12779_),
    .C(_12555_),
    .Y(_12780_));
 AO21x1_ASAP7_75t_R _32868_ (.A1(_12555_),
    .A2(_12609_),
    .B(_12737_),
    .Y(_12781_));
 AO22x1_ASAP7_75t_R _32869_ (.A1(_12683_),
    .A2(_12752_),
    .B1(_12781_),
    .B2(_12709_),
    .Y(_12782_));
 OR3x1_ASAP7_75t_R _32870_ (.A(_09270_),
    .B(_12780_),
    .C(_12782_),
    .Y(_12783_));
 OA21x2_ASAP7_75t_R _32871_ (.A1(_13255_),
    .A2(_09257_),
    .B(_12783_),
    .Y(_04477_));
 TAPCELL_ASAP7_75t_R PHY_35 ();
 AO21x1_ASAP7_75t_R _32873_ (.A1(_12696_),
    .A2(_12724_),
    .B(_12562_),
    .Y(_12785_));
 AND3x1_ASAP7_75t_R _32874_ (.A(_12600_),
    .B(_12736_),
    .C(_12703_),
    .Y(_12786_));
 AO21x1_ASAP7_75t_R _32875_ (.A1(_12562_),
    .A2(_12692_),
    .B(_12786_),
    .Y(_12787_));
 TAPCELL_ASAP7_75t_R PHY_34 ();
 OR3x1_ASAP7_75t_R _32877_ (.A(_12510_),
    .B(_12609_),
    .C(_12685_),
    .Y(_12789_));
 AO21x1_ASAP7_75t_R _32878_ (.A1(net297),
    .A2(_12787_),
    .B(_12789_),
    .Y(_12790_));
 AND3x1_ASAP7_75t_R _32879_ (.A(_12519_),
    .B(_12785_),
    .C(_12790_),
    .Y(_12791_));
 AO32x1_ASAP7_75t_R _32880_ (.A1(_12527_),
    .A2(net296),
    .A3(_12685_),
    .B1(_12740_),
    .B2(_12562_),
    .Y(_12792_));
 AND2x2_ASAP7_75t_R _32881_ (.A(net296),
    .B(_12699_),
    .Y(_12793_));
 OA21x2_ASAP7_75t_R _32882_ (.A1(_12685_),
    .A2(_12793_),
    .B(_12562_),
    .Y(_12794_));
 AO221x1_ASAP7_75t_R _32883_ (.A1(_12609_),
    .A2(_12714_),
    .B1(_12751_),
    .B2(_12600_),
    .C(_12794_),
    .Y(_12795_));
 AO22x1_ASAP7_75t_R _32884_ (.A1(_12697_),
    .A2(_12792_),
    .B1(_12795_),
    .B2(_12683_),
    .Y(_12796_));
 OR3x1_ASAP7_75t_R _32885_ (.A(_09270_),
    .B(_12791_),
    .C(_12796_),
    .Y(_12797_));
 OA21x2_ASAP7_75t_R _32886_ (.A1(_13652_),
    .A2(_09257_),
    .B(_12797_),
    .Y(_04478_));
 AO32x1_ASAP7_75t_R _32887_ (.A1(_12571_),
    .A2(net296),
    .A3(_12699_),
    .B1(_12751_),
    .B2(_12534_),
    .Y(_12798_));
 AO32x1_ASAP7_75t_R _32888_ (.A1(_12534_),
    .A2(net296),
    .A3(_12685_),
    .B1(_12740_),
    .B2(_12571_),
    .Y(_12799_));
 AO32x1_ASAP7_75t_R _32889_ (.A1(_12683_),
    .A2(_12707_),
    .A3(_12798_),
    .B1(_12799_),
    .B2(_12697_),
    .Y(_12800_));
 NAND2x2_ASAP7_75t_R _32890_ (.A(_12609_),
    .B(net297),
    .Y(_12801_));
 AO21x1_ASAP7_75t_R _32891_ (.A1(_12685_),
    .A2(_12801_),
    .B(_12519_),
    .Y(_12802_));
 NAND2x1_ASAP7_75t_R _32892_ (.A(net296),
    .B(_12626_),
    .Y(_12803_));
 AO21x1_ASAP7_75t_R _32893_ (.A1(_12724_),
    .A2(_12692_),
    .B(_12803_),
    .Y(_12804_));
 AO21x1_ASAP7_75t_R _32894_ (.A1(_12519_),
    .A2(_12804_),
    .B(_12510_),
    .Y(_12805_));
 AND3x1_ASAP7_75t_R _32895_ (.A(_12571_),
    .B(_12802_),
    .C(_12805_),
    .Y(_12806_));
 OR3x1_ASAP7_75t_R _32896_ (.A(_09270_),
    .B(_12800_),
    .C(_12806_),
    .Y(_12807_));
 OA21x2_ASAP7_75t_R _32897_ (.A1(_05548_),
    .A2(_09257_),
    .B(_12807_),
    .Y(_04479_));
 OR3x1_ASAP7_75t_R _32898_ (.A(_12618_),
    .B(_12691_),
    .C(_12741_),
    .Y(_12808_));
 OA21x2_ASAP7_75t_R _32899_ (.A1(_12519_),
    .A2(net297),
    .B(_12808_),
    .Y(_12809_));
 OR3x1_ASAP7_75t_R _32900_ (.A(_12541_),
    .B(_12685_),
    .C(_12809_),
    .Y(_12810_));
 AO21x1_ASAP7_75t_R _32901_ (.A1(_12510_),
    .A2(_12801_),
    .B(_12519_),
    .Y(_12811_));
 AO21x1_ASAP7_75t_R _32902_ (.A1(_12682_),
    .A2(_12751_),
    .B(_12579_),
    .Y(_12812_));
 AND3x1_ASAP7_75t_R _32903_ (.A(_12810_),
    .B(_12811_),
    .C(_12812_),
    .Y(_12813_));
 OR2x2_ASAP7_75t_R _32904_ (.A(_12541_),
    .B(_12626_),
    .Y(_12814_));
 OR3x1_ASAP7_75t_R _32905_ (.A(_12555_),
    .B(net297),
    .C(_12685_),
    .Y(_12815_));
 AO21x1_ASAP7_75t_R _32906_ (.A1(_12814_),
    .A2(_12815_),
    .B(_12609_),
    .Y(_12816_));
 OA211x2_ASAP7_75t_R _32907_ (.A1(_12579_),
    .A2(_12701_),
    .B(_12816_),
    .C(_12697_),
    .Y(_12817_));
 OR3x1_ASAP7_75t_R _32908_ (.A(_09270_),
    .B(_12813_),
    .C(_12817_),
    .Y(_12818_));
 OA21x2_ASAP7_75t_R _32909_ (.A1(_13950_),
    .A2(_09257_),
    .B(_12818_),
    .Y(_04480_));
 OR3x1_ASAP7_75t_R _32910_ (.A(_12541_),
    .B(_12686_),
    .C(_12691_),
    .Y(_12819_));
 OA21x2_ASAP7_75t_R _32911_ (.A1(_12519_),
    .A2(_12801_),
    .B(_12510_),
    .Y(_12820_));
 AO21x1_ASAP7_75t_R _32912_ (.A1(_12519_),
    .A2(_12819_),
    .B(_12820_),
    .Y(_12821_));
 OR3x1_ASAP7_75t_R _32913_ (.A(_12510_),
    .B(_12585_),
    .C(_12756_),
    .Y(_12822_));
 OA21x2_ASAP7_75t_R _32914_ (.A1(_12696_),
    .A2(_12724_),
    .B(_12822_),
    .Y(_12823_));
 AO221x1_ASAP7_75t_R _32915_ (.A1(_12585_),
    .A2(_12821_),
    .B1(_12823_),
    .B2(_12682_),
    .C(_09270_),
    .Y(_12824_));
 OA21x2_ASAP7_75t_R _32916_ (.A1(_14021_),
    .A2(_09257_),
    .B(_12824_),
    .Y(_04481_));
 AND3x4_ASAP7_75t_R _32917_ (.A(_12723_),
    .B(_12699_),
    .C(_12685_),
    .Y(_12825_));
 TAPCELL_ASAP7_75t_R PHY_33 ();
 AO21x1_ASAP7_75t_R _32919_ (.A1(_12592_),
    .A2(_12825_),
    .B(_12727_),
    .Y(_12827_));
 AND3x1_ASAP7_75t_R _32920_ (.A(_12696_),
    .B(_12592_),
    .C(_12771_),
    .Y(_12828_));
 AO21x1_ASAP7_75t_R _32921_ (.A1(_12510_),
    .A2(_12827_),
    .B(_12828_),
    .Y(_12829_));
 AO22x1_ASAP7_75t_R _32922_ (.A1(_12519_),
    .A2(_12819_),
    .B1(_12774_),
    .B2(_12510_),
    .Y(_12830_));
 AO221x1_ASAP7_75t_R _32923_ (.A1(_12682_),
    .A2(_12829_),
    .B1(_12830_),
    .B2(_12592_),
    .C(_09270_),
    .Y(_12831_));
 OA21x2_ASAP7_75t_R _32924_ (.A1(_14027_),
    .A2(_09257_),
    .B(_12831_),
    .Y(_04482_));
 AO21x1_ASAP7_75t_R _32925_ (.A1(_12600_),
    .A2(net297),
    .B(_12751_),
    .Y(_12832_));
 NAND2x1_ASAP7_75t_R _32926_ (.A(_12585_),
    .B(_12592_),
    .Y(_12833_));
 AO21x1_ASAP7_75t_R _32927_ (.A1(_12548_),
    .A2(_12555_),
    .B(_12600_),
    .Y(_12834_));
 OR2x2_ASAP7_75t_R _32928_ (.A(_12833_),
    .B(_12834_),
    .Y(_12835_));
 AO221x1_ASAP7_75t_R _32929_ (.A1(_12609_),
    .A2(_12832_),
    .B1(_12835_),
    .B2(_12724_),
    .C(_12519_),
    .Y(_12836_));
 AO21x1_ASAP7_75t_R _32930_ (.A1(_12527_),
    .A2(_12767_),
    .B(_12836_),
    .Y(_12837_));
 OA21x2_ASAP7_75t_R _32931_ (.A1(_12682_),
    .A2(_12600_),
    .B(_12510_),
    .Y(_12838_));
 AND2x2_ASAP7_75t_R _32932_ (.A(_12696_),
    .B(net296),
    .Y(_12839_));
 AND2x2_ASAP7_75t_R _32933_ (.A(_12600_),
    .B(_12609_),
    .Y(_12840_));
 AO21x1_ASAP7_75t_R _32934_ (.A1(_12714_),
    .A2(_12839_),
    .B(_12840_),
    .Y(_12841_));
 OA211x2_ASAP7_75t_R _32935_ (.A1(_12609_),
    .A2(_12720_),
    .B(_12696_),
    .C(_12600_),
    .Y(_12842_));
 AO221x1_ASAP7_75t_R _32936_ (.A1(_12837_),
    .A2(_12838_),
    .B1(_12841_),
    .B2(_12519_),
    .C(_12842_),
    .Y(_12843_));
 NAND2x1_ASAP7_75t_R _32937_ (.A(_00281_),
    .B(_09270_),
    .Y(_12844_));
 OA21x2_ASAP7_75t_R _32938_ (.A1(_09270_),
    .A2(_12843_),
    .B(_12844_),
    .Y(_04483_));
 AO21x1_ASAP7_75t_R _32939_ (.A1(net297),
    .A2(_12840_),
    .B(_12519_),
    .Y(_12845_));
 AO21x1_ASAP7_75t_R _32940_ (.A1(_12555_),
    .A2(_12688_),
    .B(_12840_),
    .Y(_12846_));
 OA211x2_ASAP7_75t_R _32941_ (.A1(_12687_),
    .A2(_12846_),
    .B(_12724_),
    .C(_12592_),
    .Y(_12847_));
 AOI211x1_ASAP7_75t_R _32942_ (.A1(_12534_),
    .A2(_12767_),
    .B(_12845_),
    .C(_12847_),
    .Y(_12848_));
 AO21x1_ASAP7_75t_R _32943_ (.A1(_12519_),
    .A2(net296),
    .B(_12848_),
    .Y(_12849_));
 AO221x1_ASAP7_75t_R _32944_ (.A1(net297),
    .A2(_12839_),
    .B1(_12849_),
    .B2(_12510_),
    .C(_09270_),
    .Y(_12850_));
 OAI21x1_ASAP7_75t_R _32945_ (.A1(_00282_),
    .A2(_09257_),
    .B(_12850_),
    .Y(_04484_));
 AO21x1_ASAP7_75t_R _32946_ (.A1(_12688_),
    .A2(_12690_),
    .B(_12833_),
    .Y(_12851_));
 AO221x1_ASAP7_75t_R _32947_ (.A1(_12541_),
    .A2(_12767_),
    .B1(_12851_),
    .B2(_12724_),
    .C(_12845_),
    .Y(_12852_));
 OA211x2_ASAP7_75t_R _32948_ (.A1(_12682_),
    .A2(_12618_),
    .B(_12852_),
    .C(_12510_),
    .Y(_12853_));
 AND3x1_ASAP7_75t_R _32949_ (.A(_12696_),
    .B(_12609_),
    .C(_12618_),
    .Y(_12854_));
 OR3x1_ASAP7_75t_R _32950_ (.A(_09270_),
    .B(_12853_),
    .C(_12854_),
    .Y(_12855_));
 OA21x2_ASAP7_75t_R _32951_ (.A1(_13325_),
    .A2(_09257_),
    .B(_12855_),
    .Y(_04485_));
 AND2x2_ASAP7_75t_R _32952_ (.A(_12723_),
    .B(_12618_),
    .Y(_12856_));
 AO32x1_ASAP7_75t_R _32953_ (.A1(_12562_),
    .A2(_12697_),
    .A3(_12856_),
    .B1(_12760_),
    .B2(_12626_),
    .Y(_12857_));
 AO21x1_ASAP7_75t_R _32954_ (.A1(_12724_),
    .A2(_12768_),
    .B(_12733_),
    .Y(_12858_));
 AND3x2_ASAP7_75t_R _32955_ (.A(_12548_),
    .B(_12555_),
    .C(_12688_),
    .Y(_12859_));
 AOI21x1_ASAP7_75t_R _32956_ (.A1(_12768_),
    .A2(_12834_),
    .B(_12686_),
    .Y(_12860_));
 OR3x1_ASAP7_75t_R _32957_ (.A(_12825_),
    .B(_12751_),
    .C(_12860_),
    .Y(_12861_));
 AO21x1_ASAP7_75t_R _32958_ (.A1(_12724_),
    .A2(_12859_),
    .B(_12861_),
    .Y(_12862_));
 AO222x2_ASAP7_75t_R _32959_ (.A1(_12548_),
    .A2(_12767_),
    .B1(_12858_),
    .B2(_12600_),
    .C1(_12862_),
    .C2(_12562_),
    .Y(_12863_));
 OA21x2_ASAP7_75t_R _32960_ (.A1(_12600_),
    .A2(_12736_),
    .B(_12724_),
    .Y(_12864_));
 OA21x2_ASAP7_75t_R _32961_ (.A1(_12825_),
    .A2(_12864_),
    .B(_12562_),
    .Y(_12865_));
 AO21x1_ASAP7_75t_R _32962_ (.A1(_12609_),
    .A2(_12626_),
    .B(_12865_),
    .Y(_12866_));
 AO22x1_ASAP7_75t_R _32963_ (.A1(_12683_),
    .A2(_12863_),
    .B1(_12866_),
    .B2(_12709_),
    .Y(_12867_));
 OR3x1_ASAP7_75t_R _32964_ (.A(_09270_),
    .B(_12857_),
    .C(_12867_),
    .Y(_12868_));
 OA21x2_ASAP7_75t_R _32965_ (.A1(net304),
    .A2(_09257_),
    .B(_12868_),
    .Y(_04486_));
 OR3x1_ASAP7_75t_R _32966_ (.A(_12600_),
    .B(_12686_),
    .C(_12736_),
    .Y(_12869_));
 NAND2x1_ASAP7_75t_R _32967_ (.A(net296),
    .B(net297),
    .Y(_12870_));
 AO21x1_ASAP7_75t_R _32968_ (.A1(_12571_),
    .A2(_12869_),
    .B(_12870_),
    .Y(_12871_));
 OA21x2_ASAP7_75t_R _32969_ (.A1(_12571_),
    .A2(_12758_),
    .B(_12682_),
    .Y(_12872_));
 AND2x2_ASAP7_75t_R _32970_ (.A(_00240_),
    .B(net103),
    .Y(_12873_));
 AO21x1_ASAP7_75t_R _32971_ (.A1(_06537_),
    .A2(_12311_),
    .B(_12873_),
    .Y(_12874_));
 NAND2x1_ASAP7_75t_R _32972_ (.A(_06511_),
    .B(_01813_),
    .Y(_12875_));
 OA211x2_ASAP7_75t_R _32973_ (.A1(net96),
    .A2(_06511_),
    .B(_12875_),
    .C(_06528_),
    .Y(_12876_));
 AOI21x1_ASAP7_75t_R _32974_ (.A1(net417),
    .A2(_12874_),
    .B(_12876_),
    .Y(_12877_));
 NAND2x1_ASAP7_75t_R _32975_ (.A(_12740_),
    .B(_12877_),
    .Y(_12878_));
 AO32x1_ASAP7_75t_R _32976_ (.A1(_12519_),
    .A2(net296),
    .A3(_12871_),
    .B1(_12872_),
    .B2(_12878_),
    .Y(_12879_));
 NAND2x1_ASAP7_75t_R _32977_ (.A(_12519_),
    .B(_12877_),
    .Y(_12880_));
 OR3x1_ASAP7_75t_R _32978_ (.A(_12548_),
    .B(_12555_),
    .C(_12600_),
    .Y(_12881_));
 INVx1_ASAP7_75t_R _32979_ (.A(_12877_),
    .Y(_12882_));
 AO32x1_ASAP7_75t_R _32980_ (.A1(_12600_),
    .A2(_12768_),
    .A3(_12882_),
    .B1(_12859_),
    .B2(_12571_),
    .Y(_12883_));
 AND3x1_ASAP7_75t_R _32981_ (.A(_12724_),
    .B(_12881_),
    .C(_12883_),
    .Y(_12884_));
 INVx1_ASAP7_75t_R _32982_ (.A(_12732_),
    .Y(_12885_));
 OA21x2_ASAP7_75t_R _32983_ (.A1(_12555_),
    .A2(_12885_),
    .B(_12693_),
    .Y(_12886_));
 OR3x1_ASAP7_75t_R _32984_ (.A(_12845_),
    .B(_12884_),
    .C(_12886_),
    .Y(_12887_));
 AO21x1_ASAP7_75t_R _32985_ (.A1(_12571_),
    .A2(_12861_),
    .B(_12887_),
    .Y(_12888_));
 AO22x1_ASAP7_75t_R _32986_ (.A1(_12519_),
    .A2(_12871_),
    .B1(_12888_),
    .B2(_12510_),
    .Y(_12889_));
 AO221x1_ASAP7_75t_R _32987_ (.A1(_12696_),
    .A2(_12879_),
    .B1(_12880_),
    .B2(_12889_),
    .C(_09270_),
    .Y(_12890_));
 OA21x2_ASAP7_75t_R _32988_ (.A1(_13433_),
    .A2(_09257_),
    .B(_12890_),
    .Y(_04487_));
 NAND2x1_ASAP7_75t_R _32989_ (.A(_06511_),
    .B(_01812_),
    .Y(_12891_));
 OA21x2_ASAP7_75t_R _32990_ (.A1(net107),
    .A2(_06511_),
    .B(_12891_),
    .Y(_12892_));
 NAND2x1_ASAP7_75t_R _32991_ (.A(_06537_),
    .B(_01829_),
    .Y(_12893_));
 OA211x2_ASAP7_75t_R _32992_ (.A1(_06537_),
    .A2(net104),
    .B(_12893_),
    .C(net416),
    .Y(_12894_));
 AO21x1_ASAP7_75t_R _32993_ (.A1(_06528_),
    .A2(_12892_),
    .B(_12894_),
    .Y(_12895_));
 AO32x1_ASAP7_75t_R _32994_ (.A1(_12579_),
    .A2(net296),
    .A3(_12618_),
    .B1(_12740_),
    .B2(_12895_),
    .Y(_12896_));
 AO22x1_ASAP7_75t_R _32995_ (.A1(_12631_),
    .A2(_12895_),
    .B1(_12896_),
    .B2(_12697_),
    .Y(_12897_));
 AO221x1_ASAP7_75t_R _32996_ (.A1(_12579_),
    .A2(_12864_),
    .B1(_12895_),
    .B2(_12609_),
    .C(_12825_),
    .Y(_12898_));
 AND2x2_ASAP7_75t_R _32997_ (.A(_12709_),
    .B(_12898_),
    .Y(_12899_));
 OAI21x1_ASAP7_75t_R _32998_ (.A1(_12767_),
    .A2(_12733_),
    .B(_12600_),
    .Y(_12900_));
 INVx1_ASAP7_75t_R _32999_ (.A(_12900_),
    .Y(_12901_));
 AO21x1_ASAP7_75t_R _33000_ (.A1(_12727_),
    .A2(_12895_),
    .B(_12901_),
    .Y(_12902_));
 OA21x2_ASAP7_75t_R _33001_ (.A1(_12899_),
    .A2(_12902_),
    .B(_12707_),
    .Y(_12903_));
 OA21x2_ASAP7_75t_R _33002_ (.A1(_12862_),
    .A2(_12902_),
    .B(_12683_),
    .Y(_12904_));
 OA22x2_ASAP7_75t_R _33003_ (.A1(_12579_),
    .A2(_12903_),
    .B1(_12904_),
    .B2(_12899_),
    .Y(_12905_));
 OR3x1_ASAP7_75t_R _33004_ (.A(_09270_),
    .B(_12897_),
    .C(_12905_),
    .Y(_12906_));
 OA21x2_ASAP7_75t_R _33005_ (.A1(_13397_),
    .A2(_09257_),
    .B(_12906_),
    .Y(_04488_));
 NAND2x1_ASAP7_75t_R _33006_ (.A(_06511_),
    .B(_01811_),
    .Y(_12907_));
 OA21x2_ASAP7_75t_R _33007_ (.A1(net118),
    .A2(_06511_),
    .B(_12907_),
    .Y(_12908_));
 NAND2x1_ASAP7_75t_R _33008_ (.A(_06537_),
    .B(_01828_),
    .Y(_12909_));
 OA211x2_ASAP7_75t_R _33009_ (.A1(_06537_),
    .A2(net105),
    .B(_12909_),
    .C(net416),
    .Y(_12910_));
 AO21x2_ASAP7_75t_R _33010_ (.A1(_06528_),
    .A2(_12908_),
    .B(_12910_),
    .Y(_12911_));
 AO21x1_ASAP7_75t_R _33011_ (.A1(_12771_),
    .A2(_12911_),
    .B(_12856_),
    .Y(_12912_));
 AO221x1_ASAP7_75t_R _33012_ (.A1(_12585_),
    .A2(_12864_),
    .B1(_12911_),
    .B2(_12609_),
    .C(_12825_),
    .Y(_12913_));
 OA21x2_ASAP7_75t_R _33013_ (.A1(_12750_),
    .A2(_12911_),
    .B(_12793_),
    .Y(_12914_));
 OR3x1_ASAP7_75t_R _33014_ (.A(_12751_),
    .B(_12901_),
    .C(_12914_),
    .Y(_12915_));
 AO22x1_ASAP7_75t_R _33015_ (.A1(_12709_),
    .A2(_12913_),
    .B1(_12915_),
    .B2(_12683_),
    .Y(_12916_));
 OA21x2_ASAP7_75t_R _33016_ (.A1(_12585_),
    .A2(_12707_),
    .B(_12916_),
    .Y(_12917_));
 AO21x1_ASAP7_75t_R _33017_ (.A1(_12519_),
    .A2(_12911_),
    .B(_12917_),
    .Y(_12918_));
 AO222x2_ASAP7_75t_R _33018_ (.A1(_12697_),
    .A2(_12912_),
    .B1(_12917_),
    .B2(_12519_),
    .C1(_12510_),
    .C2(_12918_),
    .Y(_12919_));
 OR2x2_ASAP7_75t_R _33019_ (.A(_09270_),
    .B(_12919_),
    .Y(_12920_));
 OA21x2_ASAP7_75t_R _33020_ (.A1(_13484_),
    .A2(_09257_),
    .B(_12920_),
    .Y(_04489_));
 TAPCELL_ASAP7_75t_R PHY_32 ();
 AND2x2_ASAP7_75t_R _33022_ (.A(_00240_),
    .B(net106),
    .Y(_12922_));
 AO21x1_ASAP7_75t_R _33023_ (.A1(_06537_),
    .A2(_12317_),
    .B(_12922_),
    .Y(_12923_));
 NAND2x1_ASAP7_75t_R _33024_ (.A(_06511_),
    .B(_01810_),
    .Y(_12924_));
 OA211x2_ASAP7_75t_R _33025_ (.A1(net121),
    .A2(_06511_),
    .B(_12924_),
    .C(_06528_),
    .Y(_12925_));
 AO21x1_ASAP7_75t_R _33026_ (.A1(net417),
    .A2(_12923_),
    .B(_12925_),
    .Y(_12926_));
 AO21x1_ASAP7_75t_R _33027_ (.A1(_12697_),
    .A2(_12740_),
    .B(_12631_),
    .Y(_12927_));
 AO221x1_ASAP7_75t_R _33028_ (.A1(_12592_),
    .A2(_12864_),
    .B1(_12926_),
    .B2(_12609_),
    .C(_12825_),
    .Y(_12928_));
 NAND2x1_ASAP7_75t_R _33029_ (.A(_12707_),
    .B(_12900_),
    .Y(_12929_));
 AO21x1_ASAP7_75t_R _33030_ (.A1(_12727_),
    .A2(_12926_),
    .B(_12929_),
    .Y(_12930_));
 AO22x1_ASAP7_75t_R _33031_ (.A1(_12709_),
    .A2(_12928_),
    .B1(_12930_),
    .B2(_12683_),
    .Y(_12931_));
 OR2x2_ASAP7_75t_R _33032_ (.A(_12592_),
    .B(_12707_),
    .Y(_12932_));
 AO221x1_ASAP7_75t_R _33033_ (.A1(_12926_),
    .A2(_12927_),
    .B1(_12931_),
    .B2(_12932_),
    .C(_09270_),
    .Y(_12933_));
 OA21x2_ASAP7_75t_R _33034_ (.A1(_13392_),
    .A2(_09257_),
    .B(_12933_),
    .Y(_04490_));
 AO21x1_ASAP7_75t_R _33035_ (.A1(_12736_),
    .A2(_12738_),
    .B(_12685_),
    .Y(_12934_));
 AO22x1_ASAP7_75t_R _33036_ (.A1(_12527_),
    .A2(_12626_),
    .B1(_12934_),
    .B2(_12699_),
    .Y(_12935_));
 AND2x2_ASAP7_75t_R _33037_ (.A(_00240_),
    .B(net108),
    .Y(_12936_));
 AO21x1_ASAP7_75t_R _33038_ (.A1(_06537_),
    .A2(_12319_),
    .B(_12936_),
    .Y(_12937_));
 TAPCELL_ASAP7_75t_R PHY_31 ();
 NAND2x1_ASAP7_75t_R _33040_ (.A(_06511_),
    .B(_01809_),
    .Y(_12939_));
 OA211x2_ASAP7_75t_R _33041_ (.A1(net122),
    .A2(_06511_),
    .B(_12939_),
    .C(_06528_),
    .Y(_12940_));
 AO21x1_ASAP7_75t_R _33042_ (.A1(net417),
    .A2(_12937_),
    .B(_12940_),
    .Y(_12941_));
 AND2x2_ASAP7_75t_R _33043_ (.A(_12609_),
    .B(_12941_),
    .Y(_12942_));
 AO21x1_ASAP7_75t_R _33044_ (.A1(_12723_),
    .A2(_12935_),
    .B(_12942_),
    .Y(_12943_));
 NAND2x1_ASAP7_75t_R _33045_ (.A(_12600_),
    .B(_12768_),
    .Y(_12944_));
 AND3x2_ASAP7_75t_R _33046_ (.A(net296),
    .B(_12618_),
    .C(_12685_),
    .Y(_12945_));
 AO21x1_ASAP7_75t_R _33047_ (.A1(_12724_),
    .A2(_12944_),
    .B(_12945_),
    .Y(_12946_));
 AO221x1_ASAP7_75t_R _33048_ (.A1(_12727_),
    .A2(_12941_),
    .B1(_12946_),
    .B2(_12527_),
    .C(_12929_),
    .Y(_12947_));
 AO22x1_ASAP7_75t_R _33049_ (.A1(_12709_),
    .A2(_12943_),
    .B1(_12947_),
    .B2(_12683_),
    .Y(_12948_));
 OA21x2_ASAP7_75t_R _33050_ (.A1(_12527_),
    .A2(_12707_),
    .B(_12948_),
    .Y(_12949_));
 AO22x1_ASAP7_75t_R _33051_ (.A1(_12527_),
    .A2(_12856_),
    .B1(_12941_),
    .B2(_12699_),
    .Y(_12950_));
 AO21x1_ASAP7_75t_R _33052_ (.A1(_12626_),
    .A2(_12950_),
    .B(_12942_),
    .Y(_12951_));
 AO22x1_ASAP7_75t_R _33053_ (.A1(_12631_),
    .A2(_12941_),
    .B1(_12951_),
    .B2(_12697_),
    .Y(_12952_));
 OR3x1_ASAP7_75t_R _33054_ (.A(_09270_),
    .B(_12949_),
    .C(_12952_),
    .Y(_12953_));
 OA21x2_ASAP7_75t_R _33055_ (.A1(net309),
    .A2(_09257_),
    .B(_12953_),
    .Y(_04491_));
 AND2x2_ASAP7_75t_R _33056_ (.A(_00240_),
    .B(net109),
    .Y(_12954_));
 AO21x1_ASAP7_75t_R _33057_ (.A1(_06537_),
    .A2(_12321_),
    .B(_12954_),
    .Y(_12955_));
 NAND2x1_ASAP7_75t_R _33058_ (.A(_06511_),
    .B(_01808_),
    .Y(_12956_));
 OA211x2_ASAP7_75t_R _33059_ (.A1(net123),
    .A2(_06511_),
    .B(_12956_),
    .C(_06528_),
    .Y(_12957_));
 AO21x1_ASAP7_75t_R _33060_ (.A1(net416),
    .A2(_12955_),
    .B(_12957_),
    .Y(_12958_));
 OA211x2_ASAP7_75t_R _33061_ (.A1(_12720_),
    .A2(_12741_),
    .B(_12958_),
    .C(_12777_),
    .Y(_12959_));
 AO21x1_ASAP7_75t_R _33062_ (.A1(_12724_),
    .A2(_12859_),
    .B(_12945_),
    .Y(_12960_));
 AND3x2_ASAP7_75t_R _33063_ (.A(_12600_),
    .B(_12693_),
    .C(_12732_),
    .Y(_12961_));
 AO221x1_ASAP7_75t_R _33064_ (.A1(_12727_),
    .A2(_12958_),
    .B1(_12960_),
    .B2(_12534_),
    .C(_12961_),
    .Y(_12962_));
 AO21x1_ASAP7_75t_R _33065_ (.A1(_12519_),
    .A2(_12699_),
    .B(_12751_),
    .Y(_12963_));
 AO21x1_ASAP7_75t_R _33066_ (.A1(_12699_),
    .A2(_12686_),
    .B(_12860_),
    .Y(_12964_));
 AO32x1_ASAP7_75t_R _33067_ (.A1(_12696_),
    .A2(net296),
    .A3(_12963_),
    .B1(_12964_),
    .B2(_12683_),
    .Y(_12965_));
 AO32x1_ASAP7_75t_R _33068_ (.A1(_12683_),
    .A2(_12707_),
    .A3(_12962_),
    .B1(_12965_),
    .B2(_12534_),
    .Y(_12966_));
 OR3x1_ASAP7_75t_R _33069_ (.A(_09270_),
    .B(_12959_),
    .C(_12966_),
    .Y(_12967_));
 OA21x2_ASAP7_75t_R _33070_ (.A1(_13127_),
    .A2(_09257_),
    .B(_12967_),
    .Y(_04492_));
 AND2x2_ASAP7_75t_R _33071_ (.A(_00240_),
    .B(net110),
    .Y(_12968_));
 AO21x1_ASAP7_75t_R _33072_ (.A1(_06537_),
    .A2(_12323_),
    .B(_12968_),
    .Y(_12969_));
 NAND2x1_ASAP7_75t_R _33073_ (.A(_06511_),
    .B(_01807_),
    .Y(_12970_));
 OA211x2_ASAP7_75t_R _33074_ (.A1(net124),
    .A2(_06511_),
    .B(_12970_),
    .C(_06528_),
    .Y(_12971_));
 AO21x2_ASAP7_75t_R _33075_ (.A1(_00662_),
    .A2(_12969_),
    .B(_12971_),
    .Y(_12972_));
 OR3x1_ASAP7_75t_R _33076_ (.A(_12541_),
    .B(net297),
    .C(_12685_),
    .Y(_12973_));
 OA21x2_ASAP7_75t_R _33077_ (.A1(_12555_),
    .A2(_12626_),
    .B(_12973_),
    .Y(_12974_));
 OA21x2_ASAP7_75t_R _33078_ (.A1(_12609_),
    .A2(_12974_),
    .B(_12972_),
    .Y(_12975_));
 AO21x1_ASAP7_75t_R _33079_ (.A1(_12701_),
    .A2(_12974_),
    .B(_12975_),
    .Y(_12976_));
 AO22x1_ASAP7_75t_R _33080_ (.A1(_12631_),
    .A2(_12972_),
    .B1(_12976_),
    .B2(_12697_),
    .Y(_12977_));
 OR3x1_ASAP7_75t_R _33081_ (.A(_12541_),
    .B(_12609_),
    .C(_12714_),
    .Y(_12978_));
 OA211x2_ASAP7_75t_R _33082_ (.A1(net296),
    .A2(_12972_),
    .B(_12978_),
    .C(_12709_),
    .Y(_12979_));
 OR3x1_ASAP7_75t_R _33083_ (.A(_12733_),
    .B(_12756_),
    .C(_12860_),
    .Y(_12980_));
 AO32x1_ASAP7_75t_R _33084_ (.A1(_12600_),
    .A2(_12768_),
    .A3(_12972_),
    .B1(_12859_),
    .B2(_12541_),
    .Y(_12981_));
 AO221x1_ASAP7_75t_R _33085_ (.A1(_12541_),
    .A2(_12980_),
    .B1(_12981_),
    .B2(_12724_),
    .C(_12825_),
    .Y(_12982_));
 OA21x2_ASAP7_75t_R _33086_ (.A1(_12961_),
    .A2(_12982_),
    .B(_12683_),
    .Y(_12983_));
 OA22x2_ASAP7_75t_R _33087_ (.A1(_12541_),
    .A2(_12707_),
    .B1(_12979_),
    .B2(_12983_),
    .Y(_12984_));
 OR3x1_ASAP7_75t_R _33088_ (.A(_09270_),
    .B(_12977_),
    .C(_12984_),
    .Y(_12985_));
 OA21x2_ASAP7_75t_R _33089_ (.A1(_13132_),
    .A2(_09257_),
    .B(_12985_),
    .Y(_04493_));
 NAND2x1_ASAP7_75t_R _33090_ (.A(_06511_),
    .B(_01806_),
    .Y(_12986_));
 OA211x2_ASAP7_75t_R _33091_ (.A1(net125),
    .A2(_06511_),
    .B(_12986_),
    .C(_06528_),
    .Y(_12987_));
 NAND2x1_ASAP7_75t_R _33092_ (.A(_06537_),
    .B(_01823_),
    .Y(_12988_));
 OA211x2_ASAP7_75t_R _33093_ (.A1(_06537_),
    .A2(net111),
    .B(_12988_),
    .C(net417),
    .Y(_12989_));
 OR2x2_ASAP7_75t_R _33094_ (.A(_12987_),
    .B(_12989_),
    .Y(_12990_));
 OAI21x1_ASAP7_75t_R _33095_ (.A1(_12944_),
    .A2(_12990_),
    .B(_12724_),
    .Y(_12991_));
 INVx1_ASAP7_75t_R _33096_ (.A(_12991_),
    .Y(_12992_));
 AO21x1_ASAP7_75t_R _33097_ (.A1(_12768_),
    .A2(_12992_),
    .B(_12548_),
    .Y(_12993_));
 OA21x2_ASAP7_75t_R _33098_ (.A1(_12945_),
    .A2(_12992_),
    .B(_12993_),
    .Y(_12994_));
 OA211x2_ASAP7_75t_R _33099_ (.A1(_12961_),
    .A2(_12994_),
    .B(_12683_),
    .C(_12707_),
    .Y(_12995_));
 OR2x2_ASAP7_75t_R _33100_ (.A(_12548_),
    .B(_12618_),
    .Y(_12996_));
 OA21x2_ASAP7_75t_R _33101_ (.A1(_12585_),
    .A2(_12699_),
    .B(_12996_),
    .Y(_12997_));
 OA21x2_ASAP7_75t_R _33102_ (.A1(_12771_),
    .A2(_12997_),
    .B(_12697_),
    .Y(_12998_));
 AO21x1_ASAP7_75t_R _33103_ (.A1(_12742_),
    .A2(_12990_),
    .B(_12998_),
    .Y(_12999_));
 OA21x2_ASAP7_75t_R _33104_ (.A1(_12701_),
    .A2(_12990_),
    .B(_12999_),
    .Y(_13000_));
 AND3x1_ASAP7_75t_R _33105_ (.A(_12696_),
    .B(_12519_),
    .C(net296),
    .Y(_13001_));
 AND4x1_ASAP7_75t_R _33106_ (.A(_12510_),
    .B(_12682_),
    .C(_12699_),
    .D(_12803_),
    .Y(_13002_));
 OA21x2_ASAP7_75t_R _33107_ (.A1(_13001_),
    .A2(_13002_),
    .B(_12548_),
    .Y(_13003_));
 OR4x1_ASAP7_75t_R _33108_ (.A(_09270_),
    .B(_12995_),
    .C(_13000_),
    .D(_13003_),
    .Y(_13004_));
 OA21x2_ASAP7_75t_R _33109_ (.A1(_13598_),
    .A2(_09257_),
    .B(_13004_),
    .Y(_04494_));
 AND2x2_ASAP7_75t_R _33110_ (.A(_00240_),
    .B(net112),
    .Y(_13005_));
 AO21x1_ASAP7_75t_R _33111_ (.A1(_06537_),
    .A2(_12327_),
    .B(_13005_),
    .Y(_13006_));
 NAND2x1_ASAP7_75t_R _33112_ (.A(_06511_),
    .B(_01805_),
    .Y(_13007_));
 OA211x2_ASAP7_75t_R _33113_ (.A1(net126),
    .A2(_06511_),
    .B(_13007_),
    .C(_06528_),
    .Y(_13008_));
 AO21x2_ASAP7_75t_R _33114_ (.A1(net417),
    .A2(_13006_),
    .B(_13008_),
    .Y(_13009_));
 AO32x1_ASAP7_75t_R _33115_ (.A1(_12592_),
    .A2(net296),
    .A3(_12685_),
    .B1(_12740_),
    .B2(_13009_),
    .Y(_13010_));
 AO22x1_ASAP7_75t_R _33116_ (.A1(_12631_),
    .A2(_13009_),
    .B1(_13010_),
    .B2(_12697_),
    .Y(_13011_));
 AND3x2_ASAP7_75t_R _33117_ (.A(_12571_),
    .B(_12693_),
    .C(_12731_),
    .Y(_13012_));
 OA21x2_ASAP7_75t_R _33118_ (.A1(_12756_),
    .A2(_13012_),
    .B(_12555_),
    .Y(_13013_));
 AO21x1_ASAP7_75t_R _33119_ (.A1(_12555_),
    .A2(_12833_),
    .B(_12803_),
    .Y(_13014_));
 OR2x2_ASAP7_75t_R _33120_ (.A(_12592_),
    .B(net296),
    .Y(_13015_));
 AO32x1_ASAP7_75t_R _33121_ (.A1(_12699_),
    .A2(_13014_),
    .A3(_13015_),
    .B1(_12727_),
    .B2(_13009_),
    .Y(_13016_));
 OR3x1_ASAP7_75t_R _33122_ (.A(_12961_),
    .B(_13013_),
    .C(_13016_),
    .Y(_13017_));
 OR3x1_ASAP7_75t_R _33123_ (.A(_12555_),
    .B(_12609_),
    .C(_12714_),
    .Y(_13018_));
 OA211x2_ASAP7_75t_R _33124_ (.A1(net296),
    .A2(_13009_),
    .B(_13018_),
    .C(_12709_),
    .Y(_13019_));
 AO21x1_ASAP7_75t_R _33125_ (.A1(_12683_),
    .A2(_13017_),
    .B(_13019_),
    .Y(_13020_));
 OA21x2_ASAP7_75t_R _33126_ (.A1(_12555_),
    .A2(_12707_),
    .B(_13020_),
    .Y(_13021_));
 OR3x1_ASAP7_75t_R _33127_ (.A(_09270_),
    .B(_13011_),
    .C(_13021_),
    .Y(_13022_));
 OA21x2_ASAP7_75t_R _33128_ (.A1(_13174_),
    .A2(_09257_),
    .B(_13022_),
    .Y(_04495_));
 OA21x2_ASAP7_75t_R _33129_ (.A1(_12600_),
    .A2(_12707_),
    .B(_12683_),
    .Y(_13023_));
 OA21x2_ASAP7_75t_R _33130_ (.A1(_12752_),
    .A2(_13012_),
    .B(_12527_),
    .Y(_13024_));
 AND2x2_ASAP7_75t_R _33131_ (.A(_00240_),
    .B(net113),
    .Y(_13025_));
 AO21x1_ASAP7_75t_R _33132_ (.A1(_06537_),
    .A2(_12329_),
    .B(_13025_),
    .Y(_13026_));
 NAND2x1_ASAP7_75t_R _33133_ (.A(_06511_),
    .B(_01804_),
    .Y(_13027_));
 OA211x2_ASAP7_75t_R _33134_ (.A1(net127),
    .A2(_06511_),
    .B(_13027_),
    .C(_06528_),
    .Y(_13028_));
 AOI21x1_ASAP7_75t_R _33135_ (.A1(net417),
    .A2(_13026_),
    .B(_13028_),
    .Y(_13029_));
 INVx1_ASAP7_75t_R _33136_ (.A(_13029_),
    .Y(_13030_));
 AND3x2_ASAP7_75t_R _33137_ (.A(_12592_),
    .B(_12600_),
    .C(_12724_),
    .Y(_13031_));
 OA21x2_ASAP7_75t_R _33138_ (.A1(_12687_),
    .A2(_13030_),
    .B(_13031_),
    .Y(_13032_));
 OA21x2_ASAP7_75t_R _33139_ (.A1(_12767_),
    .A2(_12945_),
    .B(_12600_),
    .Y(_13033_));
 OR4x1_ASAP7_75t_R _33140_ (.A(_12825_),
    .B(_13024_),
    .C(_13032_),
    .D(_13033_),
    .Y(_13034_));
 AND2x2_ASAP7_75t_R _33141_ (.A(_12740_),
    .B(_13030_),
    .Y(_13035_));
 AO21x1_ASAP7_75t_R _33142_ (.A1(_12600_),
    .A2(_12701_),
    .B(_13035_),
    .Y(_13036_));
 AND4x1_ASAP7_75t_R _33143_ (.A(_12600_),
    .B(net296),
    .C(_12618_),
    .D(_12709_),
    .Y(_13037_));
 AO221x1_ASAP7_75t_R _33144_ (.A1(_12742_),
    .A2(_13030_),
    .B1(_13036_),
    .B2(_12697_),
    .C(_13037_),
    .Y(_13038_));
 AO21x1_ASAP7_75t_R _33145_ (.A1(_13023_),
    .A2(_13034_),
    .B(_13038_),
    .Y(_13039_));
 NAND2x1_ASAP7_75t_R _33146_ (.A(_01743_),
    .B(_09270_),
    .Y(_13040_));
 OA21x2_ASAP7_75t_R _33147_ (.A1(_09270_),
    .A2(_13039_),
    .B(_13040_),
    .Y(_04496_));
 OR3x1_ASAP7_75t_R _33148_ (.A(_12562_),
    .B(_12618_),
    .C(_12626_),
    .Y(_13041_));
 OA211x2_ASAP7_75t_R _33149_ (.A1(_12548_),
    .A2(net297),
    .B(_13041_),
    .C(_12682_),
    .Y(_13042_));
 AND2x2_ASAP7_75t_R _33150_ (.A(_00240_),
    .B(net114),
    .Y(_13043_));
 AO21x1_ASAP7_75t_R _33151_ (.A1(_06537_),
    .A2(_12331_),
    .B(_13043_),
    .Y(_13044_));
 NAND2x1_ASAP7_75t_R _33152_ (.A(_06511_),
    .B(_01803_),
    .Y(_13045_));
 OA211x2_ASAP7_75t_R _33153_ (.A1(net97),
    .A2(_06511_),
    .B(_13045_),
    .C(_06528_),
    .Y(_13046_));
 AOI21x1_ASAP7_75t_R _33154_ (.A1(net417),
    .A2(_13044_),
    .B(_13046_),
    .Y(_13047_));
 OAI21x1_ASAP7_75t_R _33155_ (.A1(_12519_),
    .A2(_12740_),
    .B(_13047_),
    .Y(_13048_));
 OA211x2_ASAP7_75t_R _33156_ (.A1(_12741_),
    .A2(_13042_),
    .B(_13048_),
    .C(_12777_),
    .Y(_13049_));
 AND2x2_ASAP7_75t_R _33157_ (.A(_12527_),
    .B(_12685_),
    .Y(_13050_));
 AO21x1_ASAP7_75t_R _33158_ (.A1(_12562_),
    .A2(_12626_),
    .B(_13050_),
    .Y(_13051_));
 AND3x1_ASAP7_75t_R _33159_ (.A(_12709_),
    .B(_12856_),
    .C(_13051_),
    .Y(_13052_));
 OA211x2_ASAP7_75t_R _33160_ (.A1(_12767_),
    .A2(_12756_),
    .B(_12600_),
    .C(_12683_),
    .Y(_13053_));
 NAND2x1_ASAP7_75t_R _33161_ (.A(_12585_),
    .B(_13047_),
    .Y(_13054_));
 OA21x2_ASAP7_75t_R _33162_ (.A1(_12751_),
    .A2(_13012_),
    .B(_12548_),
    .Y(_13055_));
 AO221x1_ASAP7_75t_R _33163_ (.A1(_12562_),
    .A2(_12733_),
    .B1(_13031_),
    .B2(_13054_),
    .C(_13055_),
    .Y(_13056_));
 AND3x1_ASAP7_75t_R _33164_ (.A(_12683_),
    .B(_12707_),
    .C(_13056_),
    .Y(_13057_));
 OR5x1_ASAP7_75t_R _33165_ (.A(_09270_),
    .B(_13049_),
    .C(_13052_),
    .D(_13053_),
    .E(_13057_),
    .Y(_13058_));
 OA21x2_ASAP7_75t_R _33166_ (.A1(_14141_),
    .A2(_09257_),
    .B(_13058_),
    .Y(_04497_));
 AND2x2_ASAP7_75t_R _33167_ (.A(_00240_),
    .B(net115),
    .Y(_13059_));
 AO21x1_ASAP7_75t_R _33168_ (.A1(_06537_),
    .A2(_12333_),
    .B(_13059_),
    .Y(_13060_));
 NAND2x1_ASAP7_75t_R _33169_ (.A(_06511_),
    .B(_01802_),
    .Y(_13061_));
 OA211x2_ASAP7_75t_R _33170_ (.A1(net98),
    .A2(_06511_),
    .B(_13061_),
    .C(_06528_),
    .Y(_13062_));
 AO21x2_ASAP7_75t_R _33171_ (.A1(net417),
    .A2(_13060_),
    .B(_13062_),
    .Y(_13063_));
 AO32x1_ASAP7_75t_R _33172_ (.A1(_12571_),
    .A2(_12685_),
    .A3(_12793_),
    .B1(_12740_),
    .B2(_13063_),
    .Y(_13064_));
 AND2x2_ASAP7_75t_R _33173_ (.A(_12534_),
    .B(_12685_),
    .Y(_13065_));
 AO21x1_ASAP7_75t_R _33174_ (.A1(_12571_),
    .A2(_12626_),
    .B(_13065_),
    .Y(_13066_));
 AO221x1_ASAP7_75t_R _33175_ (.A1(_12609_),
    .A2(_13063_),
    .B1(_13066_),
    .B2(_12856_),
    .C(_12682_),
    .Y(_13067_));
 AO22x1_ASAP7_75t_R _33176_ (.A1(_12631_),
    .A2(_13063_),
    .B1(_13067_),
    .B2(_12696_),
    .Y(_13068_));
 OA21x2_ASAP7_75t_R _33177_ (.A1(_12687_),
    .A2(_13063_),
    .B(_13031_),
    .Y(_13069_));
 AO221x1_ASAP7_75t_R _33178_ (.A1(_12555_),
    .A2(_12752_),
    .B1(_13012_),
    .B2(_12534_),
    .C(_13069_),
    .Y(_13070_));
 AND3x1_ASAP7_75t_R _33179_ (.A(_12683_),
    .B(_12707_),
    .C(_13070_),
    .Y(_13071_));
 OA33x2_ASAP7_75t_R _33180_ (.A1(_12510_),
    .A2(_12519_),
    .A3(_13064_),
    .B1(_13068_),
    .B2(_13071_),
    .B3(_13053_),
    .Y(_13072_));
 AND2x2_ASAP7_75t_R _33181_ (.A(_14199_),
    .B(_09270_),
    .Y(_13073_));
 AO21x1_ASAP7_75t_R _33182_ (.A1(_09257_),
    .A2(_13072_),
    .B(_13073_),
    .Y(_04498_));
 AND2x2_ASAP7_75t_R _33183_ (.A(net414),
    .B(net116),
    .Y(_13074_));
 AO21x1_ASAP7_75t_R _33184_ (.A1(_06537_),
    .A2(_12335_),
    .B(_13074_),
    .Y(_13075_));
 NAND2x1_ASAP7_75t_R _33185_ (.A(_06511_),
    .B(_01801_),
    .Y(_13076_));
 OA211x2_ASAP7_75t_R _33186_ (.A1(net99),
    .A2(_06511_),
    .B(_13076_),
    .C(_06528_),
    .Y(_13077_));
 AO21x1_ASAP7_75t_R _33187_ (.A1(net416),
    .A2(_13075_),
    .B(_13077_),
    .Y(_13078_));
 AO32x1_ASAP7_75t_R _33188_ (.A1(_12579_),
    .A2(_12697_),
    .A3(_12825_),
    .B1(_12743_),
    .B2(_13078_),
    .Y(_13079_));
 AO21x1_ASAP7_75t_R _33189_ (.A1(_12579_),
    .A2(_12609_),
    .B(_12756_),
    .Y(_13080_));
 OA21x2_ASAP7_75t_R _33190_ (.A1(_12687_),
    .A2(_13078_),
    .B(_13031_),
    .Y(_13081_));
 AO21x1_ASAP7_75t_R _33191_ (.A1(_12541_),
    .A2(_13012_),
    .B(_13081_),
    .Y(_13082_));
 AO221x1_ASAP7_75t_R _33192_ (.A1(_12600_),
    .A2(_12751_),
    .B1(_13080_),
    .B2(net297),
    .C(_13082_),
    .Y(_13083_));
 OA21x2_ASAP7_75t_R _33193_ (.A1(_13033_),
    .A2(_13083_),
    .B(_13023_),
    .Y(_13084_));
 OR3x1_ASAP7_75t_R _33194_ (.A(_09270_),
    .B(_13079_),
    .C(_13084_),
    .Y(_13085_));
 OA21x2_ASAP7_75t_R _33195_ (.A1(_14318_),
    .A2(_09257_),
    .B(_13085_),
    .Y(_04499_));
 AND2x2_ASAP7_75t_R _33196_ (.A(net414),
    .B(net117),
    .Y(_13086_));
 AO21x1_ASAP7_75t_R _33197_ (.A1(_06537_),
    .A2(_12337_),
    .B(_13086_),
    .Y(_13087_));
 NAND2x1_ASAP7_75t_R _33198_ (.A(_06511_),
    .B(_01800_),
    .Y(_13088_));
 OA211x2_ASAP7_75t_R _33199_ (.A1(net100),
    .A2(_06511_),
    .B(_13088_),
    .C(_06528_),
    .Y(_13089_));
 AO21x1_ASAP7_75t_R _33200_ (.A1(net416),
    .A2(_13087_),
    .B(_13089_),
    .Y(_13090_));
 AO32x1_ASAP7_75t_R _33201_ (.A1(_12585_),
    .A2(_12685_),
    .A3(_12793_),
    .B1(_12740_),
    .B2(_13090_),
    .Y(_13091_));
 AO21x1_ASAP7_75t_R _33202_ (.A1(_12600_),
    .A2(_12618_),
    .B(_12825_),
    .Y(_13092_));
 AO21x1_ASAP7_75t_R _33203_ (.A1(_12585_),
    .A2(_12733_),
    .B(_13092_),
    .Y(_13093_));
 OA21x2_ASAP7_75t_R _33204_ (.A1(_12687_),
    .A2(_13090_),
    .B(_13031_),
    .Y(_13094_));
 OA21x2_ASAP7_75t_R _33205_ (.A1(_13093_),
    .A2(_13094_),
    .B(_13023_),
    .Y(_13095_));
 AO221x1_ASAP7_75t_R _33206_ (.A1(_12742_),
    .A2(_13090_),
    .B1(_13091_),
    .B2(_12697_),
    .C(_13095_),
    .Y(_13096_));
 AND2x2_ASAP7_75t_R _33207_ (.A(_09257_),
    .B(_13096_),
    .Y(_13097_));
 AO21x1_ASAP7_75t_R _33208_ (.A1(_14375_),
    .A2(_09270_),
    .B(_13097_),
    .Y(_04500_));
 AND2x2_ASAP7_75t_R _33209_ (.A(_00240_),
    .B(net119),
    .Y(_13098_));
 AO21x1_ASAP7_75t_R _33210_ (.A1(_06537_),
    .A2(_12339_),
    .B(_13098_),
    .Y(_13099_));
 NAND2x1_ASAP7_75t_R _33211_ (.A(_06511_),
    .B(_01799_),
    .Y(_13100_));
 OA211x2_ASAP7_75t_R _33212_ (.A1(net101),
    .A2(_06511_),
    .B(_13100_),
    .C(_06528_),
    .Y(_13101_));
 AOI21x1_ASAP7_75t_R _33213_ (.A1(net417),
    .A2(_13099_),
    .B(_13101_),
    .Y(_13102_));
 INVx1_ASAP7_75t_R _33214_ (.A(_13102_),
    .Y(_13103_));
 AND2x2_ASAP7_75t_R _33215_ (.A(_12687_),
    .B(_12592_),
    .Y(_13104_));
 AO21x1_ASAP7_75t_R _33216_ (.A1(_12585_),
    .A2(_13103_),
    .B(_13104_),
    .Y(_13105_));
 AOI21x1_ASAP7_75t_R _33217_ (.A1(_12592_),
    .A2(_12881_),
    .B(_12687_),
    .Y(_13106_));
 AO21x1_ASAP7_75t_R _33218_ (.A1(_12600_),
    .A2(_13105_),
    .B(_13106_),
    .Y(_13107_));
 AO221x1_ASAP7_75t_R _33219_ (.A1(_12571_),
    .A2(_12733_),
    .B1(_13107_),
    .B2(_12724_),
    .C(_13092_),
    .Y(_13108_));
 AO221x1_ASAP7_75t_R _33220_ (.A1(_12743_),
    .A2(_13103_),
    .B1(_13108_),
    .B2(_13023_),
    .C(_09270_),
    .Y(_13109_));
 OA21x2_ASAP7_75t_R _33221_ (.A1(_13369_),
    .A2(_09257_),
    .B(_13109_),
    .Y(_04501_));
 AND2x2_ASAP7_75t_R _33222_ (.A(net414),
    .B(net120),
    .Y(_13110_));
 AO21x1_ASAP7_75t_R _33223_ (.A1(_06537_),
    .A2(_12340_),
    .B(_13110_),
    .Y(_13111_));
 NAND2x1_ASAP7_75t_R _33224_ (.A(_06511_),
    .B(_01798_),
    .Y(_13112_));
 OA211x2_ASAP7_75t_R _33225_ (.A1(net102),
    .A2(_06511_),
    .B(_13112_),
    .C(_06528_),
    .Y(_13113_));
 AOI21x1_ASAP7_75t_R _33226_ (.A1(net416),
    .A2(_13111_),
    .B(_13113_),
    .Y(_13114_));
 INVx1_ASAP7_75t_R _33227_ (.A(_13114_),
    .Y(_13115_));
 NAND2x1_ASAP7_75t_R _33228_ (.A(_12585_),
    .B(_13114_),
    .Y(_13116_));
 AO221x1_ASAP7_75t_R _33229_ (.A1(_12600_),
    .A2(_12609_),
    .B1(_13031_),
    .B2(_13116_),
    .C(_13092_),
    .Y(_13117_));
 AO221x1_ASAP7_75t_R _33230_ (.A1(_12743_),
    .A2(_13115_),
    .B1(_13117_),
    .B2(_13023_),
    .C(_09270_),
    .Y(_13118_));
 OA21x2_ASAP7_75t_R _33231_ (.A1(_14597_),
    .A2(_09257_),
    .B(_13118_),
    .Y(_04502_));
 INVx1_ASAP7_75t_R _33232_ (.A(_17871_),
    .Y(_17079_));
 INVx1_ASAP7_75t_R _33233_ (.A(_17763_),
    .Y(_16820_));
 INVx1_ASAP7_75t_R _33234_ (.A(_17787_),
    .Y(_16835_));
 INVx1_ASAP7_75t_R _33235_ (.A(_17767_),
    .Y(_16836_));
 INVx1_ASAP7_75t_R _33236_ (.A(_17786_),
    .Y(_16822_));
 INVx1_ASAP7_75t_R _33237_ (.A(_17805_),
    .Y(_16882_));
 INVx1_ASAP7_75t_R _33238_ (.A(_17785_),
    .Y(_16883_));
 INVx1_ASAP7_75t_R _33239_ (.A(_17783_),
    .Y(_16829_));
 INVx1_ASAP7_75t_R _33240_ (.A(_17766_),
    .Y(_16830_));
 INVx1_ASAP7_75t_R _33241_ (.A(_17764_),
    .Y(_16779_));
 INVx1_ASAP7_75t_R _33242_ (.A(_17782_),
    .Y(_16819_));
 INVx1_ASAP7_75t_R _33243_ (.A(_17830_),
    .Y(_16999_));
 INVx1_ASAP7_75t_R _33244_ (.A(_17858_),
    .Y(_16998_));
 INVx1_ASAP7_75t_R _33245_ (.A(_17730_),
    .Y(_16747_));
 INVx1_ASAP7_75t_R _33246_ (.A(_17748_),
    .Y(_16746_));
 INVx1_ASAP7_75t_R _33247_ (.A(_17820_),
    .Y(_16976_));
 INVx1_ASAP7_75t_R _33248_ (.A(_17852_),
    .Y(_16975_));
 INVx1_ASAP7_75t_R _33249_ (.A(_17821_),
    .Y(_16979_));
 INVx1_ASAP7_75t_R _33250_ (.A(_17848_),
    .Y(_16978_));
 INVx1_ASAP7_75t_R _33251_ (.A(_01362_),
    .Y(_17624_));
 INVx1_ASAP7_75t_R _33252_ (.A(_17825_),
    .Y(_16990_));
 INVx1_ASAP7_75t_R _33253_ (.A(_17854_),
    .Y(_16989_));
 INVx1_ASAP7_75t_R _33254_ (.A(_17804_),
    .Y(_16933_));
 INVx1_ASAP7_75t_R _33255_ (.A(_17826_),
    .Y(_16932_));
 INVx1_ASAP7_75t_R _33256_ (.A(_17731_),
    .Y(_16714_));
 INVx1_ASAP7_75t_R _33257_ (.A(_17827_),
    .Y(_16991_));
 INVx1_ASAP7_75t_R _33258_ (.A(_17828_),
    .Y(_16994_));
 INVx1_ASAP7_75t_R _33259_ (.A(_17857_),
    .Y(_16993_));
 INVx1_ASAP7_75t_R _33260_ (.A(_17788_),
    .Y(_16884_));
 INVx1_ASAP7_75t_R _33261_ (.A(_17781_),
    .Y(_16815_));
 INVx1_ASAP7_75t_R _33262_ (.A(_01367_),
    .Y(_17634_));
 INVx1_ASAP7_75t_R _33263_ (.A(_18000_),
    .Y(_17289_));
 INVx1_ASAP7_75t_R _33264_ (.A(_17982_),
    .Y(_17290_));
 INVx1_ASAP7_75t_R _33265_ (.A(_17977_),
    .Y(_17241_));
 INVx1_ASAP7_75t_R _33266_ (.A(_01428_),
    .Y(_17697_));
 INVx1_ASAP7_75t_R _33267_ (.A(_00010_),
    .Y(_17744_));
 INVx1_ASAP7_75t_R _33268_ (.A(_17768_),
    .Y(_16793_));
 INVx1_ASAP7_75t_R _33269_ (.A(_17750_),
    .Y(_16794_));
 INVx1_ASAP7_75t_R _33270_ (.A(_00066_),
    .Y(_17506_));
 INVx1_ASAP7_75t_R _33271_ (.A(_17956_),
    .Y(_17242_));
 INVx1_ASAP7_75t_R _33272_ (.A(_17942_),
    .Y(_17162_));
 INVx1_ASAP7_75t_R _33273_ (.A(_17917_),
    .Y(_17163_));
 INVx1_ASAP7_75t_R _33274_ (.A(_02297_),
    .Y(_17618_));
 INVx1_ASAP7_75t_R _33275_ (.A(_02298_),
    .Y(_17620_));
 INVx1_ASAP7_75t_R _33276_ (.A(_01361_),
    .Y(_17621_));
 INVx1_ASAP7_75t_R _33277_ (.A(_17939_),
    .Y(_17157_));
 INVx1_ASAP7_75t_R _33278_ (.A(_17915_),
    .Y(_17158_));
 INVx1_ASAP7_75t_R _33279_ (.A(_01435_),
    .Y(_16723_));
 INVx1_ASAP7_75t_R _33280_ (.A(_17809_),
    .Y(_16944_));
 INVx1_ASAP7_75t_R _33281_ (.A(_17831_),
    .Y(_16943_));
 INVx1_ASAP7_75t_R _33282_ (.A(_17806_),
    .Y(_16935_));
 INVx1_ASAP7_75t_R _33283_ (.A(_17834_),
    .Y(_16934_));
 INVx1_ASAP7_75t_R _33284_ (.A(_17807_),
    .Y(_16939_));
 INVx1_ASAP7_75t_R _33285_ (.A(_17829_),
    .Y(_16938_));
 INVx1_ASAP7_75t_R _33286_ (.A(_17811_),
    .Y(_16954_));
 INVx1_ASAP7_75t_R _33287_ (.A(_17837_),
    .Y(_16953_));
 INVx1_ASAP7_75t_R _33288_ (.A(_17813_),
    .Y(_16956_));
 INVx1_ASAP7_75t_R _33289_ (.A(_17835_),
    .Y(_17004_));
 INVx1_ASAP7_75t_R _33290_ (.A(_17863_),
    .Y(_17003_));
 INVx1_ASAP7_75t_R _33291_ (.A(_17836_),
    .Y(_17006_));
 INVx1_ASAP7_75t_R _33292_ (.A(_17862_),
    .Y(_17005_));
 INVx1_ASAP7_75t_R _33293_ (.A(_02340_),
    .Y(_16921_));
 INVx1_ASAP7_75t_R _33294_ (.A(_00022_),
    .Y(_16870_));
 INVx1_ASAP7_75t_R _33295_ (.A(_00021_),
    .Y(_16863_));
 INVx1_ASAP7_75t_R _33296_ (.A(_17721_),
    .Y(_16700_));
 INVx1_ASAP7_75t_R _33297_ (.A(_17981_),
    .Y(_17246_));
 INVx1_ASAP7_75t_R _33298_ (.A(_17958_),
    .Y(_17247_));
 INVx1_ASAP7_75t_R _33299_ (.A(_01363_),
    .Y(_17625_));
 INVx1_ASAP7_75t_R _33300_ (.A(_02296_),
    .Y(_17616_));
 INVx1_ASAP7_75t_R _33301_ (.A(_01359_),
    .Y(_17617_));
 INVx1_ASAP7_75t_R _33302_ (.A(_17943_),
    .Y(_17213_));
 INVx1_ASAP7_75t_R _33303_ (.A(_17967_),
    .Y(_17212_));
 INVx1_ASAP7_75t_R _33304_ (.A(_02295_),
    .Y(_17613_));
 INVx1_ASAP7_75t_R _33305_ (.A(_01358_),
    .Y(_17614_));
 INVx1_ASAP7_75t_R _33306_ (.A(_17983_),
    .Y(_17253_));
 INVx1_ASAP7_75t_R _33307_ (.A(_17962_),
    .Y(_17254_));
 INVx1_ASAP7_75t_R _33308_ (.A(_17961_),
    .Y(_17203_));
 INVx1_ASAP7_75t_R _33309_ (.A(_17937_),
    .Y(_17204_));
 INVx1_ASAP7_75t_R _33310_ (.A(_02333_),
    .Y(_16806_));
 INVx1_ASAP7_75t_R _33311_ (.A(_17913_),
    .Y(_17106_));
 INVx1_ASAP7_75t_R _33312_ (.A(_17889_),
    .Y(_17107_));
 INVx1_ASAP7_75t_R _33313_ (.A(_02351_),
    .Y(_17269_));
 INVx1_ASAP7_75t_R _33314_ (.A(_00048_),
    .Y(_17229_));
 INVx1_ASAP7_75t_R _33315_ (.A(_17914_),
    .Y(_17156_));
 INVx1_ASAP7_75t_R _33316_ (.A(_17940_),
    .Y(_17155_));
 INVx1_ASAP7_75t_R _33317_ (.A(_17936_),
    .Y(_17150_));
 INVx1_ASAP7_75t_R _33318_ (.A(_17912_),
    .Y(_17151_));
 INVx1_ASAP7_75t_R _33319_ (.A(_01365_),
    .Y(_17628_));
 INVx1_ASAP7_75t_R _33320_ (.A(_02300_),
    .Y(_16560_));
 INVx1_ASAP7_75t_R _33321_ (.A(_17339_),
    .Y(_17298_));
 INVx2_ASAP7_75t_R _33322_ (.A(_17301_),
    .Y(_17299_));
 INVx1_ASAP7_75t_R _33323_ (.A(_02294_),
    .Y(_17610_));
 INVx1_ASAP7_75t_R _33324_ (.A(_17957_),
    .Y(_17198_));
 INVx1_ASAP7_75t_R _33325_ (.A(_17935_),
    .Y(_17199_));
 INVx1_ASAP7_75t_R _33326_ (.A(_17997_),
    .Y(_17284_));
 INVx1_ASAP7_75t_R _33327_ (.A(_17979_),
    .Y(_17285_));
 INVx1_ASAP7_75t_R _33328_ (.A(_17998_),
    .Y(_17282_));
 INVx1_ASAP7_75t_R _33329_ (.A(_17978_),
    .Y(_17283_));
 INVx1_ASAP7_75t_R _33330_ (.A(_17994_),
    .Y(_17277_));
 INVx1_ASAP7_75t_R _33331_ (.A(_17976_),
    .Y(_17278_));
 INVx1_ASAP7_75t_R _33332_ (.A(_02308_),
    .Y(_16584_));
 INVx1_ASAP7_75t_R _33333_ (.A(_01373_),
    .Y(_16561_));
 INVx1_ASAP7_75t_R _33334_ (.A(_02302_),
    .Y(_17633_));
 INVx1_ASAP7_75t_R _33335_ (.A(_17824_),
    .Y(_16920_));
 INVx1_ASAP7_75t_R _33336_ (.A(_17867_),
    .Y(_17017_));
 INVx1_ASAP7_75t_R _33337_ (.A(_01400_),
    .Y(_16609_));
 INVx1_ASAP7_75t_R _33338_ (.A(_17776_),
    .Y(_16810_));
 INVx1_ASAP7_75t_R _33339_ (.A(_17757_),
    .Y(_16811_));
 INVx1_ASAP7_75t_R _33340_ (.A(_02332_),
    .Y(_16796_));
 INVx1_ASAP7_75t_R _33341_ (.A(_01440_),
    .Y(_16755_));
 INVx1_ASAP7_75t_R _33342_ (.A(_02331_),
    .Y(_16782_));
 INVx1_ASAP7_75t_R _33343_ (.A(_17842_),
    .Y(_17018_));
 INVx1_ASAP7_75t_R _33344_ (.A(_17789_),
    .Y(_16841_));
 INVx1_ASAP7_75t_R _33345_ (.A(_02311_),
    .Y(_17652_));
 INVx1_ASAP7_75t_R _33346_ (.A(_01380_),
    .Y(_17653_));
 INVx1_ASAP7_75t_R _33347_ (.A(_02304_),
    .Y(_16574_));
 INVx1_ASAP7_75t_R _33348_ (.A(_17955_),
    .Y(_17192_));
 INVx1_ASAP7_75t_R _33349_ (.A(_17931_),
    .Y(_17193_));
 INVx1_ASAP7_75t_R _33350_ (.A(_17796_),
    .Y(_16900_));
 INVx1_ASAP7_75t_R _33351_ (.A(_17812_),
    .Y(_16899_));
 INVx1_ASAP7_75t_R _33352_ (.A(_17801_),
    .Y(_16927_));
 INVx1_ASAP7_75t_R _33353_ (.A(_17823_),
    .Y(_16926_));
 INVx1_ASAP7_75t_R _33354_ (.A(_16565_),
    .Y(_17637_));
 INVx1_ASAP7_75t_R _33355_ (.A(_01414_),
    .Y(_17675_));
 INVx1_ASAP7_75t_R _33356_ (.A(_02319_),
    .Y(_17666_));
 INVx1_ASAP7_75t_R _33357_ (.A(_01401_),
    .Y(_17667_));
 INVx1_ASAP7_75t_R _33358_ (.A(_17792_),
    .Y(_16846_));
 INVx1_ASAP7_75t_R _33359_ (.A(_02321_),
    .Y(_16650_));
 INVx1_ASAP7_75t_R _33360_ (.A(_01405_),
    .Y(_16618_));
 INVx1_ASAP7_75t_R _33361_ (.A(_02316_),
    .Y(_17661_));
 INVx1_ASAP7_75t_R _33362_ (.A(_01392_),
    .Y(_17662_));
 INVx1_ASAP7_75t_R _33363_ (.A(_02306_),
    .Y(_17644_));
 INVx1_ASAP7_75t_R _33364_ (.A(_01371_),
    .Y(_17645_));
 INVx1_ASAP7_75t_R _33365_ (.A(_00242_),
    .Y(_17535_));
 INVx1_ASAP7_75t_R _33366_ (.A(_17522_),
    .Y(_17521_));
 INVx1_ASAP7_75t_R _33367_ (.A(_17841_),
    .Y(_16961_));
 INVx1_ASAP7_75t_R _33368_ (.A(_02345_),
    .Y(_17098_));
 INVx1_ASAP7_75t_R _33369_ (.A(_00035_),
    .Y(_17051_));
 INVx1_ASAP7_75t_R _33370_ (.A(_17815_),
    .Y(_16962_));
 INVx1_ASAP7_75t_R _33371_ (.A(_17799_),
    .Y(_16918_));
 INVx1_ASAP7_75t_R _33372_ (.A(_17819_),
    .Y(_16917_));
 INVx1_ASAP7_75t_R _33373_ (.A(_02299_),
    .Y(_17623_));
 INVx1_ASAP7_75t_R _33374_ (.A(_17929_),
    .Y(_17135_));
 INVx1_ASAP7_75t_R _33375_ (.A(_01430_),
    .Y(_16689_));
 INVx1_ASAP7_75t_R _33376_ (.A(_17905_),
    .Y(_17136_));
 INVx1_ASAP7_75t_R _33377_ (.A(_01369_),
    .Y(_17640_));
 INVx1_ASAP7_75t_R _33378_ (.A(_17897_),
    .Y(_17078_));
 INVx1_ASAP7_75t_R _33379_ (.A(_18057_),
    .Y(_17429_));
 INVx1_ASAP7_75t_R _33380_ (.A(_17904_),
    .Y(_17134_));
 INVx1_ASAP7_75t_R _33381_ (.A(_17671_),
    .Y(_16594_));
 INVx1_ASAP7_75t_R _33382_ (.A(_17658_),
    .Y(_16595_));
 INVx1_ASAP7_75t_R _33383_ (.A(_17678_),
    .Y(_16613_));
 INVx1_ASAP7_75t_R _33384_ (.A(_17670_),
    .Y(_16614_));
 INVx1_ASAP7_75t_R _33385_ (.A(_18005_),
    .Y(_17342_));
 INVx1_ASAP7_75t_R _33386_ (.A(_17907_),
    .Y(_17088_));
 INVx1_ASAP7_75t_R _33387_ (.A(_17784_),
    .Y(_16877_));
 INVx1_ASAP7_75t_R _33388_ (.A(_02325_),
    .Y(_16701_));
 INVx1_ASAP7_75t_R _33389_ (.A(_01424_),
    .Y(_16673_));
 INVx1_ASAP7_75t_R _33390_ (.A(_17740_),
    .Y(_16737_));
 INVx1_ASAP7_75t_R _33391_ (.A(_17720_),
    .Y(_16738_));
 INVx1_ASAP7_75t_R _33392_ (.A(_01381_),
    .Y(_16581_));
 INVx1_ASAP7_75t_R _33393_ (.A(_02312_),
    .Y(_16602_));
 INVx1_ASAP7_75t_R _33394_ (.A(_17954_),
    .Y(_17233_));
 INVx1_ASAP7_75t_R _33395_ (.A(_17973_),
    .Y(_17232_));
 INVx1_ASAP7_75t_R _33396_ (.A(_17875_),
    .Y(_17089_));
 INVx1_ASAP7_75t_R _33397_ (.A(_17741_),
    .Y(_16733_));
 INVx1_ASAP7_75t_R _33398_ (.A(_17719_),
    .Y(_16734_));
 INVx1_ASAP7_75t_R _33399_ (.A(_17756_),
    .Y(_16771_));
 INVx1_ASAP7_75t_R _33400_ (.A(_17739_),
    .Y(_16772_));
 INVx1_ASAP7_75t_R _33401_ (.A(_18080_),
    .Y(_17448_));
 INVx1_ASAP7_75t_R _33402_ (.A(_17758_),
    .Y(_16767_));
 INVx1_ASAP7_75t_R _33403_ (.A(_17738_),
    .Y(_16768_));
 INVx1_ASAP7_75t_R _33404_ (.A(_17502_),
    .Y(_17499_));
 INVx1_ASAP7_75t_R _33405_ (.A(_17524_),
    .Y(_17498_));
 INVx1_ASAP7_75t_R _33406_ (.A(_17816_),
    .Y(_16906_));
 INVx1_ASAP7_75t_R _33407_ (.A(_17817_),
    .Y(_16968_));
 INVx1_ASAP7_75t_R _33408_ (.A(_17843_),
    .Y(_16967_));
 INVx1_ASAP7_75t_R _33409_ (.A(_17851_),
    .Y(_17038_));
 INVx1_ASAP7_75t_R _33410_ (.A(_17847_),
    .Y(_17028_));
 INVx1_ASAP7_75t_R _33411_ (.A(_17872_),
    .Y(_17027_));
 INVx1_ASAP7_75t_R _33412_ (.A(_17765_),
    .Y(_16787_));
 INVx1_ASAP7_75t_R _33413_ (.A(_17932_),
    .Y(_17141_));
 INVx1_ASAP7_75t_R _33414_ (.A(_17910_),
    .Y(_17142_));
 INVx1_ASAP7_75t_R _33415_ (.A(_17749_),
    .Y(_16788_));
 INVx1_ASAP7_75t_R _33416_ (.A(_17906_),
    .Y(_17093_));
 INVx1_ASAP7_75t_R _33417_ (.A(_17880_),
    .Y(_17094_));
 INVx1_ASAP7_75t_R _33418_ (.A(_17879_),
    .Y(_17092_));
 INVx1_ASAP7_75t_R _33419_ (.A(_17850_),
    .Y(_16983_));
 INVx1_ASAP7_75t_R _33420_ (.A(_17822_),
    .Y(_16984_));
 INVx1_ASAP7_75t_R _33421_ (.A(_17882_),
    .Y(_17037_));
 INVx1_ASAP7_75t_R _33422_ (.A(_17876_),
    .Y(_17025_));
 INVx1_ASAP7_75t_R _33423_ (.A(_17846_),
    .Y(_17026_));
 INVx1_ASAP7_75t_R _33424_ (.A(_17845_),
    .Y(_16972_));
 INVx1_ASAP7_75t_R _33425_ (.A(_17818_),
    .Y(_16973_));
 INVx1_ASAP7_75t_R _33426_ (.A(_17707_),
    .Y(_16672_));
 INVx1_ASAP7_75t_R _33427_ (.A(_18026_),
    .Y(_17343_));
 INVx1_ASAP7_75t_R _33428_ (.A(_18006_),
    .Y(_17344_));
 INVx1_ASAP7_75t_R _33429_ (.A(_00011_),
    .Y(_16780_));
 INVx1_ASAP7_75t_R _33430_ (.A(_02334_),
    .Y(_16823_));
 INVx1_ASAP7_75t_R _33431_ (.A(_17869_),
    .Y(_17022_));
 INVx1_ASAP7_75t_R _33432_ (.A(_17844_),
    .Y(_17023_));
 INVx1_ASAP7_75t_R _33433_ (.A(_17505_),
    .Y(_17472_));
 INVx1_ASAP7_75t_R _33434_ (.A(_00018_),
    .Y(_16850_));
 INVx1_ASAP7_75t_R _33435_ (.A(_02338_),
    .Y(_16896_));
 INVx1_ASAP7_75t_R _33436_ (.A(_02324_),
    .Y(_16688_));
 INVx1_ASAP7_75t_R _33437_ (.A(_01421_),
    .Y(_17683_));
 INVx1_ASAP7_75t_R _33438_ (.A(_02328_),
    .Y(_16722_));
 INVx1_ASAP7_75t_R _33439_ (.A(_01429_),
    .Y(_16687_));
 INVx1_ASAP7_75t_R _33440_ (.A(_02337_),
    .Y(_16871_));
 INVx1_ASAP7_75t_R _33441_ (.A(_18081_),
    .Y(_17480_));
 INVx1_ASAP7_75t_R _33442_ (.A(_18090_),
    .Y(_17479_));
 INVx1_ASAP7_75t_R _33443_ (.A(_17802_),
    .Y(_16876_));
 INVx1_ASAP7_75t_R _33444_ (.A(_17711_),
    .Y(_16715_));
 INVx1_ASAP7_75t_R _33445_ (.A(_17732_),
    .Y(_16753_));
 INVx1_ASAP7_75t_R _33446_ (.A(_17751_),
    .Y(_16752_));
 INVx1_ASAP7_75t_R _33447_ (.A(_01408_),
    .Y(_16623_));
 INVx2_ASAP7_75t_R _33448_ (.A(_01419_),
    .Y(_16622_));
 INVx1_ASAP7_75t_R _33449_ (.A(_18084_),
    .Y(_17481_));
 INVx1_ASAP7_75t_R _33450_ (.A(_01431_),
    .Y(_16690_));
 INVx1_ASAP7_75t_R _33451_ (.A(_17769_),
    .Y(_16838_));
 INVx1_ASAP7_75t_R _33452_ (.A(_00043_),
    .Y(_17189_));
 INVx1_ASAP7_75t_R _33453_ (.A(_02339_),
    .Y(_16912_));
 INVx1_ASAP7_75t_R _33454_ (.A(_17700_),
    .Y(_16657_));
 INVx1_ASAP7_75t_R _33455_ (.A(_17684_),
    .Y(_16658_));
 INVx1_ASAP7_75t_R _33456_ (.A(_18082_),
    .Y(_17452_));
 INVx1_ASAP7_75t_R _33457_ (.A(_02320_),
    .Y(_16647_));
 INVx1_ASAP7_75t_R _33458_ (.A(_17903_),
    .Y(_17090_));
 INVx1_ASAP7_75t_R _33459_ (.A(_17877_),
    .Y(_17091_));
 INVx1_ASAP7_75t_R _33460_ (.A(_01403_),
    .Y(_16616_));
 INVx1_ASAP7_75t_R _33461_ (.A(_17870_),
    .Y(_17077_));
 INVx1_ASAP7_75t_R _33462_ (.A(_17901_),
    .Y(_17076_));
 INVx1_ASAP7_75t_R _33463_ (.A(_18100_),
    .Y(_17529_));
 INVx1_ASAP7_75t_R _33464_ (.A(_18102_),
    .Y(_17531_));
 INVx1_ASAP7_75t_R _33465_ (.A(_17523_),
    .Y(_17497_));
 INVx1_ASAP7_75t_R _33466_ (.A(_17849_),
    .Y(_17033_));
 INVx1_ASAP7_75t_R _33467_ (.A(_18031_),
    .Y(_17391_));
 INVx1_ASAP7_75t_R _33468_ (.A(_18052_),
    .Y(_17390_));
 INVx1_ASAP7_75t_R _33469_ (.A(_18012_),
    .Y(_17354_));
 INVx1_ASAP7_75t_R _33470_ (.A(_18030_),
    .Y(_17353_));
 INVx1_ASAP7_75t_R _33471_ (.A(_17874_),
    .Y(_17032_));
 INVx1_ASAP7_75t_R _33472_ (.A(_01378_),
    .Y(_16579_));
 INVx1_ASAP7_75t_R _33473_ (.A(_02310_),
    .Y(_16598_));
 INVx1_ASAP7_75t_R _33474_ (.A(_01415_),
    .Y(_16646_));
 INVx1_ASAP7_75t_R _33475_ (.A(_02323_),
    .Y(_16674_));
 INVx1_ASAP7_75t_R _33476_ (.A(_02327_),
    .Y(_17696_));
 INVx1_ASAP7_75t_R _33477_ (.A(_01423_),
    .Y(_17687_));
 INVx1_ASAP7_75t_R _33478_ (.A(_00014_),
    .Y(_16804_));
 INVx1_ASAP7_75t_R _33479_ (.A(_00017_),
    .Y(_16825_));
 INVx1_ASAP7_75t_R _33480_ (.A(_02335_),
    .Y(_16851_));
 INVx1_ASAP7_75t_R _33481_ (.A(_17853_),
    .Y(_17040_));
 INVx1_ASAP7_75t_R _33482_ (.A(_17878_),
    .Y(_17039_));
 INVx1_ASAP7_75t_R _33483_ (.A(_17941_),
    .Y(_17211_));
 INVx1_ASAP7_75t_R _33484_ (.A(_17963_),
    .Y(_17210_));
 INVx1_ASAP7_75t_R _33485_ (.A(_17984_),
    .Y(_17292_));
 INVx1_ASAP7_75t_R _33486_ (.A(_18004_),
    .Y(_17291_));
 INVx1_ASAP7_75t_R _33487_ (.A(_17959_),
    .Y(_17249_));
 INVx1_ASAP7_75t_R _33488_ (.A(_17980_),
    .Y(_17248_));
 INVx1_ASAP7_75t_R _33489_ (.A(_17770_),
    .Y(_16842_));
 INVx1_ASAP7_75t_R _33490_ (.A(_17985_),
    .Y(_17294_));
 INVx1_ASAP7_75t_R _33491_ (.A(_18003_),
    .Y(_17293_));
 INVx1_ASAP7_75t_R _33492_ (.A(_17938_),
    .Y(_17206_));
 INVx1_ASAP7_75t_R _33493_ (.A(_17960_),
    .Y(_17205_));
 INVx1_ASAP7_75t_R _33494_ (.A(_17775_),
    .Y(_16855_));
 INVx1_ASAP7_75t_R _33495_ (.A(_17795_),
    .Y(_16854_));
 INVx1_ASAP7_75t_R _33496_ (.A(_17944_),
    .Y(_17215_));
 INVx1_ASAP7_75t_R _33497_ (.A(_17966_),
    .Y(_17214_));
 INVx1_ASAP7_75t_R _33498_ (.A(_17893_),
    .Y(_17118_));
 INVx1_ASAP7_75t_R _33499_ (.A(_17918_),
    .Y(_17117_));
 INVx1_ASAP7_75t_R _33500_ (.A(_17919_),
    .Y(_17166_));
 INVx1_ASAP7_75t_R _33501_ (.A(_17948_),
    .Y(_17165_));
 INVx1_ASAP7_75t_R _33502_ (.A(_17946_),
    .Y(_17219_));
 INVx1_ASAP7_75t_R _33503_ (.A(_17685_),
    .Y(_16627_));
 INVx1_ASAP7_75t_R _33504_ (.A(_17864_),
    .Y(_17063_));
 INVx1_ASAP7_75t_R _33505_ (.A(_17890_),
    .Y(_17062_));
 INVx1_ASAP7_75t_R _33506_ (.A(_18014_),
    .Y(_17359_));
 INVx1_ASAP7_75t_R _33507_ (.A(_17891_),
    .Y(_17113_));
 INVx1_ASAP7_75t_R _33508_ (.A(_17916_),
    .Y(_17112_));
 INVx1_ASAP7_75t_R _33509_ (.A(_18034_),
    .Y(_17358_));
 INVx1_ASAP7_75t_R _33510_ (.A(_18018_),
    .Y(_17365_));
 INVx1_ASAP7_75t_R _33511_ (.A(_18035_),
    .Y(_17364_));
 INVx1_ASAP7_75t_R _33512_ (.A(_18036_),
    .Y(_17401_));
 INVx1_ASAP7_75t_R _33513_ (.A(_18056_),
    .Y(_17400_));
 INVx1_ASAP7_75t_R _33514_ (.A(_17771_),
    .Y(_16847_));
 INVx1_ASAP7_75t_R _33515_ (.A(_01366_),
    .Y(_17632_));
 INVx1_ASAP7_75t_R _33516_ (.A(_02301_),
    .Y(_17631_));
 INVx1_ASAP7_75t_R _33517_ (.A(_01372_),
    .Y(_17647_));
 INVx1_ASAP7_75t_R _33518_ (.A(_02307_),
    .Y(_17646_));
 INVx1_ASAP7_75t_R _33519_ (.A(_01368_),
    .Y(_17636_));
 INVx1_ASAP7_75t_R _33520_ (.A(_02303_),
    .Y(_17635_));
 INVx1_ASAP7_75t_R _33521_ (.A(_16564_),
    .Y(_17649_));
 INVx1_ASAP7_75t_R _33522_ (.A(_02309_),
    .Y(_17648_));
 INVx1_ASAP7_75t_R _33523_ (.A(_01370_),
    .Y(_16559_));
 INVx1_ASAP7_75t_R _33524_ (.A(_02305_),
    .Y(_16580_));
 INVx1_ASAP7_75t_R _33525_ (.A(_01418_),
    .Y(_16652_));
 INVx1_ASAP7_75t_R _33526_ (.A(_01425_),
    .Y(_16651_));
 INVx1_ASAP7_75t_R _33527_ (.A(_17920_),
    .Y(_17168_));
 INVx1_ASAP7_75t_R _33528_ (.A(_17945_),
    .Y(_17167_));
 INVx1_ASAP7_75t_R _33529_ (.A(_17964_),
    .Y(_17256_));
 INVx1_ASAP7_75t_R _33530_ (.A(_17987_),
    .Y(_17255_));
 INVx1_ASAP7_75t_R _33531_ (.A(_01416_),
    .Y(_16649_));
 INVx1_ASAP7_75t_R _33532_ (.A(_17752_),
    .Y(_16802_));
 INVx1_ASAP7_75t_R _33533_ (.A(_17772_),
    .Y(_16801_));
 INVx1_ASAP7_75t_R _33534_ (.A(_00040_),
    .Y(_17138_));
 INVx1_ASAP7_75t_R _33535_ (.A(_02348_),
    .Y(_17190_));
 INVx1_ASAP7_75t_R _33536_ (.A(_17988_),
    .Y(_17304_));
 INVx1_ASAP7_75t_R _33537_ (.A(_17715_),
    .Y(_16728_));
 INVx1_ASAP7_75t_R _33538_ (.A(_17735_),
    .Y(_16727_));
 INVx1_ASAP7_75t_R _33539_ (.A(_17922_),
    .Y(_17173_));
 INVx1_ASAP7_75t_R _33540_ (.A(_17947_),
    .Y(_17172_));
 INVx1_ASAP7_75t_R _33541_ (.A(_17949_),
    .Y(_17221_));
 INVx1_ASAP7_75t_R _33542_ (.A(_17968_),
    .Y(_17220_));
 INVx1_ASAP7_75t_R _33543_ (.A(_17965_),
    .Y(_17258_));
 INVx1_ASAP7_75t_R _33544_ (.A(_17986_),
    .Y(_17257_));
 INVx1_ASAP7_75t_R _33545_ (.A(_00037_),
    .Y(_17097_));
 INVx1_ASAP7_75t_R _33546_ (.A(_02346_),
    .Y(_17139_));
 INVx1_ASAP7_75t_R _33547_ (.A(_17989_),
    .Y(_17306_));
 INVx1_ASAP7_75t_R _33548_ (.A(_18007_),
    .Y(_17305_));
 INVx1_ASAP7_75t_R _33549_ (.A(_02343_),
    .Y(_17052_));
 INVx1_ASAP7_75t_R _33550_ (.A(_17703_),
    .Y(_16695_));
 INVx1_ASAP7_75t_R _33551_ (.A(_17716_),
    .Y(_16694_));
 INVx1_ASAP7_75t_R _33552_ (.A(_17999_),
    .Y(_17332_));
 INVx1_ASAP7_75t_R _33553_ (.A(_18019_),
    .Y(_17331_));
 INVx1_ASAP7_75t_R _33554_ (.A(_17699_),
    .Y(_16682_));
 INVx1_ASAP7_75t_R _33555_ (.A(_17712_),
    .Y(_16681_));
 INVx1_ASAP7_75t_R _33556_ (.A(_18064_),
    .Y(_17447_));
 INVx1_ASAP7_75t_R _33557_ (.A(_17969_),
    .Y(_17264_));
 INVx1_ASAP7_75t_R _33558_ (.A(_17733_),
    .Y(_16720_));
 INVx1_ASAP7_75t_R _33559_ (.A(_18001_),
    .Y(_17334_));
 INVx1_ASAP7_75t_R _33560_ (.A(_01434_),
    .Y(_16721_));
 INVx1_ASAP7_75t_R _33561_ (.A(_02329_),
    .Y(_16756_));
 INVx1_ASAP7_75t_R _33562_ (.A(_18023_),
    .Y(_17333_));
 INVx1_ASAP7_75t_R _33563_ (.A(_18062_),
    .Y(_17444_));
 INVx1_ASAP7_75t_R _33564_ (.A(_17475_),
    .Y(_17443_));
 INVx1_ASAP7_75t_R _33565_ (.A(_17898_),
    .Y(_17128_));
 INVx1_ASAP7_75t_R _33566_ (.A(_17923_),
    .Y(_17127_));
 INVx1_ASAP7_75t_R _33567_ (.A(_17925_),
    .Y(_17181_));
 INVx1_ASAP7_75t_R _33568_ (.A(_17950_),
    .Y(_17180_));
 INVx1_ASAP7_75t_R _33569_ (.A(_18047_),
    .Y(_17416_));
 INVx1_ASAP7_75t_R _33570_ (.A(_18063_),
    .Y(_17415_));
 INVx1_ASAP7_75t_R _33571_ (.A(_01393_),
    .Y(_16599_));
 INVx1_ASAP7_75t_R _33572_ (.A(_02317_),
    .Y(_16621_));
 INVx1_ASAP7_75t_R _33573_ (.A(_18065_),
    .Y(_17449_));
 INVx1_ASAP7_75t_R _33574_ (.A(_17780_),
    .Y(_16868_));
 INVx1_ASAP7_75t_R _33575_ (.A(_17800_),
    .Y(_16867_));
 INVx1_ASAP7_75t_R _33576_ (.A(_17970_),
    .Y(_17266_));
 INVx1_ASAP7_75t_R _33577_ (.A(_17990_),
    .Y(_17265_));
 INVx1_ASAP7_75t_R _33578_ (.A(_17993_),
    .Y(_17320_));
 INVx1_ASAP7_75t_R _33579_ (.A(_18013_),
    .Y(_17319_));
 INVx1_ASAP7_75t_R _33580_ (.A(_17995_),
    .Y(_17325_));
 INVx1_ASAP7_75t_R _33581_ (.A(_18017_),
    .Y(_17324_));
 INVx1_ASAP7_75t_R _33582_ (.A(_17996_),
    .Y(_17327_));
 INVx1_ASAP7_75t_R _33583_ (.A(_18016_),
    .Y(_17326_));
 INVx1_ASAP7_75t_R _33584_ (.A(_18058_),
    .Y(_17431_));
 INVx1_ASAP7_75t_R _33585_ (.A(_18074_),
    .Y(_17430_));
 INVx1_ASAP7_75t_R _33586_ (.A(_17803_),
    .Y(_16869_));
 INVx1_ASAP7_75t_R _33587_ (.A(_18060_),
    .Y(_17435_));
 INVx1_ASAP7_75t_R _33588_ (.A(_18076_),
    .Y(_17434_));
 INVx1_ASAP7_75t_R _33589_ (.A(_18002_),
    .Y(_17336_));
 INVx1_ASAP7_75t_R _33590_ (.A(_18022_),
    .Y(_17335_));
 INVx1_ASAP7_75t_R _33591_ (.A(_17474_),
    .Y(_17465_));
 INVx1_ASAP7_75t_R _33592_ (.A(_17873_),
    .Y(_17084_));
 INVx1_ASAP7_75t_R _33593_ (.A(_17899_),
    .Y(_17083_));
 INVx1_ASAP7_75t_R _33594_ (.A(_18079_),
    .Y(_17473_));
 INVx1_ASAP7_75t_R _33595_ (.A(_17900_),
    .Y(_17131_));
 INVx1_ASAP7_75t_R _33596_ (.A(_18089_),
    .Y(_17504_));
 INVx1_ASAP7_75t_R _33597_ (.A(_18097_),
    .Y(_17503_));
 INVx1_ASAP7_75t_R _33598_ (.A(_01412_),
    .Y(_16631_));
 INVx1_ASAP7_75t_R _33599_ (.A(_17734_),
    .Y(_16762_));
 INVx1_ASAP7_75t_R _33600_ (.A(_17753_),
    .Y(_16761_));
 INVx1_ASAP7_75t_R _33601_ (.A(_02349_),
    .Y(_17230_));
 INVx1_ASAP7_75t_R _33602_ (.A(_18091_),
    .Y(_17510_));
 INVx1_ASAP7_75t_R _33603_ (.A(_18099_),
    .Y(_17509_));
 INVx1_ASAP7_75t_R _33604_ (.A(_17902_),
    .Y(_17133_));
 INVx1_ASAP7_75t_R _33605_ (.A(_18049_),
    .Y(_17421_));
 INVx1_ASAP7_75t_R _33606_ (.A(_17926_),
    .Y(_17132_));
 INVx1_ASAP7_75t_R _33607_ (.A(_01390_),
    .Y(_16597_));
 INVx1_ASAP7_75t_R _33608_ (.A(_02315_),
    .Y(_16617_));
 INVx1_ASAP7_75t_R _33609_ (.A(_01406_),
    .Y(_16620_));
 INVx1_ASAP7_75t_R _33610_ (.A(_01417_),
    .Y(_16619_));
 INVx1_ASAP7_75t_R _33611_ (.A(_18067_),
    .Y(_17420_));
 INVx1_ASAP7_75t_R _33612_ (.A(_17868_),
    .Y(_17074_));
 INVx1_ASAP7_75t_R _33613_ (.A(_17894_),
    .Y(_17073_));
 INVx1_ASAP7_75t_R _33614_ (.A(_18068_),
    .Y(_17451_));
 INVx1_ASAP7_75t_R _33615_ (.A(_18083_),
    .Y(_17450_));
 INVx1_ASAP7_75t_R _33616_ (.A(_17895_),
    .Y(_17121_));
 INVx1_ASAP7_75t_R _33617_ (.A(_17692_),
    .Y(_16645_));
 INVx1_ASAP7_75t_R _33618_ (.A(_17924_),
    .Y(_17120_));
 INVx1_ASAP7_75t_R _33619_ (.A(_00023_),
    .Y(_16897_));
 INVx1_ASAP7_75t_R _33620_ (.A(_02341_),
    .Y(_16951_));
 INVx1_ASAP7_75t_R _33621_ (.A(_17927_),
    .Y(_17182_));
 INVx1_ASAP7_75t_R _33622_ (.A(_18029_),
    .Y(_17386_));
 INVx1_ASAP7_75t_R _33623_ (.A(_18048_),
    .Y(_17385_));
 INVx1_ASAP7_75t_R _33624_ (.A(_17991_),
    .Y(_17311_));
 INVx1_ASAP7_75t_R _33625_ (.A(_18009_),
    .Y(_17310_));
 INVx1_ASAP7_75t_R _33626_ (.A(_18050_),
    .Y(_17423_));
 INVx1_ASAP7_75t_R _33627_ (.A(_18066_),
    .Y(_17422_));
 INVx1_ASAP7_75t_R _33628_ (.A(_18069_),
    .Y(_17453_));
 INVx1_ASAP7_75t_R _33629_ (.A(_01399_),
    .Y(_17665_));
 INVx1_ASAP7_75t_R _33630_ (.A(_02318_),
    .Y(_16633_));
 INVx1_ASAP7_75t_R _33631_ (.A(_18085_),
    .Y(_17483_));
 INVx1_ASAP7_75t_R _33632_ (.A(_18092_),
    .Y(_17482_));
 INVx1_ASAP7_75t_R _33633_ (.A(_18093_),
    .Y(_17514_));
 INVx1_ASAP7_75t_R _33634_ (.A(_18101_),
    .Y(_17513_));
 INVx1_ASAP7_75t_R _33635_ (.A(_01413_),
    .Y(_16635_));
 INVx1_ASAP7_75t_R _33636_ (.A(_01422_),
    .Y(_16634_));
 INVx1_ASAP7_75t_R _33637_ (.A(_18098_),
    .Y(_17527_));
 INVx2_ASAP7_75t_R _33638_ (.A(net278),
    .Y(_17338_));
 INVx2_ASAP7_75t_R _33639_ (.A(_17370_),
    .Y(_17337_));
 INVx1_ASAP7_75t_R _33640_ (.A(_17840_),
    .Y(_17012_));
 INVx1_ASAP7_75t_R _33641_ (.A(_17865_),
    .Y(_17011_));
 INVx1_ASAP7_75t_R _33642_ (.A(_17866_),
    .Y(_17069_));
 INVx1_ASAP7_75t_R _33643_ (.A(_17892_),
    .Y(_17068_));
 INVx1_ASAP7_75t_R _33644_ (.A(_18015_),
    .Y(_17361_));
 INVx1_ASAP7_75t_R _33645_ (.A(_18033_),
    .Y(_17360_));
 INVx1_ASAP7_75t_R _33646_ (.A(_18037_),
    .Y(_17403_));
 INVx1_ASAP7_75t_R _33647_ (.A(_18055_),
    .Y(_17402_));
 INVx1_ASAP7_75t_R _33648_ (.A(_18020_),
    .Y(_17367_));
 INVx1_ASAP7_75t_R _33649_ (.A(_18039_),
    .Y(_17366_));
 INVx1_ASAP7_75t_R _33650_ (.A(_18040_),
    .Y(_17404_));
 INVx1_ASAP7_75t_R _33651_ (.A(_18021_),
    .Y(_17369_));
 INVx1_ASAP7_75t_R _33652_ (.A(_18038_),
    .Y(_17368_));
 INVx1_ASAP7_75t_R _33653_ (.A(_18041_),
    .Y(_17406_));
 INVx1_ASAP7_75t_R _33654_ (.A(_18059_),
    .Y(_17405_));
 INVx1_ASAP7_75t_R _33655_ (.A(_18024_),
    .Y(_17371_));
 INVx1_ASAP7_75t_R _33656_ (.A(_18025_),
    .Y(_17373_));
 INVx1_ASAP7_75t_R _33657_ (.A(_18042_),
    .Y(_17372_));
 INVx1_ASAP7_75t_R _33658_ (.A(_18043_),
    .Y(_17410_));
 INVx1_ASAP7_75t_R _33659_ (.A(_18061_),
    .Y(_17409_));
 INVx1_ASAP7_75t_R _33660_ (.A(_18027_),
    .Y(_17377_));
 INVx1_ASAP7_75t_R _33661_ (.A(_18044_),
    .Y(_17376_));
 INVx1_ASAP7_75t_R _33662_ (.A(_17688_),
    .Y(_16667_));
 INVx1_ASAP7_75t_R _33663_ (.A(_17704_),
    .Y(_16666_));
 INVx1_ASAP7_75t_R _33664_ (.A(_17677_),
    .Y(_16640_));
 INVx1_ASAP7_75t_R _33665_ (.A(_17689_),
    .Y(_16639_));
 INVx1_ASAP7_75t_R _33666_ (.A(_18008_),
    .Y(_17348_));
 INVx1_ASAP7_75t_R _33667_ (.A(_18028_),
    .Y(_17347_));
 INVx1_ASAP7_75t_R _33668_ (.A(_17855_),
    .Y(_17041_));
 INVx1_ASAP7_75t_R _33669_ (.A(_17856_),
    .Y(_17043_));
 INVx1_ASAP7_75t_R _33670_ (.A(_17881_),
    .Y(_17042_));
 INVx1_ASAP7_75t_R _33671_ (.A(_17885_),
    .Y(_17101_));
 INVx1_ASAP7_75t_R _33672_ (.A(_17911_),
    .Y(_17100_));
 INVx1_ASAP7_75t_R _33673_ (.A(_17861_),
    .Y(_17055_));
 INVx1_ASAP7_75t_R _33674_ (.A(_17886_),
    .Y(_17054_));
 INVx1_ASAP7_75t_R _33675_ (.A(_17896_),
    .Y(_17123_));
 INVx1_ASAP7_75t_R _33676_ (.A(_17921_),
    .Y(_17122_));
 INVx1_ASAP7_75t_R _33677_ (.A(_18053_),
    .Y(_17426_));
 INVx1_ASAP7_75t_R _33678_ (.A(_18071_),
    .Y(_17425_));
 INVx1_ASAP7_75t_R _33679_ (.A(_17928_),
    .Y(_17184_));
 INVx1_ASAP7_75t_R _33680_ (.A(_17953_),
    .Y(_17183_));
 INVx1_ASAP7_75t_R _33681_ (.A(_18032_),
    .Y(_17393_));
 INVx1_ASAP7_75t_R _33682_ (.A(_18051_),
    .Y(_17392_));
 INVx1_ASAP7_75t_R _33683_ (.A(_17951_),
    .Y(_17222_));
 INVx1_ASAP7_75t_R _33684_ (.A(_17952_),
    .Y(_17224_));
 INVx1_ASAP7_75t_R _33685_ (.A(_17971_),
    .Y(_17223_));
 INVx1_ASAP7_75t_R _33686_ (.A(_18054_),
    .Y(_17428_));
 INVx1_ASAP7_75t_R _33687_ (.A(_18070_),
    .Y(_17427_));
 INVx1_ASAP7_75t_R _33688_ (.A(_17972_),
    .Y(_17272_));
 INVx1_ASAP7_75t_R _33689_ (.A(_17992_),
    .Y(_17271_));
 INVx1_ASAP7_75t_R _33690_ (.A(_18072_),
    .Y(_17454_));
 INVx1_ASAP7_75t_R _33691_ (.A(_18087_),
    .Y(_17487_));
 INVx1_ASAP7_75t_R _33692_ (.A(_18103_),
    .Y(_17516_));
 INVx1_ASAP7_75t_R _33693_ (.A(_18086_),
    .Y(_17455_));
 INVx1_ASAP7_75t_R _33694_ (.A(_18073_),
    .Y(_17456_));
 INVx1_ASAP7_75t_R _33695_ (.A(_18094_),
    .Y(_17486_));
 INVx1_ASAP7_75t_R _33696_ (.A(_17814_),
    .Y(_16902_));
 INVx1_ASAP7_75t_R _33697_ (.A(_17790_),
    .Y(_16888_));
 INVx1_ASAP7_75t_R _33698_ (.A(_17808_),
    .Y(_16887_));
 INVx1_ASAP7_75t_R _33699_ (.A(_00013_),
    .Y(_16783_));
 INVx1_ASAP7_75t_R _33700_ (.A(_17791_),
    .Y(_16893_));
 INVx1_ASAP7_75t_R _33701_ (.A(_17810_),
    .Y(_16892_));
 INVx1_ASAP7_75t_R _33702_ (.A(_01389_),
    .Y(_17656_));
 INVx1_ASAP7_75t_R _33703_ (.A(_02314_),
    .Y(_17655_));
 INVx1_ASAP7_75t_R _33704_ (.A(_01402_),
    .Y(_17668_));
 INVx1_ASAP7_75t_R _33705_ (.A(_17659_),
    .Y(_16573_));
 INVx1_ASAP7_75t_R _33706_ (.A(_01394_),
    .Y(_16601_));
 INVx1_ASAP7_75t_R _33707_ (.A(_01407_),
    .Y(_16600_));
 INVx1_ASAP7_75t_R _33708_ (.A(_01391_),
    .Y(_16577_));
 INVx1_ASAP7_75t_R _33709_ (.A(_01384_),
    .Y(_16586_));
 INVx2_ASAP7_75t_R _33710_ (.A(_01397_),
    .Y(_16585_));
 INVx1_ASAP7_75t_R _33711_ (.A(_01388_),
    .Y(_16590_));
 INVx1_ASAP7_75t_R _33712_ (.A(_01396_),
    .Y(_16604_));
 INVx1_ASAP7_75t_R _33713_ (.A(_01409_),
    .Y(_16603_));
 INVx1_ASAP7_75t_R _33714_ (.A(_00027_),
    .Y(_16913_));
 INVx1_ASAP7_75t_R _33715_ (.A(_01404_),
    .Y(_17674_));
 INVx1_ASAP7_75t_R _33716_ (.A(_01374_),
    .Y(_16563_));
 INVx1_ASAP7_75t_R _33717_ (.A(_01383_),
    .Y(_16562_));
 INVx1_ASAP7_75t_R _33718_ (.A(_01377_),
    .Y(_16569_));
 INVx1_ASAP7_75t_R _33719_ (.A(_00012_),
    .Y(_16781_));
 INVx1_ASAP7_75t_R _33720_ (.A(_18075_),
    .Y(_17460_));
 INVx1_ASAP7_75t_R _33721_ (.A(_18088_),
    .Y(_17459_));
 FAx1_ASAP7_75t_R _33722_ (.SN(\ex_block_i.alu_adder_result_ex_o[1] ),
    .A(_16496_),
    .B(_16497_),
    .CI(_16498_),
    .CON(_02222_));
 FAx1_ASAP7_75t_R _33723_ (.SN(\ex_block_i.alu_adder_result_ex_o[0] ),
    .A(_16500_),
    .B(_16501_),
    .CI(_13781_),
    .CON(_17539_));
 FAx1_ASAP7_75t_R _33724_ (.SN(net174),
    .A(_16504_),
    .B(_16505_),
    .CI(_16506_),
    .CON(_02223_));
 FAx1_ASAP7_75t_R _33725_ (.SN(net176),
    .A(_16507_),
    .B(_16508_),
    .CI(_16509_),
    .CON(_02224_));
 FAx1_ASAP7_75t_R _33726_ (.SN(_00676_),
    .A(_16510_),
    .B(_16511_),
    .CI(_16512_),
    .CON(_00679_));
 FAx1_ASAP7_75t_R _33727_ (.SN(net180),
    .A(_16513_),
    .B(_16514_),
    .CI(_16515_),
    .CON(_02225_));
 FAx1_ASAP7_75t_R _33728_ (.SN(net152),
    .A(_16516_),
    .B(_16517_),
    .CI(_16518_),
    .CON(_02226_));
 FAx1_ASAP7_75t_R _33729_ (.SN(net154),
    .A(_16519_),
    .B(_16520_),
    .CI(_16521_),
    .CON(_02227_));
 FAx1_ASAP7_75t_R _33730_ (.SN(_00785_),
    .A(_16522_),
    .B(_16523_),
    .CI(_16524_),
    .CON(_00818_));
 FAx1_ASAP7_75t_R _33731_ (.SN(net158),
    .A(_16525_),
    .B(_16526_),
    .CI(_16527_),
    .CON(_02228_));
 FAx1_ASAP7_75t_R _33732_ (.SN(net160),
    .A(_16528_),
    .B(_16529_),
    .CI(_16530_),
    .CON(_02229_));
 FAx1_ASAP7_75t_R _33733_ (.SN(net162),
    .A(_16531_),
    .B(_16532_),
    .CI(_16533_),
    .CON(_01014_));
 FAx1_ASAP7_75t_R _33734_ (.SN(net164),
    .A(_16534_),
    .B(_16535_),
    .CI(_16536_),
    .CON(_02230_));
 FAx1_ASAP7_75t_R _33735_ (.SN(net166),
    .A(_16537_),
    .B(_16538_),
    .CI(_16539_),
    .CON(_01145_));
 FAx1_ASAP7_75t_R _33736_ (.SN(net168),
    .A(_16540_),
    .B(_16541_),
    .CI(_16542_),
    .CON(_01211_));
 FAx1_ASAP7_75t_R _33737_ (.SN(net170),
    .A(_16543_),
    .B(_16544_),
    .CI(_16545_),
    .CON(_01277_));
 FAx1_ASAP7_75t_R _33738_ (.SN(_17619_),
    .A(_16546_),
    .B(_16547_),
    .CI(_16548_),
    .CON(_17630_));
 FAx1_ASAP7_75t_R _33739_ (.SN(_17629_),
    .A(_16549_),
    .B(_16550_),
    .CI(_16551_),
    .CON(_17643_));
 FAx1_ASAP7_75t_R _33740_ (.SN(_02231_),
    .A(_16552_),
    .B(_16553_),
    .CI(_16554_),
    .CON(_17650_));
 FAx1_ASAP7_75t_R _33741_ (.SN(_17642_),
    .A(_16556_),
    .B(_16557_),
    .CI(_16558_),
    .CON(_16576_));
 FAx1_ASAP7_75t_R _33742_ (.SN(_01374_),
    .A(_16559_),
    .B(_16560_),
    .CI(_16561_),
    .CON(_01383_));
 FAx1_ASAP7_75t_R _33743_ (.SN(_01376_),
    .A(_16564_),
    .B(_16565_),
    .CI(_16555_),
    .CON(_01387_));
 FAx1_ASAP7_75t_R _33744_ (.SN(_01377_),
    .A(_16566_),
    .B(_16567_),
    .CI(_16568_),
    .CON(_16596_));
 FAx1_ASAP7_75t_R _33745_ (.SN(_16575_),
    .A(_16570_),
    .B(_16571_),
    .CI(_16572_),
    .CON(_17659_));
 FAx1_ASAP7_75t_R _33746_ (.SN(_01379_),
    .A(_16574_),
    .B(_16575_),
    .CI(_16576_),
    .CON(_01391_));
 FAx1_ASAP7_75t_R _33747_ (.SN(_01382_),
    .A(_16579_),
    .B(_16580_),
    .CI(_16581_),
    .CON(_01395_));
 FAx1_ASAP7_75t_R _33748_ (.SN(_01384_),
    .A(_16583_),
    .B(_16562_),
    .CI(_16584_),
    .CON(_01397_));
 FAx1_ASAP7_75t_R _33749_ (.SN(_01388_),
    .A(_16587_),
    .B(_16588_),
    .CI(_16589_),
    .CON(_16615_));
 FAx1_ASAP7_75t_R _33750_ (.SN(_17658_),
    .A(_16591_),
    .B(_16592_),
    .CI(_16593_),
    .CON(_17671_));
 FAx1_ASAP7_75t_R _33751_ (.SN(_17660_),
    .A(_16596_),
    .B(_16595_),
    .CI(_16573_),
    .CON(_17673_));
 FAx1_ASAP7_75t_R _33752_ (.SN(_01394_),
    .A(_16597_),
    .B(_16598_),
    .CI(_16599_),
    .CON(_01407_));
 FAx1_ASAP7_75t_R _33753_ (.SN(_01396_),
    .A(_16601_),
    .B(_16582_),
    .CI(_16602_),
    .CON(_01409_));
 FAx1_ASAP7_75t_R _33754_ (.SN(_02233_),
    .A(_16604_),
    .B(_16585_),
    .CI(_16605_),
    .CON(_02232_));
 FAx1_ASAP7_75t_R _33755_ (.SN(_01400_),
    .A(_16606_),
    .B(_16607_),
    .CI(_16608_),
    .CON(_16641_));
 FAx1_ASAP7_75t_R _33756_ (.SN(_17670_),
    .A(_16610_),
    .B(_16611_),
    .CI(_16612_),
    .CON(_17678_));
 FAx1_ASAP7_75t_R _33757_ (.SN(_17672_),
    .A(_16615_),
    .B(_16614_),
    .CI(_16594_),
    .CON(_17680_));
 FAx1_ASAP7_75t_R _33758_ (.SN(_01406_),
    .A(_16616_),
    .B(_16617_),
    .CI(_16618_),
    .CON(_01417_));
 FAx1_ASAP7_75t_R _33759_ (.SN(_01408_),
    .A(_16620_),
    .B(_16600_),
    .CI(_16621_),
    .CON(_01419_));
 FAx1_ASAP7_75t_R _33760_ (.SN(_16632_),
    .A(_16624_),
    .B(_16625_),
    .CI(_16626_),
    .CON(_17685_));
 FAx1_ASAP7_75t_R _33761_ (.SN(_01412_),
    .A(_16628_),
    .B(_16629_),
    .CI(_16630_),
    .CON(_16668_));
 FAx1_ASAP7_75t_R _33762_ (.SN(_01413_),
    .A(_16632_),
    .B(_16633_),
    .CI(_16631_),
    .CON(_01422_));
 FAx1_ASAP7_75t_R _33763_ (.SN(_17677_),
    .A(_16636_),
    .B(_16637_),
    .CI(_16638_),
    .CON(_17689_));
 FAx1_ASAP7_75t_R _33764_ (.SN(_17679_),
    .A(_16641_),
    .B(_16640_),
    .CI(_16613_),
    .CON(_17691_));
 FAx1_ASAP7_75t_R _33765_ (.SN(_16648_),
    .A(_16642_),
    .B(_16643_),
    .CI(_16644_),
    .CON(_17692_));
 FAx1_ASAP7_75t_R _33766_ (.SN(_01416_),
    .A(_16646_),
    .B(_16647_),
    .CI(_16648_),
    .CON(_16677_));
 FAx1_ASAP7_75t_R _33767_ (.SN(_01418_),
    .A(_16649_),
    .B(_16619_),
    .CI(_16650_),
    .CON(_01425_));
 FAx1_ASAP7_75t_R _33768_ (.SN(_02235_),
    .A(_16652_),
    .B(_16622_),
    .CI(_16653_),
    .CON(_02234_));
 FAx1_ASAP7_75t_R _33769_ (.SN(_17684_),
    .A(_16654_),
    .B(_16655_),
    .CI(_16656_),
    .CON(_17700_));
 FAx1_ASAP7_75t_R _33770_ (.SN(_16662_),
    .A(_16659_),
    .B(_16660_),
    .CI(_16661_),
    .CON(_16696_));
 FAx1_ASAP7_75t_R _33771_ (.SN(_17686_),
    .A(_16658_),
    .B(_16627_),
    .CI(_16662_),
    .CON(_17702_));
 FAx1_ASAP7_75t_R _33772_ (.SN(_17688_),
    .A(_16663_),
    .B(_16664_),
    .CI(_16665_),
    .CON(_17704_));
 FAx1_ASAP7_75t_R _33773_ (.SN(_17690_),
    .A(_16668_),
    .B(_16667_),
    .CI(_16639_),
    .CON(_17706_));
 FAx1_ASAP7_75t_R _33774_ (.SN(_16675_),
    .A(_16669_),
    .B(_16670_),
    .CI(_16671_),
    .CON(_17707_));
 FAx1_ASAP7_75t_R _33775_ (.SN(_16676_),
    .A(_16673_),
    .B(_16674_),
    .CI(_16675_),
    .CON(_16704_));
 FAx1_ASAP7_75t_R _33776_ (.SN(_17693_),
    .A(_16676_),
    .B(_16677_),
    .CI(_16645_),
    .CON(_16706_));
 FAx1_ASAP7_75t_R _33777_ (.SN(_17699_),
    .A(_16678_),
    .B(_16679_),
    .CI(_16680_),
    .CON(_17712_));
 FAx1_ASAP7_75t_R _33778_ (.SN(_16686_),
    .A(_16683_),
    .B(_16684_),
    .CI(_16685_),
    .CON(_16729_));
 FAx1_ASAP7_75t_R _33779_ (.SN(_17701_),
    .A(_16682_),
    .B(_16657_),
    .CI(_16686_),
    .CON(_17714_));
 FAx1_ASAP7_75t_R _33780_ (.SN(_01431_),
    .A(_16687_),
    .B(_16688_),
    .CI(_16689_),
    .CON(_16736_));
 FAx1_ASAP7_75t_R _33781_ (.SN(_17703_),
    .A(_16691_),
    .B(_16692_),
    .CI(_16693_),
    .CON(_17716_));
 FAx1_ASAP7_75t_R _33782_ (.SN(_17705_),
    .A(_16696_),
    .B(_16695_),
    .CI(_16666_),
    .CON(_17718_));
 FAx1_ASAP7_75t_R _33783_ (.SN(_16702_),
    .A(_16697_),
    .B(_16698_),
    .CI(_16699_),
    .CON(_17721_));
 FAx1_ASAP7_75t_R _33784_ (.SN(_16703_),
    .A(_16690_),
    .B(_16701_),
    .CI(_16702_),
    .CON(_16739_));
 FAx1_ASAP7_75t_R _33785_ (.SN(_16705_),
    .A(_16703_),
    .B(_16704_),
    .CI(_16672_),
    .CON(_17723_));
 FAx1_ASAP7_75t_R _33786_ (.SN(_02237_),
    .A(_16705_),
    .B(_16706_),
    .CI(_16707_),
    .CON(_02236_));
 FAx1_ASAP7_75t_R _33787_ (.SN(_17708_),
    .A(_16708_),
    .B(_16709_),
    .CI(_16710_),
    .CON(_17728_));
 FAx1_ASAP7_75t_R _33788_ (.SN(_17711_),
    .A(_16711_),
    .B(_16712_),
    .CI(_16713_),
    .CON(_17731_));
 FAx1_ASAP7_75t_R _33789_ (.SN(_16719_),
    .A(_16716_),
    .B(_16717_),
    .CI(_16718_),
    .CON(_16763_));
 FAx1_ASAP7_75t_R _33790_ (.SN(_17713_),
    .A(_16715_),
    .B(_16681_),
    .CI(_16719_),
    .CON(_17733_));
 FAx1_ASAP7_75t_R _33791_ (.SN(_16735_),
    .A(_16721_),
    .B(_16722_),
    .CI(_16723_),
    .CON(_16770_));
 FAx1_ASAP7_75t_R _33792_ (.SN(_17715_),
    .A(_16724_),
    .B(_16725_),
    .CI(_16726_),
    .CON(_17735_));
 FAx1_ASAP7_75t_R _33793_ (.SN(_17717_),
    .A(_16729_),
    .B(_16728_),
    .CI(_16694_),
    .CON(_17737_));
 FAx1_ASAP7_75t_R _33794_ (.SN(_17719_),
    .A(_16730_),
    .B(_16731_),
    .CI(_16732_),
    .CON(_17741_));
 FAx1_ASAP7_75t_R _33795_ (.SN(_17720_),
    .A(_16735_),
    .B(_16736_),
    .CI(_16734_),
    .CON(_17740_));
 FAx1_ASAP7_75t_R _33796_ (.SN(_17722_),
    .A(_16738_),
    .B(_16739_),
    .CI(_16700_),
    .CON(_16775_));
 FAx1_ASAP7_75t_R _33797_ (.SN(_17727_),
    .A(_16740_),
    .B(_16741_),
    .CI(_16742_),
    .CON(_17747_));
 FAx1_ASAP7_75t_R _33798_ (.SN(_17730_),
    .A(_16743_),
    .B(_16744_),
    .CI(_16745_),
    .CON(_17748_));
 FAx1_ASAP7_75t_R _33799_ (.SN(_16751_),
    .A(_16748_),
    .B(_16749_),
    .CI(_16750_),
    .CON(_16803_));
 FAx1_ASAP7_75t_R _33800_ (.SN(_17732_),
    .A(_16747_),
    .B(_16714_),
    .CI(_16751_),
    .CON(_17751_));
 FAx1_ASAP7_75t_R _33801_ (.SN(_16757_),
    .A(_16754_),
    .B(_16753_),
    .CI(_16720_),
    .CON(_16805_));
 FAx1_ASAP7_75t_R _33802_ (.SN(_16769_),
    .A(_16755_),
    .B(_16756_),
    .CI(_16757_),
    .CON(_16809_));
 FAx1_ASAP7_75t_R _33803_ (.SN(_17734_),
    .A(_16758_),
    .B(_16759_),
    .CI(_16760_),
    .CON(_17753_));
 FAx1_ASAP7_75t_R _33804_ (.SN(_17736_),
    .A(_16763_),
    .B(_16762_),
    .CI(_16727_),
    .CON(_17755_));
 FAx1_ASAP7_75t_R _33805_ (.SN(_17738_),
    .A(_16764_),
    .B(_16765_),
    .CI(_16766_),
    .CON(_17758_));
 FAx1_ASAP7_75t_R _33806_ (.SN(_17739_),
    .A(_16769_),
    .B(_16770_),
    .CI(_16768_),
    .CON(_17756_));
 FAx1_ASAP7_75t_R _33807_ (.SN(_16773_),
    .A(_16772_),
    .B(_16737_),
    .CI(_16733_),
    .CON(_17759_));
 FAx1_ASAP7_75t_R _33808_ (.SN(_02239_),
    .A(_16773_),
    .B(_16774_),
    .CI(_16775_),
    .CON(_02238_));
 FAx1_ASAP7_75t_R _33809_ (.SN(_17746_),
    .A(_16776_),
    .B(_16777_),
    .CI(_16778_),
    .CON(_17764_));
 FAx1_ASAP7_75t_R _33810_ (.SN(_00013_),
    .A(_16780_),
    .B(_16781_),
    .CI(_16782_),
    .CON(_16839_));
 FAx1_ASAP7_75t_R _33811_ (.SN(_17749_),
    .A(_16784_),
    .B(_16785_),
    .CI(_16786_),
    .CON(_17765_));
 FAx1_ASAP7_75t_R _33812_ (.SN(_16792_),
    .A(_16789_),
    .B(_16790_),
    .CI(_16791_),
    .CON(_16848_));
 FAx1_ASAP7_75t_R _33813_ (.SN(_17750_),
    .A(_16746_),
    .B(_16792_),
    .CI(_16788_),
    .CON(_17768_));
 FAx1_ASAP7_75t_R _33814_ (.SN(_16797_),
    .A(_16752_),
    .B(_16795_),
    .CI(_16794_),
    .CON(_16849_));
 FAx1_ASAP7_75t_R _33815_ (.SN(_16808_),
    .A(_16796_),
    .B(_16797_),
    .CI(_16783_),
    .CON(_16852_));
 FAx1_ASAP7_75t_R _33816_ (.SN(_17752_),
    .A(_16798_),
    .B(_16799_),
    .CI(_16800_),
    .CON(_17772_));
 FAx1_ASAP7_75t_R _33817_ (.SN(_17754_),
    .A(_16802_),
    .B(_16803_),
    .CI(_16761_),
    .CON(_17773_));
 FAx1_ASAP7_75t_R _33818_ (.SN(_16807_),
    .A(_16804_),
    .B(_16805_),
    .CI(_16806_),
    .CON(_16856_));
 FAx1_ASAP7_75t_R _33819_ (.SN(_17757_),
    .A(_16807_),
    .B(_16808_),
    .CI(_16809_),
    .CON(_17776_));
 FAx1_ASAP7_75t_R _33820_ (.SN(_17760_),
    .A(_16771_),
    .B(_16767_),
    .CI(_16811_),
    .CON(_16858_));
 FAx1_ASAP7_75t_R _33821_ (.SN(_17762_),
    .A(_16812_),
    .B(_16813_),
    .CI(_16814_),
    .CON(_17781_));
 FAx1_ASAP7_75t_R _33822_ (.SN(_17763_),
    .A(_16816_),
    .B(_16817_),
    .CI(_16818_),
    .CON(_17782_));
 FAx1_ASAP7_75t_R _33823_ (.SN(_16824_),
    .A(_16821_),
    .B(_16779_),
    .CI(_16820_),
    .CON(_17786_));
 FAx1_ASAP7_75t_R _33824_ (.SN(_16840_),
    .A(_16823_),
    .B(_16824_),
    .CI(_16825_),
    .CON(_16885_));
 FAx1_ASAP7_75t_R _33825_ (.SN(_17766_),
    .A(_16826_),
    .B(_16827_),
    .CI(_16828_),
    .CON(_17783_));
 FAx1_ASAP7_75t_R _33826_ (.SN(_16834_),
    .A(_16831_),
    .B(_16832_),
    .CI(_16833_),
    .CON(_16894_));
 FAx1_ASAP7_75t_R _33827_ (.SN(_17767_),
    .A(_16834_),
    .B(_16787_),
    .CI(_16830_),
    .CON(_17787_));
 FAx1_ASAP7_75t_R _33828_ (.SN(_17769_),
    .A(_16836_),
    .B(_16793_),
    .CI(_16837_),
    .CON(_16895_));
 FAx1_ASAP7_75t_R _33829_ (.SN(_17770_),
    .A(_16839_),
    .B(_16838_),
    .CI(_16840_),
    .CON(_17789_));
 FAx1_ASAP7_75t_R _33830_ (.SN(_17771_),
    .A(_16843_),
    .B(_16844_),
    .CI(_16845_),
    .CON(_17792_));
 FAx1_ASAP7_75t_R _33831_ (.SN(_17774_),
    .A(_16848_),
    .B(_16847_),
    .CI(_16801_),
    .CON(_17793_));
 FAx1_ASAP7_75t_R _33832_ (.SN(_16853_),
    .A(_16849_),
    .B(_16850_),
    .CI(_16851_),
    .CON(_16901_));
 FAx1_ASAP7_75t_R _33833_ (.SN(_17775_),
    .A(_16842_),
    .B(_16852_),
    .CI(_16853_),
    .CON(_17795_));
 FAx1_ASAP7_75t_R _33834_ (.SN(_16859_),
    .A(_16855_),
    .B(_16810_),
    .CI(_16856_),
    .CON(_17797_));
 FAx1_ASAP7_75t_R _33835_ (.SN(_02241_),
    .A(_16857_),
    .B(_16858_),
    .CI(_16859_),
    .CON(_02240_));
 FAx1_ASAP7_75t_R _33836_ (.SN(_00021_),
    .A(_16860_),
    .B(_16861_),
    .CI(_16862_),
    .CON(_16919_));
 FAx1_ASAP7_75t_R _33837_ (.SN(_17780_),
    .A(_16864_),
    .B(_16865_),
    .CI(_16866_),
    .CON(_17800_));
 FAx1_ASAP7_75t_R _33838_ (.SN(_16872_),
    .A(_16868_),
    .B(_16819_),
    .CI(_16815_),
    .CON(_17803_));
 FAx1_ASAP7_75t_R _33839_ (.SN(_16886_),
    .A(_16870_),
    .B(_16871_),
    .CI(_16872_),
    .CON(_16936_));
 FAx1_ASAP7_75t_R _33840_ (.SN(_17784_),
    .A(_16873_),
    .B(_16874_),
    .CI(_16875_),
    .CON(_17802_));
 FAx1_ASAP7_75t_R _33841_ (.SN(_16881_),
    .A(_16878_),
    .B(_16879_),
    .CI(_16880_),
    .CON(_16945_));
 FAx1_ASAP7_75t_R _33842_ (.SN(_17785_),
    .A(_16881_),
    .B(_16829_),
    .CI(_16877_),
    .CON(_17805_));
 FAx1_ASAP7_75t_R _33843_ (.SN(_17788_),
    .A(_16835_),
    .B(_16883_),
    .CI(_16822_),
    .CON(_16950_));
 FAx1_ASAP7_75t_R _33844_ (.SN(_17790_),
    .A(_16884_),
    .B(_16885_),
    .CI(_16886_),
    .CON(_17808_));
 FAx1_ASAP7_75t_R _33845_ (.SN(_17791_),
    .A(_16889_),
    .B(_16890_),
    .CI(_16891_),
    .CON(_17810_));
 FAx1_ASAP7_75t_R _33846_ (.SN(_17794_),
    .A(_16893_),
    .B(_16846_),
    .CI(_16894_),
    .CON(_16947_));
 FAx1_ASAP7_75t_R _33847_ (.SN(_16898_),
    .A(_16895_),
    .B(_16896_),
    .CI(_16897_),
    .CON(_16955_));
 FAx1_ASAP7_75t_R _33848_ (.SN(_17796_),
    .A(_16898_),
    .B(_16841_),
    .CI(_16888_),
    .CON(_17812_));
 FAx1_ASAP7_75t_R _33849_ (.SN(_17798_),
    .A(_16901_),
    .B(_16854_),
    .CI(_16900_),
    .CON(_17814_));
 FAx1_ASAP7_75t_R _33850_ (.SN(_16911_),
    .A(_05911_),
    .B(_16904_),
    .CI(_16905_),
    .CON(_17816_));
 FAx1_ASAP7_75t_R _33851_ (.SN(_00026_),
    .A(_16907_),
    .B(_16908_),
    .CI(_16909_),
    .CON(_16974_));
 FAx1_ASAP7_75t_R _33852_ (.SN(_00027_),
    .A(_16911_),
    .B(_16912_),
    .CI(_16910_),
    .CON(_16977_));
 FAx1_ASAP7_75t_R _33853_ (.SN(_17799_),
    .A(_16914_),
    .B(_16915_),
    .CI(_16916_),
    .CON(_17819_));
 FAx1_ASAP7_75t_R _33854_ (.SN(_16922_),
    .A(_16919_),
    .B(_16918_),
    .CI(_16867_),
    .CON(_17824_));
 FAx1_ASAP7_75t_R _33855_ (.SN(_16937_),
    .A(_16913_),
    .B(_16921_),
    .CI(_16922_),
    .CON(_16992_));
 FAx1_ASAP7_75t_R _33856_ (.SN(_17801_),
    .A(_16923_),
    .B(_16924_),
    .CI(_16925_),
    .CON(_17823_));
 FAx1_ASAP7_75t_R _33857_ (.SN(_16931_),
    .A(_16928_),
    .B(_16929_),
    .CI(_16930_),
    .CON(_17000_));
 FAx1_ASAP7_75t_R _33858_ (.SN(_17804_),
    .A(_16927_),
    .B(_16876_),
    .CI(_16931_),
    .CON(_17826_));
 FAx1_ASAP7_75t_R _33859_ (.SN(_17806_),
    .A(_16869_),
    .B(_16933_),
    .CI(_16882_),
    .CON(_17834_));
 FAx1_ASAP7_75t_R _33860_ (.SN(_17807_),
    .A(_16936_),
    .B(_16935_),
    .CI(_16937_),
    .CON(_17829_));
 FAx1_ASAP7_75t_R _33861_ (.SN(_17809_),
    .A(_16940_),
    .B(_16941_),
    .CI(_16942_),
    .CON(_17831_));
 FAx1_ASAP7_75t_R _33862_ (.SN(_16946_),
    .A(_16945_),
    .B(_16944_),
    .CI(_16892_),
    .CON(_17833_));
 FAx1_ASAP7_75t_R _33863_ (.SN(_00028_),
    .A(_16946_),
    .B(_16947_),
    .CI(_16948_),
    .CON(_17002_));
 FAx1_ASAP7_75t_R _33864_ (.SN(_16952_),
    .A(_16950_),
    .B(_16949_),
    .CI(_16951_),
    .CON(_17007_));
 FAx1_ASAP7_75t_R _33865_ (.SN(_17811_),
    .A(_16939_),
    .B(_16887_),
    .CI(_16952_),
    .CON(_17837_));
 FAx1_ASAP7_75t_R _33866_ (.SN(_17813_),
    .A(_16954_),
    .B(_16899_),
    .CI(_16955_),
    .CON(_17839_));
 FAx1_ASAP7_75t_R _33867_ (.SN(_00030_),
    .A(_16956_),
    .B(_16902_),
    .CI(_16957_),
    .CON(_00033_));
 FAx1_ASAP7_75t_R _33868_ (.SN(_17815_),
    .A(_16958_),
    .B(_16959_),
    .CI(_16960_),
    .CON(_17841_));
 FAx1_ASAP7_75t_R _33869_ (.SN(_16966_),
    .A(_16963_),
    .B(_16964_),
    .CI(_16965_),
    .CON(_17024_));
 FAx1_ASAP7_75t_R _33870_ (.SN(_17817_),
    .A(_16962_),
    .B(_16906_),
    .CI(_16966_),
    .CON(_17843_));
 FAx1_ASAP7_75t_R _33871_ (.SN(_17818_),
    .A(_16969_),
    .B(_16970_),
    .CI(_16971_),
    .CON(_17845_));
 FAx1_ASAP7_75t_R _33872_ (.SN(_17820_),
    .A(_16974_),
    .B(_16973_),
    .CI(_16917_),
    .CON(_17852_));
 FAx1_ASAP7_75t_R _33873_ (.SN(_17821_),
    .A(_16968_),
    .B(_16977_),
    .CI(_16976_),
    .CON(_17848_));
 FAx1_ASAP7_75t_R _33874_ (.SN(_17822_),
    .A(_16980_),
    .B(_16981_),
    .CI(_16982_),
    .CON(_17850_));
 FAx1_ASAP7_75t_R _33875_ (.SN(_16988_),
    .A(_16985_),
    .B(_16986_),
    .CI(_16987_),
    .CON(_17048_));
 FAx1_ASAP7_75t_R _33876_ (.SN(_17825_),
    .A(_16984_),
    .B(_16926_),
    .CI(_16988_),
    .CON(_17854_));
 FAx1_ASAP7_75t_R _33877_ (.SN(_17827_),
    .A(_16920_),
    .B(_16990_),
    .CI(_16932_),
    .CON(_17050_));
 FAx1_ASAP7_75t_R _33878_ (.SN(_17828_),
    .A(_16979_),
    .B(_16992_),
    .CI(_16991_),
    .CON(_17857_));
 FAx1_ASAP7_75t_R _33879_ (.SN(_17830_),
    .A(_16995_),
    .B(_16996_),
    .CI(_16997_),
    .CON(_17858_));
 FAx1_ASAP7_75t_R _33880_ (.SN(_17832_),
    .A(_17000_),
    .B(_16999_),
    .CI(_16943_),
    .CON(_17860_));
 FAx1_ASAP7_75t_R _33881_ (.SN(_17835_),
    .A(_16934_),
    .B(_17001_),
    .CI(_17002_),
    .CON(_17863_));
 FAx1_ASAP7_75t_R _33882_ (.SN(_17836_),
    .A(_16994_),
    .B(_16938_),
    .CI(_17004_),
    .CON(_17862_));
 FAx1_ASAP7_75t_R _33883_ (.SN(_17838_),
    .A(_17006_),
    .B(_16953_),
    .CI(_17007_),
    .CON(_17057_));
 FAx1_ASAP7_75t_R _33884_ (.SN(_17840_),
    .A(_17008_),
    .B(_17009_),
    .CI(_17010_),
    .CON(_17865_));
 FAx1_ASAP7_75t_R _33885_ (.SN(_17016_),
    .A(_17013_),
    .B(_17014_),
    .CI(_17015_),
    .CON(_17075_));
 FAx1_ASAP7_75t_R _33886_ (.SN(_17842_),
    .A(_17012_),
    .B(_16961_),
    .CI(_17016_),
    .CON(_17867_));
 FAx1_ASAP7_75t_R _33887_ (.SN(_17844_),
    .A(_17019_),
    .B(_17020_),
    .CI(_17021_),
    .CON(_17869_));
 FAx1_ASAP7_75t_R _33888_ (.SN(_17846_),
    .A(_17024_),
    .B(_17023_),
    .CI(_16972_),
    .CON(_17876_));
 FAx1_ASAP7_75t_R _33889_ (.SN(_17847_),
    .A(_17018_),
    .B(_16967_),
    .CI(_17026_),
    .CON(_17872_));
 FAx1_ASAP7_75t_R _33890_ (.SN(_17849_),
    .A(_17029_),
    .B(_17030_),
    .CI(_17031_),
    .CON(_17874_));
 FAx1_ASAP7_75t_R _33891_ (.SN(_17851_),
    .A(_17034_),
    .B(_17035_),
    .CI(_17036_),
    .CON(_17882_));
 FAx1_ASAP7_75t_R _33892_ (.SN(_17853_),
    .A(_17033_),
    .B(_16983_),
    .CI(_17038_),
    .CON(_17878_));
 FAx1_ASAP7_75t_R _33893_ (.SN(_17855_),
    .A(_16975_),
    .B(_17040_),
    .CI(_16989_),
    .CON(_17096_));
 FAx1_ASAP7_75t_R _33894_ (.SN(_17856_),
    .A(_17028_),
    .B(_16978_),
    .CI(_17041_),
    .CON(_17881_));
 FAx1_ASAP7_75t_R _33895_ (.SN(_17049_),
    .A(_16948_),
    .B(_17044_),
    .CI(_17045_),
    .CON(_17095_));
 FAx1_ASAP7_75t_R _33896_ (.SN(_17859_),
    .A(_17048_),
    .B(_17049_),
    .CI(_16998_),
    .CON(_17884_));
 FAx1_ASAP7_75t_R _33897_ (.SN(_17053_),
    .A(_17050_),
    .B(_17051_),
    .CI(_17052_),
    .CON(_17102_));
 FAx1_ASAP7_75t_R _33898_ (.SN(_17861_),
    .A(_17043_),
    .B(_16993_),
    .CI(_17053_),
    .CON(_17886_));
 FAx1_ASAP7_75t_R _33899_ (.SN(_17056_),
    .A(_17055_),
    .B(_17005_),
    .CI(_17003_),
    .CON(_17888_));
 FAx1_ASAP7_75t_R _33900_ (.SN(_02243_),
    .A(_17056_),
    .B(_17057_),
    .CI(_17058_),
    .CON(_02242_));
 FAx1_ASAP7_75t_R _33901_ (.SN(_17864_),
    .A(_17059_),
    .B(_17060_),
    .CI(_17061_),
    .CON(_17890_));
 FAx1_ASAP7_75t_R _33902_ (.SN(_17067_),
    .A(_17064_),
    .B(_17065_),
    .CI(_17066_),
    .CON(_17119_));
 FAx1_ASAP7_75t_R _33903_ (.SN(_17866_),
    .A(_17063_),
    .B(_17011_),
    .CI(_17067_),
    .CON(_17892_));
 FAx1_ASAP7_75t_R _33904_ (.SN(_17868_),
    .A(_17070_),
    .B(_17071_),
    .CI(_17072_),
    .CON(_17894_));
 FAx1_ASAP7_75t_R _33905_ (.SN(_17870_),
    .A(_17075_),
    .B(_17074_),
    .CI(_17022_),
    .CON(_17901_));
 FAx1_ASAP7_75t_R _33906_ (.SN(_17871_),
    .A(_17069_),
    .B(_17017_),
    .CI(_17077_),
    .CON(_17897_));
 FAx1_ASAP7_75t_R _33907_ (.SN(_17873_),
    .A(_17080_),
    .B(_17081_),
    .CI(_17082_),
    .CON(_17899_));
 FAx1_ASAP7_75t_R _33908_ (.SN(_17875_),
    .A(_17085_),
    .B(_17086_),
    .CI(_17087_),
    .CON(_17907_));
 FAx1_ASAP7_75t_R _33909_ (.SN(_17877_),
    .A(_17084_),
    .B(_17032_),
    .CI(_17089_),
    .CON(_17903_));
 FAx1_ASAP7_75t_R _33910_ (.SN(_17879_),
    .A(_17025_),
    .B(_17091_),
    .CI(_17039_),
    .CON(_17137_));
 FAx1_ASAP7_75t_R _33911_ (.SN(_17880_),
    .A(_17079_),
    .B(_17027_),
    .CI(_17092_),
    .CON(_17906_));
 FAx1_ASAP7_75t_R _33912_ (.SN(_17883_),
    .A(_17049_),
    .B(_17037_),
    .CI(_17095_),
    .CON(_17909_));
 FAx1_ASAP7_75t_R _33913_ (.SN(_17099_),
    .A(_17096_),
    .B(_17097_),
    .CI(_17098_),
    .CON(_17143_));
 FAx1_ASAP7_75t_R _33914_ (.SN(_17885_),
    .A(_17094_),
    .B(_17042_),
    .CI(_17099_),
    .CON(_17911_));
 FAx1_ASAP7_75t_R _33915_ (.SN(_17887_),
    .A(_17101_),
    .B(_17054_),
    .CI(_17102_),
    .CON(_17145_));
 FAx1_ASAP7_75t_R _33916_ (.SN(_17889_),
    .A(_17103_),
    .B(_17104_),
    .CI(_17105_),
    .CON(_17913_));
 FAx1_ASAP7_75t_R _33917_ (.SN(_17111_),
    .A(_17108_),
    .B(_17109_),
    .CI(_17110_),
    .CON(_17164_));
 FAx1_ASAP7_75t_R _33918_ (.SN(_17891_),
    .A(_17107_),
    .B(_17062_),
    .CI(_17111_),
    .CON(_17916_));
 FAx1_ASAP7_75t_R _33919_ (.SN(_17893_),
    .A(_17114_),
    .B(_17115_),
    .CI(_17116_),
    .CON(_17918_));
 FAx1_ASAP7_75t_R _33920_ (.SN(_17895_),
    .A(_17119_),
    .B(_17118_),
    .CI(_17073_),
    .CON(_17924_));
 FAx1_ASAP7_75t_R _33921_ (.SN(_17896_),
    .A(_17113_),
    .B(_17068_),
    .CI(_17121_),
    .CON(_17921_));
 FAx1_ASAP7_75t_R _33922_ (.SN(_17898_),
    .A(_17124_),
    .B(_17125_),
    .CI(_17126_),
    .CON(_17923_));
 FAx1_ASAP7_75t_R _33923_ (.SN(_17900_),
    .A(_17087_),
    .B(_17129_),
    .CI(_17130_),
    .CON(_17185_));
 FAx1_ASAP7_75t_R _33924_ (.SN(_17902_),
    .A(_17128_),
    .B(_17083_),
    .CI(_17131_),
    .CON(_17926_));
 FAx1_ASAP7_75t_R _33925_ (.SN(_17904_),
    .A(_17076_),
    .B(_17133_),
    .CI(_17090_),
    .CON(_17188_));
 FAx1_ASAP7_75t_R _33926_ (.SN(_17905_),
    .A(_17123_),
    .B(_17078_),
    .CI(_17134_),
    .CON(_17929_));
 FAx1_ASAP7_75t_R _33927_ (.SN(_17908_),
    .A(_17049_),
    .B(_17095_),
    .CI(_17088_),
    .CON(_17930_));
 FAx1_ASAP7_75t_R _33928_ (.SN(_17140_),
    .A(_17137_),
    .B(_17138_),
    .CI(_17139_),
    .CON(_17194_));
 FAx1_ASAP7_75t_R _33929_ (.SN(_17910_),
    .A(_17136_),
    .B(_17093_),
    .CI(_17140_),
    .CON(_17932_));
 FAx1_ASAP7_75t_R _33930_ (.SN(_17144_),
    .A(_17142_),
    .B(_17100_),
    .CI(_17143_),
    .CON(_17934_));
 FAx1_ASAP7_75t_R _33931_ (.SN(_02245_),
    .A(_17144_),
    .B(_17145_),
    .CI(_17146_),
    .CON(_02244_));
 FAx1_ASAP7_75t_R _33932_ (.SN(_17912_),
    .A(_17147_),
    .B(_17148_),
    .CI(_17149_),
    .CON(_17936_));
 FAx1_ASAP7_75t_R _33933_ (.SN(_17914_),
    .A(_17152_),
    .B(_17153_),
    .CI(_17154_),
    .CON(_17940_));
 FAx1_ASAP7_75t_R _33934_ (.SN(_17915_),
    .A(_17151_),
    .B(_17106_),
    .CI(_17156_),
    .CON(_17939_));
 FAx1_ASAP7_75t_R _33935_ (.SN(_17917_),
    .A(_17159_),
    .B(_17160_),
    .CI(_17161_),
    .CON(_17942_));
 FAx1_ASAP7_75t_R _33936_ (.SN(_17919_),
    .A(_17164_),
    .B(_17163_),
    .CI(_17117_),
    .CON(_17948_));
 FAx1_ASAP7_75t_R _33937_ (.SN(_17920_),
    .A(_17158_),
    .B(_17112_),
    .CI(_17166_),
    .CON(_17945_));
 FAx1_ASAP7_75t_R _33938_ (.SN(_17922_),
    .A(_17169_),
    .B(_17170_),
    .CI(_17171_),
    .CON(_17947_));
 FAx1_ASAP7_75t_R _33939_ (.SN(_17179_),
    .A(_17174_),
    .B(_17175_),
    .CI(_17176_),
    .CON(_17227_));
 FAx1_ASAP7_75t_R _33940_ (.SN(_17925_),
    .A(_17173_),
    .B(_17127_),
    .CI(_17179_),
    .CON(_17950_));
 FAx1_ASAP7_75t_R _33941_ (.SN(_17927_),
    .A(_17120_),
    .B(_17181_),
    .CI(_17132_),
    .CON(_17228_));
 FAx1_ASAP7_75t_R _33942_ (.SN(_17928_),
    .A(_17168_),
    .B(_17122_),
    .CI(_17182_),
    .CON(_17953_));
 FAx1_ASAP7_75t_R _33943_ (.SN(_00042_),
    .A(_17047_),
    .B(_17046_),
    .CI(_17185_),
    .CON(_00047_));
 FAx1_ASAP7_75t_R _33944_ (.SN(_17191_),
    .A(_17188_),
    .B(_17189_),
    .CI(_17190_),
    .CON(_17234_));
 FAx1_ASAP7_75t_R _33945_ (.SN(_17931_),
    .A(_17184_),
    .B(_17135_),
    .CI(_17191_),
    .CON(_17955_));
 FAx1_ASAP7_75t_R _33946_ (.SN(_17933_),
    .A(_17193_),
    .B(_17141_),
    .CI(_17194_),
    .CON(_17236_));
 FAx1_ASAP7_75t_R _33947_ (.SN(_17935_),
    .A(_17195_),
    .B(_17196_),
    .CI(_17197_),
    .CON(_17957_));
 FAx1_ASAP7_75t_R _33948_ (.SN(_17937_),
    .A(_17200_),
    .B(_17201_),
    .CI(_17202_),
    .CON(_17961_));
 FAx1_ASAP7_75t_R _33949_ (.SN(_17938_),
    .A(_17199_),
    .B(_17150_),
    .CI(_17204_),
    .CON(_17960_));
 FAx1_ASAP7_75t_R _33950_ (.SN(_17941_),
    .A(_17207_),
    .B(_17208_),
    .CI(_17209_),
    .CON(_17963_));
 FAx1_ASAP7_75t_R _33951_ (.SN(_17943_),
    .A(_17155_),
    .B(_17211_),
    .CI(_17162_),
    .CON(_17967_));
 FAx1_ASAP7_75t_R _33952_ (.SN(_17944_),
    .A(_17206_),
    .B(_17157_),
    .CI(_17213_),
    .CON(_17966_));
 FAx1_ASAP7_75t_R _33953_ (.SN(_17946_),
    .A(_17216_),
    .B(_17217_),
    .CI(_17218_),
    .CON(_17262_));
 FAx1_ASAP7_75t_R _33954_ (.SN(_17949_),
    .A(_17179_),
    .B(_17219_),
    .CI(_17172_),
    .CON(_17968_));
 FAx1_ASAP7_75t_R _33955_ (.SN(_17951_),
    .A(_17165_),
    .B(_17221_),
    .CI(_17180_),
    .CON(_17267_));
 FAx1_ASAP7_75t_R _33956_ (.SN(_17952_),
    .A(_17215_),
    .B(_17167_),
    .CI(_17222_),
    .CON(_17971_));
 FAx1_ASAP7_75t_R _33957_ (.SN(_00046_),
    .A(_17047_),
    .B(_17046_),
    .CI(_17177_),
    .CON(_00050_));
 FAx1_ASAP7_75t_R _33958_ (.SN(_17231_),
    .A(_17228_),
    .B(_17229_),
    .CI(_17230_),
    .CON(_17273_));
 FAx1_ASAP7_75t_R _33959_ (.SN(_17954_),
    .A(_17224_),
    .B(_17183_),
    .CI(_17231_),
    .CON(_17973_));
 FAx1_ASAP7_75t_R _33960_ (.SN(_17235_),
    .A(_17233_),
    .B(_17192_),
    .CI(_17234_),
    .CON(_17975_));
 FAx1_ASAP7_75t_R _33961_ (.SN(_02247_),
    .A(_17235_),
    .B(_17236_),
    .CI(_17237_),
    .CON(_02246_));
 FAx1_ASAP7_75t_R _33962_ (.SN(_17956_),
    .A(_17238_),
    .B(_17239_),
    .CI(_17240_),
    .CON(_17977_));
 FAx1_ASAP7_75t_R _33963_ (.SN(_17958_),
    .A(_17243_),
    .B(_17244_),
    .CI(_17245_),
    .CON(_17981_));
 FAx1_ASAP7_75t_R _33964_ (.SN(_17959_),
    .A(_17242_),
    .B(_17198_),
    .CI(_17247_),
    .CON(_17980_));
 FAx1_ASAP7_75t_R _33965_ (.SN(_17962_),
    .A(_17250_),
    .B(_17251_),
    .CI(_17252_),
    .CON(_17983_));
 FAx1_ASAP7_75t_R _33966_ (.SN(_17964_),
    .A(_17203_),
    .B(_17254_),
    .CI(_17210_),
    .CON(_17987_));
 FAx1_ASAP7_75t_R _33967_ (.SN(_17965_),
    .A(_17249_),
    .B(_17205_),
    .CI(_17256_),
    .CON(_17986_));
 FAx1_ASAP7_75t_R _33968_ (.SN(_17261_),
    .A(_17218_),
    .B(_17259_),
    .CI(_17260_),
    .CON(_17300_));
 FAx1_ASAP7_75t_R _33969_ (.SN(_17263_),
    .A(_17178_),
    .B(_17261_),
    .CI(_17262_),
    .CON(_17303_));
 FAx1_ASAP7_75t_R _33970_ (.SN(_17969_),
    .A(_17212_),
    .B(_17263_),
    .CI(_17220_),
    .CON(_17307_));
 FAx1_ASAP7_75t_R _33971_ (.SN(_17970_),
    .A(_17258_),
    .B(_17214_),
    .CI(_17264_),
    .CON(_17990_));
 FAx1_ASAP7_75t_R _33972_ (.SN(_17270_),
    .A(_17267_),
    .B(_17268_),
    .CI(_17269_),
    .CON(_17312_));
 FAx1_ASAP7_75t_R _33973_ (.SN(_17972_),
    .A(_17266_),
    .B(_17223_),
    .CI(_17270_),
    .CON(_17992_));
 FAx1_ASAP7_75t_R _33974_ (.SN(_17974_),
    .A(_17272_),
    .B(_17232_),
    .CI(_17273_),
    .CON(_17314_));
 FAx1_ASAP7_75t_R _33975_ (.SN(_17976_),
    .A(_17274_),
    .B(_17275_),
    .CI(_17276_),
    .CON(_17994_));
 FAx1_ASAP7_75t_R _33976_ (.SN(_17978_),
    .A(_17279_),
    .B(_17280_),
    .CI(_17281_),
    .CON(_17998_));
 FAx1_ASAP7_75t_R _33977_ (.SN(_17979_),
    .A(_17278_),
    .B(_17241_),
    .CI(_17283_),
    .CON(_17997_));
 FAx1_ASAP7_75t_R _33978_ (.SN(_17982_),
    .A(_17286_),
    .B(_17287_),
    .CI(_17288_),
    .CON(_18000_));
 FAx1_ASAP7_75t_R _33979_ (.SN(_17984_),
    .A(_17246_),
    .B(_17290_),
    .CI(_17253_),
    .CON(_18004_));
 FAx1_ASAP7_75t_R _33980_ (.SN(_17985_),
    .A(_17285_),
    .B(_17248_),
    .CI(_17292_),
    .CON(_18003_));
 FAx1_ASAP7_75t_R _33981_ (.SN(_17301_),
    .A(_17295_),
    .B(_17296_),
    .CI(_17297_),
    .CON(_17339_));
 FAx1_ASAP7_75t_R _33982_ (.SN(_17302_),
    .A(_17178_),
    .B(_17299_),
    .CI(_17300_),
    .CON(_17341_));
 FAx1_ASAP7_75t_R _33983_ (.SN(_17988_),
    .A(_17255_),
    .B(_17302_),
    .CI(_17303_),
    .CON(_17345_));
 FAx1_ASAP7_75t_R _33984_ (.SN(_17989_),
    .A(_17294_),
    .B(_17257_),
    .CI(_17304_),
    .CON(_18007_));
 FAx1_ASAP7_75t_R _33985_ (.SN(_17309_),
    .A(_17268_),
    .B(_17307_),
    .CI(_17308_),
    .CON(_17349_));
 FAx1_ASAP7_75t_R _33986_ (.SN(_17991_),
    .A(_17306_),
    .B(_17265_),
    .CI(_17309_),
    .CON(_18009_));
 FAx1_ASAP7_75t_R _33987_ (.SN(_17313_),
    .A(_17311_),
    .B(_17271_),
    .CI(_17312_),
    .CON(_18011_));
 FAx1_ASAP7_75t_R _33988_ (.SN(_02249_),
    .A(_17313_),
    .B(_17314_),
    .CI(_17315_),
    .CON(_02248_));
 FAx1_ASAP7_75t_R _33989_ (.SN(_17993_),
    .A(_17316_),
    .B(_17317_),
    .CI(_17318_),
    .CON(_18013_));
 FAx1_ASAP7_75t_R _33990_ (.SN(_17995_),
    .A(_17321_),
    .B(_17322_),
    .CI(_17323_),
    .CON(_18017_));
 FAx1_ASAP7_75t_R _33991_ (.SN(_17996_),
    .A(_17320_),
    .B(_17277_),
    .CI(_17325_),
    .CON(_18016_));
 FAx1_ASAP7_75t_R _33992_ (.SN(_17999_),
    .A(_17328_),
    .B(_17329_),
    .CI(_17330_),
    .CON(_18019_));
 FAx1_ASAP7_75t_R _33993_ (.SN(_18001_),
    .A(_17282_),
    .B(_17332_),
    .CI(_17289_),
    .CON(_18023_));
 FAx1_ASAP7_75t_R _33994_ (.SN(_18002_),
    .A(_17327_),
    .B(_17284_),
    .CI(_17334_),
    .CON(_18022_));
 FAx1_ASAP7_75t_R _33995_ (.SN(_17340_),
    .A(_17178_),
    .B(_17299_),
    .CI(_17298_),
    .CON(_17370_));
 FAx1_ASAP7_75t_R _33996_ (.SN(_18005_),
    .A(_17291_),
    .B(_17340_),
    .CI(_17341_),
    .CON(_17374_));
 FAx1_ASAP7_75t_R _33997_ (.SN(_18006_),
    .A(_17336_),
    .B(_17293_),
    .CI(_17342_),
    .CON(_18026_));
 FAx1_ASAP7_75t_R _33998_ (.SN(_17346_),
    .A(_17268_),
    .B(_17308_),
    .CI(_17345_),
    .CON(_17378_));
 FAx1_ASAP7_75t_R _33999_ (.SN(_18008_),
    .A(_17344_),
    .B(_17305_),
    .CI(_17346_),
    .CON(_18028_));
 FAx1_ASAP7_75t_R _34000_ (.SN(_18010_),
    .A(_17348_),
    .B(_17310_),
    .CI(_17349_),
    .CON(_17380_));
 FAx1_ASAP7_75t_R _34001_ (.SN(_18012_),
    .A(_17350_),
    .B(_17351_),
    .CI(_17352_),
    .CON(_18030_));
 FAx1_ASAP7_75t_R _34002_ (.SN(_18014_),
    .A(_17355_),
    .B(_17356_),
    .CI(_17357_),
    .CON(_18034_));
 FAx1_ASAP7_75t_R _34003_ (.SN(_18015_),
    .A(_17354_),
    .B(_17319_),
    .CI(_17359_),
    .CON(_18033_));
 FAx1_ASAP7_75t_R _34004_ (.SN(_18018_),
    .A(_17330_),
    .B(_17362_),
    .CI(_17363_),
    .CON(_18035_));
 FAx1_ASAP7_75t_R _34005_ (.SN(_18020_),
    .A(_17324_),
    .B(_17365_),
    .CI(_17331_),
    .CON(_18039_));
 FAx1_ASAP7_75t_R _34006_ (.SN(_18021_),
    .A(_17361_),
    .B(_17326_),
    .CI(_17367_),
    .CON(_18038_));
 FAx1_ASAP7_75t_R _34007_ (.SN(_18024_),
    .A(_17340_),
    .B(_17333_),
    .CI(_17370_),
    .CON(_17407_));
 FAx1_ASAP7_75t_R _34008_ (.SN(_18025_),
    .A(_17369_),
    .B(_17335_),
    .CI(_17371_),
    .CON(_18042_));
 FAx1_ASAP7_75t_R _34009_ (.SN(_17375_),
    .A(_17268_),
    .B(_17308_),
    .CI(_17374_),
    .CON(_17411_));
 FAx1_ASAP7_75t_R _34010_ (.SN(_18027_),
    .A(_17373_),
    .B(_17343_),
    .CI(_17375_),
    .CON(_18044_));
 FAx1_ASAP7_75t_R _34011_ (.SN(_17379_),
    .A(_17377_),
    .B(_17347_),
    .CI(_17378_),
    .CON(_18046_));
 FAx1_ASAP7_75t_R _34012_ (.SN(_02251_),
    .A(_17379_),
    .B(_17380_),
    .CI(_17381_),
    .CON(_02250_));
 FAx1_ASAP7_75t_R _34013_ (.SN(_18029_),
    .A(_17382_),
    .B(_17383_),
    .CI(_17384_),
    .CON(_18048_));
 FAx1_ASAP7_75t_R _34014_ (.SN(_18031_),
    .A(_17387_),
    .B(_17388_),
    .CI(_17389_),
    .CON(_18052_));
 FAx1_ASAP7_75t_R _34015_ (.SN(_18032_),
    .A(_17386_),
    .B(_17353_),
    .CI(_17391_),
    .CON(_18051_));
 FAx1_ASAP7_75t_R _34016_ (.SN(_17399_),
    .A(_17394_),
    .B(_17395_),
    .CI(_17396_),
    .CON(_17424_));
 FAx1_ASAP7_75t_R _34017_ (.SN(_18036_),
    .A(_17358_),
    .B(_17399_),
    .CI(_17364_),
    .CON(_18056_));
 FAx1_ASAP7_75t_R _34018_ (.SN(_18037_),
    .A(_17393_),
    .B(_17360_),
    .CI(_17401_),
    .CON(_18055_));
 FAx1_ASAP7_75t_R _34019_ (.SN(_18040_),
    .A(net278),
    .B(_17370_),
    .CI(_17366_),
    .CON(_17432_));
 FAx1_ASAP7_75t_R _34020_ (.SN(_18041_),
    .A(_17403_),
    .B(_17368_),
    .CI(_17404_),
    .CON(_18059_));
 FAx1_ASAP7_75t_R _34021_ (.SN(_17408_),
    .A(_17268_),
    .B(_17308_),
    .CI(_17407_),
    .CON(_17436_));
 FAx1_ASAP7_75t_R _34022_ (.SN(_18043_),
    .A(_17406_),
    .B(_17372_),
    .CI(_17408_),
    .CON(_18061_));
 FAx1_ASAP7_75t_R _34023_ (.SN(_18045_),
    .A(_17410_),
    .B(_17376_),
    .CI(_17411_),
    .CON(_17438_));
 FAx1_ASAP7_75t_R _34024_ (.SN(_18047_),
    .A(_17412_),
    .B(_17413_),
    .CI(_17414_),
    .CON(_18063_));
 FAx1_ASAP7_75t_R _34025_ (.SN(_18049_),
    .A(_17417_),
    .B(_17418_),
    .CI(_17419_),
    .CON(_18067_));
 FAx1_ASAP7_75t_R _34026_ (.SN(_18050_),
    .A(_17416_),
    .B(_17385_),
    .CI(_17421_),
    .CON(_18066_));
 FAx1_ASAP7_75t_R _34027_ (.SN(_18053_),
    .A(_17399_),
    .B(_17390_),
    .CI(_17424_),
    .CON(_18071_));
 FAx1_ASAP7_75t_R _34028_ (.SN(_18054_),
    .A(_17423_),
    .B(_17392_),
    .CI(_17426_),
    .CON(_18070_));
 FAx1_ASAP7_75t_R _34029_ (.SN(_18057_),
    .A(net278),
    .B(_17370_),
    .CI(_17400_),
    .CON(_17457_));
 FAx1_ASAP7_75t_R _34030_ (.SN(_18058_),
    .A(_17428_),
    .B(_17402_),
    .CI(_17429_),
    .CON(_18074_));
 FAx1_ASAP7_75t_R _34031_ (.SN(_17433_),
    .A(_17268_),
    .B(_17308_),
    .CI(_17432_),
    .CON(_17461_));
 FAx1_ASAP7_75t_R _34032_ (.SN(_18060_),
    .A(_17431_),
    .B(_17405_),
    .CI(_17433_),
    .CON(_18076_));
 FAx1_ASAP7_75t_R _34033_ (.SN(_17437_),
    .A(_17435_),
    .B(_17409_),
    .CI(_17436_),
    .CON(_18078_));
 FAx1_ASAP7_75t_R _34034_ (.SN(_02253_),
    .A(_17437_),
    .B(_17438_),
    .CI(_17439_),
    .CON(_02252_));
 FAx1_ASAP7_75t_R _34035_ (.SN(_18062_),
    .A(_17440_),
    .B(_17441_),
    .CI(_17442_),
    .CON(_17475_));
 FAx1_ASAP7_75t_R _34036_ (.SN(_18064_),
    .A(_17419_),
    .B(_17445_),
    .CI(_17446_),
    .CON(_17476_));
 FAx1_ASAP7_75t_R _34037_ (.SN(_18065_),
    .A(_17444_),
    .B(_17415_),
    .CI(_17447_),
    .CON(_18080_));
 FAx1_ASAP7_75t_R _34038_ (.SN(_18068_),
    .A(_17399_),
    .B(_17424_),
    .CI(_17420_),
    .CON(_18083_));
 FAx1_ASAP7_75t_R _34039_ (.SN(_18069_),
    .A(_17449_),
    .B(_17422_),
    .CI(_17451_),
    .CON(_18082_));
 FAx1_ASAP7_75t_R _34040_ (.SN(_18072_),
    .A(net278),
    .B(_17370_),
    .CI(_17425_),
    .CON(_17484_));
 FAx1_ASAP7_75t_R _34041_ (.SN(_18073_),
    .A(_17453_),
    .B(_17427_),
    .CI(_17454_),
    .CON(_18086_));
 FAx1_ASAP7_75t_R _34042_ (.SN(_17458_),
    .A(_17268_),
    .B(_17308_),
    .CI(_17457_),
    .CON(_17488_));
 FAx1_ASAP7_75t_R _34043_ (.SN(_18075_),
    .A(_17456_),
    .B(_17430_),
    .CI(_17458_),
    .CON(_18088_));
 FAx1_ASAP7_75t_R _34044_ (.SN(_18077_),
    .A(_17460_),
    .B(_17434_),
    .CI(_17461_),
    .CON(_17490_));
 FAx1_ASAP7_75t_R _34045_ (.SN(_17474_),
    .A(_17462_),
    .B(_17463_),
    .CI(_17464_),
    .CON(_17496_));
 FAx1_ASAP7_75t_R _34046_ (.SN(_17471_),
    .A(_17466_),
    .B(_17467_),
    .CI(_17468_),
    .CON(_17500_));
 FAx1_ASAP7_75t_R _34047_ (.SN(_18079_),
    .A(_17465_),
    .B(_17443_),
    .CI(_17471_),
    .CON(_17505_));
 FAx1_ASAP7_75t_R _34048_ (.SN(_17478_),
    .A(_17398_),
    .B(_17397_),
    .CI(_17476_),
    .CON(_17507_));
 FAx1_ASAP7_75t_R _34049_ (.SN(_18081_),
    .A(_17473_),
    .B(_17448_),
    .CI(_17478_),
    .CON(_18090_));
 FAx1_ASAP7_75t_R _34050_ (.SN(_18084_),
    .A(net278),
    .B(_17370_),
    .CI(_17450_),
    .CON(_17511_));
 FAx1_ASAP7_75t_R _34051_ (.SN(_18085_),
    .A(_17480_),
    .B(_17452_),
    .CI(_17481_),
    .CON(_18092_));
 FAx1_ASAP7_75t_R _34052_ (.SN(_17485_),
    .A(_17268_),
    .B(_17308_),
    .CI(_17484_),
    .CON(_17515_));
 FAx1_ASAP7_75t_R _34053_ (.SN(_18087_),
    .A(_17483_),
    .B(_17455_),
    .CI(_17485_),
    .CON(_18094_));
 FAx1_ASAP7_75t_R _34054_ (.SN(_17489_),
    .A(_17487_),
    .B(_17459_),
    .CI(_17488_),
    .CON(_18096_));
 FAx1_ASAP7_75t_R _34055_ (.SN(_02255_),
    .A(_17489_),
    .B(_17490_),
    .CI(_17491_),
    .CON(_02254_));
 FAx1_ASAP7_75t_R _34056_ (.SN(_17495_),
    .A(_17492_),
    .B(_17493_),
    .CI(_17494_),
    .CON(_17520_));
 FAx1_ASAP7_75t_R _34057_ (.SN(_17501_),
    .A(_17470_),
    .B(_17495_),
    .CI(_17496_),
    .CON(_17523_));
 FAx1_ASAP7_75t_R _34058_ (.SN(_17502_),
    .A(_17398_),
    .B(_17397_),
    .CI(_17469_),
    .CON(_17524_));
 FAx1_ASAP7_75t_R _34059_ (.SN(_18089_),
    .A(_17501_),
    .B(_17472_),
    .CI(_17502_),
    .CON(_18097_));
 FAx1_ASAP7_75t_R _34060_ (.SN(_17508_),
    .A(_17338_),
    .B(_17337_),
    .CI(_17477_),
    .CON(_00066_));
 FAx1_ASAP7_75t_R _34061_ (.SN(_18091_),
    .A(_17504_),
    .B(_17479_),
    .CI(_17508_),
    .CON(_18099_));
 FAx1_ASAP7_75t_R _34062_ (.SN(_17512_),
    .A(_17268_),
    .B(_17308_),
    .CI(_17511_),
    .CON(_17530_));
 FAx1_ASAP7_75t_R _34063_ (.SN(_18093_),
    .A(_17510_),
    .B(_17482_),
    .CI(_17512_),
    .CON(_18101_));
 FAx1_ASAP7_75t_R _34064_ (.SN(_18095_),
    .A(_17514_),
    .B(_17486_),
    .CI(_17515_),
    .CON(_18103_));
 FAx1_ASAP7_75t_R _34065_ (.SN(_17519_),
    .A(_17494_),
    .B(_17517_),
    .CI(_17518_),
    .CON(_02256_));
 FAx1_ASAP7_75t_R _34066_ (.SN(_17522_),
    .A(_17470_),
    .B(_17519_),
    .CI(_17520_),
    .CON(_00068_));
 FAx1_ASAP7_75t_R _34067_ (.SN(_17525_),
    .A(_17499_),
    .B(_17521_),
    .CI(_17497_),
    .CON(_00069_));
 FAx1_ASAP7_75t_R _34068_ (.SN(_17526_),
    .A(_17338_),
    .B(_17337_),
    .CI(_17498_),
    .CON(_00070_));
 FAx1_ASAP7_75t_R _34069_ (.SN(_18098_),
    .A(_17525_),
    .B(_17503_),
    .CI(_17526_),
    .CON(_02257_));
 FAx1_ASAP7_75t_R _34070_ (.SN(_17528_),
    .A(_17268_),
    .B(_17308_),
    .CI(_17506_),
    .CON(_00071_));
 FAx1_ASAP7_75t_R _34071_ (.SN(_18100_),
    .A(_17527_),
    .B(_17509_),
    .CI(_17528_),
    .CON(_02258_));
 FAx1_ASAP7_75t_R _34072_ (.SN(_18102_),
    .A(_17529_),
    .B(_17513_),
    .CI(_17530_),
    .CON(_02259_));
 FAx1_ASAP7_75t_R _34073_ (.SN(_02261_),
    .A(_17531_),
    .B(_17516_),
    .CI(_17532_),
    .CON(_02260_));
 FAx1_ASAP7_75t_R _34074_ (.SN(_00241_),
    .A(_17533_),
    .B(_17534_),
    .CI(\cs_registers_i.pc_if_i[2] ),
    .CON(_00242_));
 HAxp5_ASAP7_75t_R _34075_ (.A(_17537_),
    .B(_17538_),
    .CON(_00664_),
    .SN(_00292_));
 HAxp5_ASAP7_75t_R _34076_ (.A(_17540_),
    .B(_17541_),
    .CON(_00667_),
    .SN(_02262_));
 HAxp5_ASAP7_75t_R _34077_ (.A(_17542_),
    .B(_17543_),
    .CON(_00669_),
    .SN(_00666_));
 HAxp5_ASAP7_75t_R _34078_ (.A(_17544_),
    .B(_17545_),
    .CON(_02263_),
    .SN(_02264_));
 HAxp5_ASAP7_75t_R _34079_ (.A(_17546_),
    .B(_17547_),
    .CON(_00673_),
    .SN(_00671_));
 HAxp5_ASAP7_75t_R _34080_ (.A(_17548_),
    .B(_17549_),
    .CON(_02265_),
    .SN(_02266_));
 HAxp5_ASAP7_75t_R _34081_ (.A(_16510_),
    .B(_16511_),
    .CON(_00678_),
    .SN(_00675_));
 HAxp5_ASAP7_75t_R _34082_ (.A(_17550_),
    .B(_17551_),
    .CON(_02267_),
    .SN(_02268_));
 HAxp5_ASAP7_75t_R _34083_ (.A(_17552_),
    .B(_17553_),
    .CON(_00683_),
    .SN(_00681_));
 HAxp5_ASAP7_75t_R _34084_ (.A(_17554_),
    .B(_17555_),
    .CON(_02269_),
    .SN(_02270_));
 HAxp5_ASAP7_75t_R _34085_ (.A(_17556_),
    .B(_17557_),
    .CON(_00687_),
    .SN(_00685_));
 HAxp5_ASAP7_75t_R _34086_ (.A(_17558_),
    .B(_17559_),
    .CON(_02271_),
    .SN(_02272_));
 HAxp5_ASAP7_75t_R _34087_ (.A(_17560_),
    .B(_17561_),
    .CON(_00752_),
    .SN(_00719_));
 HAxp5_ASAP7_75t_R _34088_ (.A(_17562_),
    .B(_17563_),
    .CON(_02273_),
    .SN(_00751_));
 HAxp5_ASAP7_75t_R _34089_ (.A(_16522_),
    .B(_16524_),
    .CON(_00817_),
    .SN(_00784_));
 HAxp5_ASAP7_75t_R _34090_ (.A(_17564_),
    .B(_17565_),
    .CON(_02274_),
    .SN(_02275_));
 HAxp5_ASAP7_75t_R _34091_ (.A(_17566_),
    .B(_17567_),
    .CON(_00883_),
    .SN(_00850_));
 HAxp5_ASAP7_75t_R _34092_ (.A(_17568_),
    .B(_17569_),
    .CON(_02276_),
    .SN(_00882_));
 HAxp5_ASAP7_75t_R _34093_ (.A(_17570_),
    .B(_17571_),
    .CON(_00948_),
    .SN(_00915_));
 HAxp5_ASAP7_75t_R _34094_ (.A(_17572_),
    .B(_17573_),
    .CON(_02277_),
    .SN(_00947_));
 HAxp5_ASAP7_75t_R _34095_ (.A(_16532_),
    .B(_16533_),
    .CON(_01013_),
    .SN(_00980_));
 HAxp5_ASAP7_75t_R _34096_ (.A(_17574_),
    .B(_17575_),
    .CON(_02278_),
    .SN(_01012_));
 HAxp5_ASAP7_75t_R _34097_ (.A(_17576_),
    .B(_17577_),
    .CON(_01079_),
    .SN(_01046_));
 HAxp5_ASAP7_75t_R _34098_ (.A(_17578_),
    .B(_17579_),
    .CON(_02279_),
    .SN(_01078_));
 HAxp5_ASAP7_75t_R _34099_ (.A(_16538_),
    .B(_16539_),
    .CON(_01144_),
    .SN(_01111_));
 HAxp5_ASAP7_75t_R _34100_ (.A(_17580_),
    .B(_17581_),
    .CON(_02280_),
    .SN(_01143_));
 HAxp5_ASAP7_75t_R _34101_ (.A(_16540_),
    .B(_16542_),
    .CON(_01210_),
    .SN(_01177_));
 HAxp5_ASAP7_75t_R _34102_ (.A(_17582_),
    .B(_17583_),
    .CON(_02281_),
    .SN(_01209_));
 HAxp5_ASAP7_75t_R _34103_ (.A(_16543_),
    .B(_16544_),
    .CON(_01276_),
    .SN(_01243_));
 HAxp5_ASAP7_75t_R _34104_ (.A(_17584_),
    .B(_17585_),
    .CON(_01309_),
    .SN(_01275_));
 HAxp5_ASAP7_75t_R _34105_ (.A(_17586_),
    .B(_17587_),
    .CON(_02282_),
    .SN(_01310_));
 HAxp5_ASAP7_75t_R _34106_ (.A(_17588_),
    .B(_05478_),
    .CON(_00160_),
    .SN(_17590_));
 HAxp5_ASAP7_75t_R _34107_ (.A(_17591_),
    .B(_17592_),
    .CON(_02283_),
    .SN(_02284_));
 HAxp5_ASAP7_75t_R _34108_ (.A(_17593_),
    .B(\cs_registers_i.priv_lvl_q[0] ),
    .CON(_02285_),
    .SN(_01313_));
 HAxp5_ASAP7_75t_R _34109_ (.A(_17594_),
    .B(_14501_),
    .CON(_02286_),
    .SN(_02287_));
 HAxp5_ASAP7_75t_R _34110_ (.A(_17594_),
    .B(_14502_),
    .CON(_02288_),
    .SN(_17597_));
 HAxp5_ASAP7_75t_R _34111_ (.A(_17598_),
    .B(_14501_),
    .CON(_02289_),
    .SN(_17599_));
 HAxp5_ASAP7_75t_R _34112_ (.A(_17600_),
    .B(_17601_),
    .CON(_01321_),
    .SN(_02290_));
 HAxp5_ASAP7_75t_R _34113_ (.A(_17600_),
    .B(_17601_),
    .CON(_02291_),
    .SN(_17602_));
 HAxp5_ASAP7_75t_R _34114_ (.A(_17600_),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CON(_01326_),
    .SN(_17604_));
 HAxp5_ASAP7_75t_R _34115_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_17601_),
    .CON(_01319_),
    .SN(_17605_));
 HAxp5_ASAP7_75t_R _34116_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CON(_01320_),
    .SN(_17606_));
 HAxp5_ASAP7_75t_R _34117_ (.A(_17607_),
    .B(_17603_),
    .CON(_02292_),
    .SN(_02293_));
 HAxp5_ASAP7_75t_R _34118_ (.A(_17608_),
    .B(_17609_),
    .CON(_02294_),
    .SN(_01356_));
 HAxp5_ASAP7_75t_R _34119_ (.A(_17611_),
    .B(_17612_),
    .CON(_02295_),
    .SN(_01358_));
 HAxp5_ASAP7_75t_R _34120_ (.A(_17615_),
    .B(_17614_),
    .CON(_02296_),
    .SN(_01359_));
 HAxp5_ASAP7_75t_R _34121_ (.A(_17617_),
    .B(_17610_),
    .CON(_02297_),
    .SN(_01360_));
 HAxp5_ASAP7_75t_R _34122_ (.A(_17619_),
    .B(_17613_),
    .CON(_02298_),
    .SN(_01361_));
 HAxp5_ASAP7_75t_R _34123_ (.A(_17622_),
    .B(_17621_),
    .CON(_02299_),
    .SN(_01362_));
 HAxp5_ASAP7_75t_R _34124_ (.A(_17624_),
    .B(_17616_),
    .CON(_16553_),
    .SN(_01363_));
 HAxp5_ASAP7_75t_R _34125_ (.A(_17625_),
    .B(_17618_),
    .CON(_16554_),
    .SN(_01364_));
 HAxp5_ASAP7_75t_R _34126_ (.A(_17626_),
    .B(_17627_),
    .CON(_02300_),
    .SN(_01365_));
 HAxp5_ASAP7_75t_R _34127_ (.A(_17629_),
    .B(_17630_),
    .CON(_02301_),
    .SN(_01366_));
 HAxp5_ASAP7_75t_R _34128_ (.A(_17632_),
    .B(_17620_),
    .CON(_02302_),
    .SN(_01367_));
 HAxp5_ASAP7_75t_R _34129_ (.A(_17628_),
    .B(_17634_),
    .CON(_02303_),
    .SN(_01368_));
 HAxp5_ASAP7_75t_R _34130_ (.A(_17636_),
    .B(_17623_),
    .CON(_16565_),
    .SN(_16552_));
 HAxp5_ASAP7_75t_R _34131_ (.A(_17638_),
    .B(_17639_),
    .CON(_02304_),
    .SN(_01369_));
 HAxp5_ASAP7_75t_R _34132_ (.A(_17641_),
    .B(_17640_),
    .CON(_02305_),
    .SN(_01370_));
 HAxp5_ASAP7_75t_R _34133_ (.A(_17642_),
    .B(_17643_),
    .CON(_02306_),
    .SN(_01371_));
 HAxp5_ASAP7_75t_R _34134_ (.A(_17645_),
    .B(_17631_),
    .CON(_02307_),
    .SN(_01372_));
 HAxp5_ASAP7_75t_R _34135_ (.A(_17647_),
    .B(_17633_),
    .CON(_02308_),
    .SN(_01373_));
 HAxp5_ASAP7_75t_R _34136_ (.A(_16563_),
    .B(_17635_),
    .CON(_02309_),
    .SN(_16564_));
 HAxp5_ASAP7_75t_R _34137_ (.A(_17649_),
    .B(_17637_),
    .CON(_01386_),
    .SN(_01375_));
 HAxp5_ASAP7_75t_R _34138_ (.A(_17651_),
    .B(_16569_),
    .CON(_02310_),
    .SN(_01378_));
 HAxp5_ASAP7_75t_R _34139_ (.A(_16578_),
    .B(_17644_),
    .CON(_02311_),
    .SN(_01380_));
 HAxp5_ASAP7_75t_R _34140_ (.A(_17653_),
    .B(_17646_),
    .CON(_02312_),
    .SN(_01381_));
 HAxp5_ASAP7_75t_R _34141_ (.A(_16586_),
    .B(_17648_),
    .CON(_02313_),
    .SN(_01385_));
 HAxp5_ASAP7_75t_R _34142_ (.A(_17654_),
    .B(_16590_),
    .CON(_02314_),
    .SN(_01389_));
 HAxp5_ASAP7_75t_R _34143_ (.A(_17657_),
    .B(_17656_),
    .CON(_02315_),
    .SN(_01390_));
 HAxp5_ASAP7_75t_R _34144_ (.A(_17660_),
    .B(_16577_),
    .CON(_02316_),
    .SN(_01392_));
 HAxp5_ASAP7_75t_R _34145_ (.A(_17662_),
    .B(_17652_),
    .CON(_02317_),
    .SN(_01393_));
 HAxp5_ASAP7_75t_R _34146_ (.A(_16604_),
    .B(_16585_),
    .CON(_01411_),
    .SN(_01398_));
 HAxp5_ASAP7_75t_R _34147_ (.A(_17663_),
    .B(_17664_),
    .CON(_02318_),
    .SN(_01399_));
 HAxp5_ASAP7_75t_R _34148_ (.A(_17665_),
    .B(_16609_),
    .CON(_02319_),
    .SN(_01401_));
 HAxp5_ASAP7_75t_R _34149_ (.A(_17667_),
    .B(_17655_),
    .CON(_16642_),
    .SN(_01402_));
 HAxp5_ASAP7_75t_R _34150_ (.A(_17669_),
    .B(_17668_),
    .CON(_02320_),
    .SN(_01403_));
 HAxp5_ASAP7_75t_R _34151_ (.A(_17672_),
    .B(_17673_),
    .CON(_16644_),
    .SN(_01404_));
 HAxp5_ASAP7_75t_R _34152_ (.A(_17674_),
    .B(_17661_),
    .CON(_02321_),
    .SN(_01405_));
 HAxp5_ASAP7_75t_R _34153_ (.A(_16623_),
    .B(_16603_),
    .CON(_02322_),
    .SN(_01410_));
 HAxp5_ASAP7_75t_R _34154_ (.A(_16635_),
    .B(_17666_),
    .CON(_16669_),
    .SN(_01414_));
 HAxp5_ASAP7_75t_R _34155_ (.A(_17676_),
    .B(_17675_),
    .CON(_02323_),
    .SN(_01415_));
 HAxp5_ASAP7_75t_R _34156_ (.A(_17679_),
    .B(_17680_),
    .CON(_16671_),
    .SN(_16643_));
 HAxp5_ASAP7_75t_R _34157_ (.A(_16652_),
    .B(_16622_),
    .CON(_01427_),
    .SN(_01420_));
 HAxp5_ASAP7_75t_R _34158_ (.A(_17681_),
    .B(_17682_),
    .CON(_02324_),
    .SN(_01421_));
 HAxp5_ASAP7_75t_R _34159_ (.A(_17686_),
    .B(_16634_),
    .CON(_16697_),
    .SN(_01423_));
 HAxp5_ASAP7_75t_R _34160_ (.A(_17683_),
    .B(_17687_),
    .CON(_02325_),
    .SN(_01424_));
 HAxp5_ASAP7_75t_R _34161_ (.A(_17690_),
    .B(_17691_),
    .CON(_16699_),
    .SN(_16670_));
 HAxp5_ASAP7_75t_R _34162_ (.A(_17693_),
    .B(_16651_),
    .CON(_02326_),
    .SN(_01426_));
 HAxp5_ASAP7_75t_R _34163_ (.A(_17694_),
    .B(_17695_),
    .CON(_02327_),
    .SN(_01428_));
 HAxp5_ASAP7_75t_R _34164_ (.A(_17698_),
    .B(_17697_),
    .CON(_02328_),
    .SN(_01429_));
 HAxp5_ASAP7_75t_R _34165_ (.A(_17701_),
    .B(_17702_),
    .CON(_16730_),
    .SN(_01430_));
 HAxp5_ASAP7_75t_R _34166_ (.A(_17705_),
    .B(_17706_),
    .CON(_16732_),
    .SN(_16698_));
 HAxp5_ASAP7_75t_R _34167_ (.A(_16705_),
    .B(_16706_),
    .CON(_01437_),
    .SN(_01432_));
 HAxp5_ASAP7_75t_R _34168_ (.A(_17708_),
    .B(_17696_),
    .CON(_16754_),
    .SN(_01433_));
 HAxp5_ASAP7_75t_R _34169_ (.A(_17710_),
    .B(_17709_),
    .CON(_02329_),
    .SN(_01434_));
 HAxp5_ASAP7_75t_R _34170_ (.A(_17713_),
    .B(_17714_),
    .CON(_16764_),
    .SN(_01435_));
 HAxp5_ASAP7_75t_R _34171_ (.A(_17717_),
    .B(_17718_),
    .CON(_16766_),
    .SN(_16731_));
 HAxp5_ASAP7_75t_R _34172_ (.A(_17722_),
    .B(_17723_),
    .CON(_02330_),
    .SN(_01436_));
 HAxp5_ASAP7_75t_R _34173_ (.A(_17724_),
    .B(_17725_),
    .CON(_02331_),
    .SN(_01438_));
 HAxp5_ASAP7_75t_R _34174_ (.A(_17727_),
    .B(_17728_),
    .CON(_16795_),
    .SN(_01439_));
 HAxp5_ASAP7_75t_R _34175_ (.A(_17726_),
    .B(_17729_),
    .CON(_02332_),
    .SN(_01440_));
 HAxp5_ASAP7_75t_R _34176_ (.A(_17736_),
    .B(_17737_),
    .CON(_02333_),
    .SN(_16765_));
 HAxp5_ASAP7_75t_R _34177_ (.A(_16773_),
    .B(_16775_),
    .CON(_00016_),
    .SN(_00009_));
 HAxp5_ASAP7_75t_R _34178_ (.A(_17742_),
    .B(_17743_),
    .CON(_16821_),
    .SN(_00010_));
 HAxp5_ASAP7_75t_R _34179_ (.A(_17744_),
    .B(_17745_),
    .CON(_02334_),
    .SN(_00011_));
 HAxp5_ASAP7_75t_R _34180_ (.A(_17746_),
    .B(_17747_),
    .CON(_16837_),
    .SN(_00012_));
 HAxp5_ASAP7_75t_R _34181_ (.A(_17754_),
    .B(_17755_),
    .CON(_02335_),
    .SN(_00014_));
 HAxp5_ASAP7_75t_R _34182_ (.A(_17759_),
    .B(_17760_),
    .CON(_02336_),
    .SN(_00015_));
 HAxp5_ASAP7_75t_R _34183_ (.A(_17761_),
    .B(_17762_),
    .CON(_02337_),
    .SN(_00017_));
 HAxp5_ASAP7_75t_R _34184_ (.A(_17773_),
    .B(_17774_),
    .CON(_02338_),
    .SN(_00018_));
 HAxp5_ASAP7_75t_R _34185_ (.A(_16858_),
    .B(_16859_),
    .CON(_00025_),
    .SN(_00019_));
 HAxp5_ASAP7_75t_R _34186_ (.A(_17777_),
    .B(_17778_),
    .CON(_02339_),
    .SN(_00020_));
 HAxp5_ASAP7_75t_R _34187_ (.A(_17779_),
    .B(_16863_),
    .CON(_02340_),
    .SN(_00022_));
 HAxp5_ASAP7_75t_R _34188_ (.A(_17793_),
    .B(_17794_),
    .CON(_02341_),
    .SN(_00023_));
 HAxp5_ASAP7_75t_R _34189_ (.A(_17797_),
    .B(_17798_),
    .CON(_02342_),
    .SN(_00024_));
 HAxp5_ASAP7_75t_R _34190_ (.A(_17813_),
    .B(_17814_),
    .CON(_00032_),
    .SN(_00029_));
 HAxp5_ASAP7_75t_R _34191_ (.A(_17832_),
    .B(_17833_),
    .CON(_02343_),
    .SN(_17001_));
 HAxp5_ASAP7_75t_R _34192_ (.A(_17838_),
    .B(_17839_),
    .CON(_02344_),
    .SN(_00031_));
 HAxp5_ASAP7_75t_R _34193_ (.A(_17859_),
    .B(_17860_),
    .CON(_02345_),
    .SN(_00035_));
 HAxp5_ASAP7_75t_R _34194_ (.A(_17056_),
    .B(_17057_),
    .CON(_00039_),
    .SN(_00036_));
 HAxp5_ASAP7_75t_R _34195_ (.A(_17883_),
    .B(_17884_),
    .CON(_02346_),
    .SN(_00037_));
 HAxp5_ASAP7_75t_R _34196_ (.A(_17887_),
    .B(_17888_),
    .CON(_02347_),
    .SN(_00038_));
 HAxp5_ASAP7_75t_R _34197_ (.A(_17908_),
    .B(_17909_),
    .CON(_02348_),
    .SN(_00040_));
 HAxp5_ASAP7_75t_R _34198_ (.A(_17144_),
    .B(_17145_),
    .CON(_00045_),
    .SN(_00041_));
 HAxp5_ASAP7_75t_R _34199_ (.A(_17187_),
    .B(_17930_),
    .CON(_02349_),
    .SN(_00043_));
 HAxp5_ASAP7_75t_R _34200_ (.A(_17933_),
    .B(_17934_),
    .CON(_02350_),
    .SN(_00044_));
 HAxp5_ASAP7_75t_R _34201_ (.A(_17226_),
    .B(_17186_),
    .CON(_02351_),
    .SN(_00048_));
 HAxp5_ASAP7_75t_R _34202_ (.A(_17235_),
    .B(_17236_),
    .CON(_00053_),
    .SN(_00049_));
 HAxp5_ASAP7_75t_R _34203_ (.A(_17226_),
    .B(_17225_),
    .CON(_02352_),
    .SN(_00051_));
 HAxp5_ASAP7_75t_R _34204_ (.A(_17974_),
    .B(_17975_),
    .CON(_02353_),
    .SN(_00052_));
 HAxp5_ASAP7_75t_R _34205_ (.A(_17313_),
    .B(_17314_),
    .CON(_00056_),
    .SN(_00054_));
 HAxp5_ASAP7_75t_R _34206_ (.A(_18010_),
    .B(_18011_),
    .CON(_02354_),
    .SN(_00055_));
 HAxp5_ASAP7_75t_R _34207_ (.A(_17379_),
    .B(_17380_),
    .CON(_00059_),
    .SN(_00057_));
 HAxp5_ASAP7_75t_R _34208_ (.A(_18045_),
    .B(_18046_),
    .CON(_02355_),
    .SN(_00058_));
 HAxp5_ASAP7_75t_R _34209_ (.A(_17437_),
    .B(_17438_),
    .CON(_00062_),
    .SN(_00060_));
 HAxp5_ASAP7_75t_R _34210_ (.A(_18077_),
    .B(_18078_),
    .CON(_02356_),
    .SN(_00061_));
 HAxp5_ASAP7_75t_R _34211_ (.A(_17489_),
    .B(_17490_),
    .CON(_00065_),
    .SN(_00063_));
 HAxp5_ASAP7_75t_R _34212_ (.A(_18095_),
    .B(_18096_),
    .CON(_00067_),
    .SN(_00064_));
 HAxp5_ASAP7_75t_R _34213_ (.A(net290),
    .B(_13301_),
    .CON(_02357_),
    .SN(_00072_));
 HAxp5_ASAP7_75t_R _34214_ (.A(_13955_),
    .B(_18106_),
    .CON(_02358_),
    .SN(_00073_));
 HAxp5_ASAP7_75t_R _34215_ (.A(net290),
    .B(_18108_),
    .CON(_00074_),
    .SN(_02359_));
 HAxp5_ASAP7_75t_R _34216_ (.A(_13658_),
    .B(_13777_),
    .CON(_02360_),
    .SN(_18111_));
 HAxp5_ASAP7_75t_R _34217_ (.A(_13573_),
    .B(_13302_),
    .CON(_00076_),
    .SN(_00075_));
 HAxp5_ASAP7_75t_R _34218_ (.A(_18114_),
    .B(_13301_),
    .CON(_02361_),
    .SN(_18115_));
 HAxp5_ASAP7_75t_R _34219_ (.A(_13954_),
    .B(_18117_),
    .CON(_00078_),
    .SN(_00077_));
 HAxp5_ASAP7_75t_R _34220_ (.A(_13955_),
    .B(_14688_),
    .CON(_02362_),
    .SN(_18119_));
 HAxp5_ASAP7_75t_R _34221_ (.A(_14025_),
    .B(_18121_),
    .CON(_02363_),
    .SN(_00079_));
 HAxp5_ASAP7_75t_R _34222_ (.A(_14026_),
    .B(_14761_),
    .CON(_00080_),
    .SN(_18124_));
 HAxp5_ASAP7_75t_R _34223_ (.A(_14083_),
    .B(_14822_),
    .CON(_02364_),
    .SN(_00082_));
 HAxp5_ASAP7_75t_R _34224_ (.A(_14084_),
    .B(_18128_),
    .CON(_00083_),
    .SN(_18129_));
 HAxp5_ASAP7_75t_R _34225_ (.A(_14139_),
    .B(_18131_),
    .CON(_00086_),
    .SN(_00085_));
 HAxp5_ASAP7_75t_R _34226_ (.A(_14140_),
    .B(_18133_),
    .CON(_02365_),
    .SN(_18134_));
 HAxp5_ASAP7_75t_R _34227_ (.A(_18135_),
    .B(_14938_),
    .CON(_00089_),
    .SN(_00088_));
 HAxp5_ASAP7_75t_R _34228_ (.A(_18137_),
    .B(_18138_),
    .CON(_02366_),
    .SN(_18139_));
 HAxp5_ASAP7_75t_R _34229_ (.A(_14256_),
    .B(_18141_),
    .CON(_00092_),
    .SN(_00091_));
 HAxp5_ASAP7_75t_R _34230_ (.A(_18142_),
    .B(_18143_),
    .CON(_02367_),
    .SN(_18144_));
 HAxp5_ASAP7_75t_R _34231_ (.A(_14319_),
    .B(_18146_),
    .CON(_00094_),
    .SN(_00093_));
 HAxp5_ASAP7_75t_R _34232_ (.A(_18147_),
    .B(_18148_),
    .CON(_02368_),
    .SN(_18149_));
 HAxp5_ASAP7_75t_R _34233_ (.A(_14376_),
    .B(_15104_),
    .CON(_00097_),
    .SN(_00096_));
 HAxp5_ASAP7_75t_R _34234_ (.A(_18152_),
    .B(_18153_),
    .CON(_02369_),
    .SN(_18154_));
 HAxp5_ASAP7_75t_R _34235_ (.A(_18155_),
    .B(_15159_),
    .CON(_00100_),
    .SN(_00099_));
 HAxp5_ASAP7_75t_R _34236_ (.A(_18157_),
    .B(_18158_),
    .CON(_02370_),
    .SN(_18159_));
 HAxp5_ASAP7_75t_R _34237_ (.A(_14497_),
    .B(_14576_),
    .CON(_02371_),
    .SN(_00102_));
 HAxp5_ASAP7_75t_R _34238_ (.A(_18162_),
    .B(_18163_),
    .CON(_00103_),
    .SN(_18164_));
 HAxp5_ASAP7_75t_R _34239_ (.A(_18165_),
    .B(_18166_),
    .CON(_00105_),
    .SN(_00104_));
 HAxp5_ASAP7_75t_R _34240_ (.A(_18167_),
    .B(_18168_),
    .CON(_02372_),
    .SN(_18169_));
 HAxp5_ASAP7_75t_R _34241_ (.A(_18170_),
    .B(_18171_),
    .CON(_00107_),
    .SN(_00106_));
 HAxp5_ASAP7_75t_R _34242_ (.A(_15407_),
    .B(_18173_),
    .CON(_02373_),
    .SN(_18174_));
 HAxp5_ASAP7_75t_R _34243_ (.A(_18175_),
    .B(_15556_),
    .CON(_02374_),
    .SN(_00109_));
 HAxp5_ASAP7_75t_R _34244_ (.A(_18177_),
    .B(_18178_),
    .CON(_00110_),
    .SN(_18179_));
 HAxp5_ASAP7_75t_R _34245_ (.A(_15668_),
    .B(_18181_),
    .CON(_00113_),
    .SN(_00112_));
 HAxp5_ASAP7_75t_R _34246_ (.A(_18182_),
    .B(_15620_),
    .CON(_02375_),
    .SN(_18184_));
 HAxp5_ASAP7_75t_R _34247_ (.A(_18185_),
    .B(_18186_),
    .CON(_02376_),
    .SN(_00115_));
 HAxp5_ASAP7_75t_R _34248_ (.A(_18187_),
    .B(_15781_),
    .CON(_00116_),
    .SN(_18189_));
 HAxp5_ASAP7_75t_R _34249_ (.A(_18190_),
    .B(_15897_),
    .CON(_02377_),
    .SN(_00118_));
 HAxp5_ASAP7_75t_R _34250_ (.A(_18192_),
    .B(_18193_),
    .CON(_00119_),
    .SN(_18194_));
 HAxp5_ASAP7_75t_R _34251_ (.A(_18195_),
    .B(_18196_),
    .CON(_02378_),
    .SN(_00121_));
 HAxp5_ASAP7_75t_R _34252_ (.A(_18197_),
    .B(_18198_),
    .CON(_00122_),
    .SN(_18199_));
 HAxp5_ASAP7_75t_R _34253_ (.A(_18200_),
    .B(_18201_),
    .CON(_00125_),
    .SN(_00124_));
 HAxp5_ASAP7_75t_R _34254_ (.A(_16137_),
    .B(_18203_),
    .CON(_02379_),
    .SN(_18204_));
 HAxp5_ASAP7_75t_R _34255_ (.A(_18205_),
    .B(_18206_),
    .CON(_02380_),
    .SN(_00127_));
 HAxp5_ASAP7_75t_R _34256_ (.A(_18207_),
    .B(_16259_),
    .CON(_00128_),
    .SN(_18209_));
 HAxp5_ASAP7_75t_R _34257_ (.A(_16326_),
    .B(_18211_),
    .CON(_02381_),
    .SN(_00130_));
 HAxp5_ASAP7_75t_R _34258_ (.A(_18212_),
    .B(_18213_),
    .CON(_00131_),
    .SN(_18214_));
 HAxp5_ASAP7_75t_R _34259_ (.A(_18215_),
    .B(_18216_),
    .CON(_00134_),
    .SN(_00133_));
 HAxp5_ASAP7_75t_R _34260_ (.A(_16480_),
    .B(_18218_),
    .CON(_02382_),
    .SN(_18219_));
 HAxp5_ASAP7_75t_R _34261_ (.A(_04603_),
    .B(_18221_),
    .CON(_00137_),
    .SN(_00136_));
 HAxp5_ASAP7_75t_R _34262_ (.A(_18222_),
    .B(_18223_),
    .CON(_02383_),
    .SN(_18224_));
 HAxp5_ASAP7_75t_R _34263_ (.A(_18225_),
    .B(_18226_),
    .CON(_02384_),
    .SN(_00139_));
 HAxp5_ASAP7_75t_R _34264_ (.A(_18227_),
    .B(_04718_),
    .CON(_00140_),
    .SN(_18229_));
 HAxp5_ASAP7_75t_R _34265_ (.A(_04782_),
    .B(_18231_),
    .CON(_02385_),
    .SN(_00142_));
 HAxp5_ASAP7_75t_R _34266_ (.A(_18232_),
    .B(_04829_),
    .CON(_00143_),
    .SN(_18234_));
 HAxp5_ASAP7_75t_R _34267_ (.A(_18235_),
    .B(_18236_),
    .CON(_00146_),
    .SN(_00145_));
 HAxp5_ASAP7_75t_R _34268_ (.A(_18237_),
    .B(_18238_),
    .CON(_02386_),
    .SN(_18239_));
 HAxp5_ASAP7_75t_R _34269_ (.A(_05045_),
    .B(_18241_),
    .CON(_00149_),
    .SN(_00148_));
 HAxp5_ASAP7_75t_R _34270_ (.A(_18242_),
    .B(_04998_),
    .CON(_02387_),
    .SN(_18244_));
 HAxp5_ASAP7_75t_R _34271_ (.A(_05107_),
    .B(_18246_),
    .CON(_02388_),
    .SN(_00151_));
 HAxp5_ASAP7_75t_R _34272_ (.A(_18247_),
    .B(_18248_),
    .CON(_00152_),
    .SN(_18249_));
 HAxp5_ASAP7_75t_R _34273_ (.A(_05215_),
    .B(_18251_),
    .CON(_02389_),
    .SN(_00154_));
 HAxp5_ASAP7_75t_R _34274_ (.A(_18252_),
    .B(_18253_),
    .CON(_00155_),
    .SN(_18254_));
 HAxp5_ASAP7_75t_R _34275_ (.A(_05325_),
    .B(_18256_),
    .CON(_02390_),
    .SN(_00157_));
 HAxp5_ASAP7_75t_R _34276_ (.A(_18257_),
    .B(_05371_),
    .CON(_00158_),
    .SN(_18259_));
 HAxp5_ASAP7_75t_R _34277_ (.A(\cs_registers_i.mhpmcounter[2][0] ),
    .B(\cs_registers_i.mhpmcounter[2][1] ),
    .CON(_02391_),
    .SN(_02392_));
 HAxp5_ASAP7_75t_R _34278_ (.A(\cs_registers_i.mhpmcounter[2][2] ),
    .B(_18260_),
    .CON(_02393_),
    .SN(_02394_));
 HAxp5_ASAP7_75t_R _34279_ (.A(\cs_registers_i.mhpmcounter[2][4] ),
    .B(_18261_),
    .CON(_02395_),
    .SN(_02396_));
 HAxp5_ASAP7_75t_R _34280_ (.A(\cs_registers_i.mhpmcounter[2][6] ),
    .B(_18262_),
    .CON(_02397_),
    .SN(_02398_));
 HAxp5_ASAP7_75t_R _34281_ (.A(\cs_registers_i.mhpmcounter[2][8] ),
    .B(_18263_),
    .CON(_02399_),
    .SN(_02400_));
 HAxp5_ASAP7_75t_R _34282_ (.A(\cs_registers_i.mhpmcounter[2][10] ),
    .B(_18264_),
    .CON(_02401_),
    .SN(_02402_));
 HAxp5_ASAP7_75t_R _34283_ (.A(\cs_registers_i.mhpmcounter[2][12] ),
    .B(_18265_),
    .CON(_02403_),
    .SN(_02404_));
 HAxp5_ASAP7_75t_R _34284_ (.A(\cs_registers_i.mhpmcounter[2][14] ),
    .B(_18266_),
    .CON(_02405_),
    .SN(_02406_));
 HAxp5_ASAP7_75t_R _34285_ (.A(\cs_registers_i.mhpmcounter[2][16] ),
    .B(_18267_),
    .CON(_02407_),
    .SN(_02408_));
 HAxp5_ASAP7_75t_R _34286_ (.A(\cs_registers_i.mhpmcounter[2][18] ),
    .B(_18268_),
    .CON(_02409_),
    .SN(_02410_));
 HAxp5_ASAP7_75t_R _34287_ (.A(\cs_registers_i.mhpmcounter[2][20] ),
    .B(_18269_),
    .CON(_02411_),
    .SN(_02412_));
 HAxp5_ASAP7_75t_R _34288_ (.A(\cs_registers_i.mhpmcounter[2][22] ),
    .B(_18270_),
    .CON(_02413_),
    .SN(_02414_));
 HAxp5_ASAP7_75t_R _34289_ (.A(\cs_registers_i.mhpmcounter[2][24] ),
    .B(_18271_),
    .CON(_02415_),
    .SN(_02416_));
 HAxp5_ASAP7_75t_R _34290_ (.A(\cs_registers_i.mhpmcounter[2][26] ),
    .B(_18272_),
    .CON(_02417_),
    .SN(_02418_));
 HAxp5_ASAP7_75t_R _34291_ (.A(\cs_registers_i.mhpmcounter[2][28] ),
    .B(_18273_),
    .CON(_02419_),
    .SN(_02420_));
 HAxp5_ASAP7_75t_R _34292_ (.A(\cs_registers_i.mhpmcounter[2][30] ),
    .B(_18274_),
    .CON(_02421_),
    .SN(_02422_));
 HAxp5_ASAP7_75t_R _34293_ (.A(\cs_registers_i.mhpmcounter[2][32] ),
    .B(_18275_),
    .CON(_02423_),
    .SN(_02424_));
 HAxp5_ASAP7_75t_R _34294_ (.A(\cs_registers_i.mhpmcounter[2][34] ),
    .B(_18276_),
    .CON(_02425_),
    .SN(_02426_));
 HAxp5_ASAP7_75t_R _34295_ (.A(\cs_registers_i.mhpmcounter[2][36] ),
    .B(_18277_),
    .CON(_02427_),
    .SN(_02428_));
 HAxp5_ASAP7_75t_R _34296_ (.A(\cs_registers_i.mhpmcounter[2][38] ),
    .B(_18278_),
    .CON(_02429_),
    .SN(_02430_));
 HAxp5_ASAP7_75t_R _34297_ (.A(\cs_registers_i.mhpmcounter[2][40] ),
    .B(_18279_),
    .CON(_02431_),
    .SN(_02432_));
 HAxp5_ASAP7_75t_R _34298_ (.A(\cs_registers_i.mhpmcounter[2][42] ),
    .B(_18280_),
    .CON(_02433_),
    .SN(_02434_));
 HAxp5_ASAP7_75t_R _34299_ (.A(\cs_registers_i.mhpmcounter[2][44] ),
    .B(_18281_),
    .CON(_02435_),
    .SN(_02436_));
 HAxp5_ASAP7_75t_R _34300_ (.A(\cs_registers_i.mhpmcounter[2][46] ),
    .B(_18282_),
    .CON(_02437_),
    .SN(_02438_));
 HAxp5_ASAP7_75t_R _34301_ (.A(\cs_registers_i.mhpmcounter[2][48] ),
    .B(_18283_),
    .CON(_02439_),
    .SN(_02440_));
 HAxp5_ASAP7_75t_R _34302_ (.A(\cs_registers_i.mhpmcounter[2][50] ),
    .B(_18284_),
    .CON(_02441_),
    .SN(_02442_));
 HAxp5_ASAP7_75t_R _34303_ (.A(\cs_registers_i.mhpmcounter[2][52] ),
    .B(_18285_),
    .CON(_02443_),
    .SN(_02444_));
 HAxp5_ASAP7_75t_R _34304_ (.A(\cs_registers_i.mhpmcounter[2][54] ),
    .B(_18286_),
    .CON(_02445_),
    .SN(_02446_));
 HAxp5_ASAP7_75t_R _34305_ (.A(\cs_registers_i.mhpmcounter[2][56] ),
    .B(_18287_),
    .CON(_02447_),
    .SN(_02448_));
 HAxp5_ASAP7_75t_R _34306_ (.A(\cs_registers_i.mhpmcounter[2][58] ),
    .B(_18288_),
    .CON(_02449_),
    .SN(_02450_));
 HAxp5_ASAP7_75t_R _34307_ (.A(\cs_registers_i.mhpmcounter[2][60] ),
    .B(_18289_),
    .CON(_02451_),
    .SN(_02452_));
 HAxp5_ASAP7_75t_R _34308_ (.A(\cs_registers_i.mhpmcounter[2][62] ),
    .B(_18290_),
    .CON(_02453_),
    .SN(_02454_));
 HAxp5_ASAP7_75t_R _34309_ (.A(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .CON(_02455_),
    .SN(_02456_));
 HAxp5_ASAP7_75t_R _34310_ (.A(\cs_registers_i.mcycle_counter_i.counter[2] ),
    .B(_18291_),
    .CON(_02457_),
    .SN(_02458_));
 HAxp5_ASAP7_75t_R _34311_ (.A(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .B(_18292_),
    .CON(_02459_),
    .SN(_02460_));
 HAxp5_ASAP7_75t_R _34312_ (.A(\cs_registers_i.mcycle_counter_i.counter[6] ),
    .B(_18293_),
    .CON(_02461_),
    .SN(_02462_));
 HAxp5_ASAP7_75t_R _34313_ (.A(\cs_registers_i.mcycle_counter_i.counter[8] ),
    .B(_18294_),
    .CON(_02463_),
    .SN(_02464_));
 HAxp5_ASAP7_75t_R _34314_ (.A(\cs_registers_i.mcycle_counter_i.counter[10] ),
    .B(_18295_),
    .CON(_02465_),
    .SN(_02466_));
 HAxp5_ASAP7_75t_R _34315_ (.A(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .B(_18296_),
    .CON(_02467_),
    .SN(_02468_));
 HAxp5_ASAP7_75t_R _34316_ (.A(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .B(_18297_),
    .CON(_02469_),
    .SN(_02470_));
 HAxp5_ASAP7_75t_R _34317_ (.A(\cs_registers_i.mcycle_counter_i.counter[16] ),
    .B(_18298_),
    .CON(_02471_),
    .SN(_02472_));
 HAxp5_ASAP7_75t_R _34318_ (.A(\cs_registers_i.mcycle_counter_i.counter[18] ),
    .B(_18299_),
    .CON(_02473_),
    .SN(_02474_));
 HAxp5_ASAP7_75t_R _34319_ (.A(\cs_registers_i.mcycle_counter_i.counter[20] ),
    .B(_18300_),
    .CON(_02475_),
    .SN(_02476_));
 HAxp5_ASAP7_75t_R _34320_ (.A(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .B(_18301_),
    .CON(_02477_),
    .SN(_02478_));
 HAxp5_ASAP7_75t_R _34321_ (.A(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .B(_18302_),
    .CON(_02479_),
    .SN(_02480_));
 HAxp5_ASAP7_75t_R _34322_ (.A(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .B(_18303_),
    .CON(_02481_),
    .SN(_02482_));
 HAxp5_ASAP7_75t_R _34323_ (.A(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .B(_18304_),
    .CON(_02483_),
    .SN(_02484_));
 HAxp5_ASAP7_75t_R _34324_ (.A(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .B(_18305_),
    .CON(_02485_),
    .SN(_02486_));
 HAxp5_ASAP7_75t_R _34325_ (.A(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .B(_18306_),
    .CON(_02487_),
    .SN(_02488_));
 HAxp5_ASAP7_75t_R _34326_ (.A(\cs_registers_i.mcycle_counter_i.counter[34] ),
    .B(_18307_),
    .CON(_02489_),
    .SN(_02490_));
 HAxp5_ASAP7_75t_R _34327_ (.A(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .B(_18308_),
    .CON(_02491_),
    .SN(_02492_));
 HAxp5_ASAP7_75t_R _34328_ (.A(\cs_registers_i.mcycle_counter_i.counter[38] ),
    .B(_18309_),
    .CON(_02493_),
    .SN(_02494_));
 HAxp5_ASAP7_75t_R _34329_ (.A(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .B(_18310_),
    .CON(_02495_),
    .SN(_02496_));
 HAxp5_ASAP7_75t_R _34330_ (.A(\cs_registers_i.mcycle_counter_i.counter[42] ),
    .B(_18311_),
    .CON(_02497_),
    .SN(_02498_));
 HAxp5_ASAP7_75t_R _34331_ (.A(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .B(_18312_),
    .CON(_02499_),
    .SN(_02500_));
 HAxp5_ASAP7_75t_R _34332_ (.A(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .B(_18313_),
    .CON(_02501_),
    .SN(_02502_));
 HAxp5_ASAP7_75t_R _34333_ (.A(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .B(_18314_),
    .CON(_02503_),
    .SN(_02504_));
 HAxp5_ASAP7_75t_R _34334_ (.A(\cs_registers_i.mcycle_counter_i.counter[50] ),
    .B(_18315_),
    .CON(_02505_),
    .SN(_02506_));
 HAxp5_ASAP7_75t_R _34335_ (.A(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .B(_18316_),
    .CON(_02507_),
    .SN(_02508_));
 HAxp5_ASAP7_75t_R _34336_ (.A(\cs_registers_i.mcycle_counter_i.counter[54] ),
    .B(_18317_),
    .CON(_02509_),
    .SN(_02510_));
 HAxp5_ASAP7_75t_R _34337_ (.A(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .B(_18318_),
    .CON(_02511_),
    .SN(_02512_));
 HAxp5_ASAP7_75t_R _34338_ (.A(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .B(_18319_),
    .CON(_02513_),
    .SN(_02514_));
 HAxp5_ASAP7_75t_R _34339_ (.A(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .B(_18320_),
    .CON(_02515_),
    .SN(_02516_));
 HAxp5_ASAP7_75t_R _34340_ (.A(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .B(_18321_),
    .CON(_02517_),
    .SN(_02518_));
 HAxp5_ASAP7_75t_R _34341_ (.A(\cs_registers_i.pc_id_i[1] ),
    .B(\cs_registers_i.pc_id_i[2] ),
    .CON(_02519_),
    .SN(_00167_));
 HAxp5_ASAP7_75t_R _34342_ (.A(\cs_registers_i.pc_id_i[3] ),
    .B(_18322_),
    .CON(_02520_),
    .SN(_00171_));
 HAxp5_ASAP7_75t_R _34343_ (.A(\cs_registers_i.pc_id_i[5] ),
    .B(_18323_),
    .CON(_02521_),
    .SN(_00178_));
 HAxp5_ASAP7_75t_R _34344_ (.A(\cs_registers_i.pc_id_i[7] ),
    .B(_18324_),
    .CON(_02522_),
    .SN(_00183_));
 HAxp5_ASAP7_75t_R _34345_ (.A(\cs_registers_i.pc_id_i[9] ),
    .B(_18325_),
    .CON(_02523_),
    .SN(_00190_));
 HAxp5_ASAP7_75t_R _34346_ (.A(\cs_registers_i.pc_id_i[11] ),
    .B(_18326_),
    .CON(_02524_),
    .SN(_00197_));
 HAxp5_ASAP7_75t_R _34347_ (.A(\cs_registers_i.pc_id_i[13] ),
    .B(_18327_),
    .CON(_02525_),
    .SN(_00202_));
 HAxp5_ASAP7_75t_R _34348_ (.A(\cs_registers_i.pc_id_i[15] ),
    .B(_18328_),
    .CON(_02526_),
    .SN(_00207_));
 HAxp5_ASAP7_75t_R _34349_ (.A(\cs_registers_i.pc_id_i[17] ),
    .B(_18329_),
    .CON(_02527_),
    .SN(_00210_));
 HAxp5_ASAP7_75t_R _34350_ (.A(\cs_registers_i.pc_id_i[19] ),
    .B(_18330_),
    .CON(_02528_),
    .SN(_00213_));
 HAxp5_ASAP7_75t_R _34351_ (.A(\cs_registers_i.pc_id_i[21] ),
    .B(_18331_),
    .CON(_02529_),
    .SN(_00216_));
 HAxp5_ASAP7_75t_R _34352_ (.A(\cs_registers_i.pc_id_i[23] ),
    .B(_18332_),
    .CON(_02530_),
    .SN(_00219_));
 HAxp5_ASAP7_75t_R _34353_ (.A(\cs_registers_i.pc_id_i[25] ),
    .B(_18333_),
    .CON(_02531_),
    .SN(_00222_));
 HAxp5_ASAP7_75t_R _34354_ (.A(\cs_registers_i.pc_id_i[27] ),
    .B(_18334_),
    .CON(_02532_),
    .SN(_00225_));
 HAxp5_ASAP7_75t_R _34355_ (.A(\cs_registers_i.pc_id_i[29] ),
    .B(_18335_),
    .CON(_02533_),
    .SN(_00228_));
 HAxp5_ASAP7_75t_R _34356_ (.A(_18336_),
    .B(_18337_),
    .CON(_02534_),
    .SN(_02535_));
 HAxp5_ASAP7_75t_R _34357_ (.A(\ex_block_i.alu_adder_result_ex_o[1] ),
    .B(_18336_),
    .CON(_00236_),
    .SN(_02536_));
 HAxp5_ASAP7_75t_R _34358_ (.A(_16499_),
    .B(_18336_),
    .CON(_00233_),
    .SN(_18338_));
 HAxp5_ASAP7_75t_R _34359_ (.A(\ex_block_i.alu_adder_result_ex_o[1] ),
    .B(net280),
    .CON(_00234_),
    .SN(_00235_));
 HAxp5_ASAP7_75t_R _34360_ (.A(\ex_block_i.alu_adder_result_ex_o[1] ),
    .B(net280),
    .CON(_02537_),
    .SN(_18339_));
 HAxp5_ASAP7_75t_R _34361_ (.A(\ex_block_i.alu_adder_result_ex_o[1] ),
    .B(_16503_),
    .CON(_00231_),
    .SN(_18340_));
 HAxp5_ASAP7_75t_R _34362_ (.A(_16499_),
    .B(net280),
    .CON(_00232_),
    .SN(_18341_));
 HAxp5_ASAP7_75t_R _34363_ (.A(_16499_),
    .B(_16503_),
    .CON(_18337_),
    .SN(_18342_));
 HAxp5_ASAP7_75t_R _34364_ (.A(_17535_),
    .B(\cs_registers_i.pc_if_i[3] ),
    .CON(_02538_),
    .SN(_02539_));
 HAxp5_ASAP7_75t_R _34365_ (.A(_18343_),
    .B(\cs_registers_i.pc_if_i[5] ),
    .CON(_02540_),
    .SN(_02541_));
 HAxp5_ASAP7_75t_R _34366_ (.A(_18344_),
    .B(\cs_registers_i.pc_if_i[7] ),
    .CON(_02542_),
    .SN(_02543_));
 HAxp5_ASAP7_75t_R _34367_ (.A(_18345_),
    .B(\cs_registers_i.pc_if_i[9] ),
    .CON(_02544_),
    .SN(_02545_));
 HAxp5_ASAP7_75t_R _34368_ (.A(_18346_),
    .B(\cs_registers_i.pc_if_i[11] ),
    .CON(_02546_),
    .SN(_02547_));
 HAxp5_ASAP7_75t_R _34369_ (.A(_18347_),
    .B(\cs_registers_i.pc_if_i[13] ),
    .CON(_02548_),
    .SN(_02549_));
 HAxp5_ASAP7_75t_R _34370_ (.A(_18348_),
    .B(\cs_registers_i.pc_if_i[15] ),
    .CON(_02550_),
    .SN(_02551_));
 HAxp5_ASAP7_75t_R _34371_ (.A(_18349_),
    .B(\cs_registers_i.pc_if_i[17] ),
    .CON(_02552_),
    .SN(_02553_));
 HAxp5_ASAP7_75t_R _34372_ (.A(_18350_),
    .B(\cs_registers_i.pc_if_i[19] ),
    .CON(_02554_),
    .SN(_02555_));
 HAxp5_ASAP7_75t_R _34373_ (.A(_18351_),
    .B(\cs_registers_i.pc_if_i[21] ),
    .CON(_02556_),
    .SN(_02557_));
 HAxp5_ASAP7_75t_R _34374_ (.A(_18352_),
    .B(\cs_registers_i.pc_if_i[23] ),
    .CON(_02558_),
    .SN(_02559_));
 HAxp5_ASAP7_75t_R _34375_ (.A(_18353_),
    .B(\cs_registers_i.pc_if_i[25] ),
    .CON(_02560_),
    .SN(_02561_));
 HAxp5_ASAP7_75t_R _34376_ (.A(_18354_),
    .B(\cs_registers_i.pc_if_i[27] ),
    .CON(_02562_),
    .SN(_02563_));
 HAxp5_ASAP7_75t_R _34377_ (.A(_18355_),
    .B(\cs_registers_i.pc_if_i[29] ),
    .CON(_02564_),
    .SN(_02565_));
 HAxp5_ASAP7_75t_R _34378_ (.A(_18356_),
    .B(_18357_),
    .CON(_02566_),
    .SN(_02567_));
 HAxp5_ASAP7_75t_R _34379_ (.A(_18358_),
    .B(_18359_),
    .CON(_02568_),
    .SN(_02569_));
 HAxp5_ASAP7_75t_R _34380_ (.A(_18360_),
    .B(_18361_),
    .CON(_02570_),
    .SN(_02571_));
 HAxp5_ASAP7_75t_R _34381_ (.A(_18362_),
    .B(_18363_),
    .CON(_02572_),
    .SN(_02573_));
 HAxp5_ASAP7_75t_R _34382_ (.A(_18364_),
    .B(_18365_),
    .CON(_02574_),
    .SN(_02575_));
 HAxp5_ASAP7_75t_R _34383_ (.A(_18366_),
    .B(_18367_),
    .CON(_02576_),
    .SN(_02577_));
 HAxp5_ASAP7_75t_R _34384_ (.A(_18368_),
    .B(_18369_),
    .CON(_02578_),
    .SN(_02579_));
 HAxp5_ASAP7_75t_R _34385_ (.A(_18370_),
    .B(_18371_),
    .CON(_02580_),
    .SN(_02581_));
 HAxp5_ASAP7_75t_R _34386_ (.A(_18372_),
    .B(_18373_),
    .CON(_02582_),
    .SN(_02583_));
 HAxp5_ASAP7_75t_R _34387_ (.A(_18374_),
    .B(_18375_),
    .CON(_02584_),
    .SN(_02585_));
 HAxp5_ASAP7_75t_R _34388_ (.A(_18376_),
    .B(_18377_),
    .CON(_02586_),
    .SN(_02587_));
 HAxp5_ASAP7_75t_R _34389_ (.A(_18378_),
    .B(_18379_),
    .CON(_02588_),
    .SN(_02589_));
 HAxp5_ASAP7_75t_R _34390_ (.A(_18380_),
    .B(_18381_),
    .CON(_02590_),
    .SN(_02591_));
 HAxp5_ASAP7_75t_R _34391_ (.A(_18382_),
    .B(_18383_),
    .CON(_02592_),
    .SN(_02593_));
 HAxp5_ASAP7_75t_R _34392_ (.A(_18384_),
    .B(_18385_),
    .CON(_02594_),
    .SN(_02595_));
 HAxp5_ASAP7_75t_R _34393_ (.A(_18386_),
    .B(_18387_),
    .CON(_00243_),
    .SN(_02596_));
 DFFHQNx1_ASAP7_75t_R _34394_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02597_),
    .QN(_01723_));
 DFFHQNx1_ASAP7_75t_R _34395_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02598_),
    .QN(_00164_));
 DFFHQNx1_ASAP7_75t_R _34396_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02599_),
    .QN(_00166_));
 DFFHQNx1_ASAP7_75t_R _34397_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02600_),
    .QN(_00169_));
 DFFHQNx1_ASAP7_75t_R _34398_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02601_),
    .QN(_00173_));
 DFFHQNx1_ASAP7_75t_R _34399_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02602_),
    .QN(_00176_));
 DFFHQNx1_ASAP7_75t_R _34400_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02603_),
    .QN(_00179_));
 DFFHQNx1_ASAP7_75t_R _34401_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02604_),
    .QN(_00181_));
 DFFHQNx1_ASAP7_75t_R _34402_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02605_),
    .QN(_00185_));
 DFFHQNx1_ASAP7_75t_R _34403_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02606_),
    .QN(_00188_));
 DFFHQNx1_ASAP7_75t_R _34404_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02607_),
    .QN(_00192_));
 DFFHQNx1_ASAP7_75t_R _34405_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02608_),
    .QN(_00195_));
 DFFHQNx1_ASAP7_75t_R _34406_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02609_),
    .QN(_00198_));
 DFFHQNx1_ASAP7_75t_R _34407_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02610_),
    .QN(_00200_));
 DFFHQNx1_ASAP7_75t_R _34408_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02611_),
    .QN(_00203_));
 DFFHQNx1_ASAP7_75t_R _34409_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02612_),
    .QN(_00205_));
 DFFHQNx1_ASAP7_75t_R _34410_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02613_),
    .QN(_00385_));
 DFFHQNx1_ASAP7_75t_R _34411_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02614_),
    .QN(_01722_));
 DFFHQNx1_ASAP7_75t_R _34412_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02615_),
    .QN(_01721_));
 DFFHQNx1_ASAP7_75t_R _34413_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02616_),
    .QN(_01720_));
 DFFHQNx1_ASAP7_75t_R _34414_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02617_),
    .QN(_00162_));
 DFFHQNx1_ASAP7_75t_R _34415_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02618_),
    .QN(_00170_));
 DFFHQNx1_ASAP7_75t_R _34416_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02619_),
    .QN(_00174_));
 DFFHQNx1_ASAP7_75t_R _34417_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02620_),
    .QN(_00177_));
 DFFHQNx1_ASAP7_75t_R _34418_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02621_),
    .QN(_00180_));
 DFFHQNx1_ASAP7_75t_R _34419_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02622_),
    .QN(_00182_));
 DFFHQNx1_ASAP7_75t_R _34420_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02623_),
    .QN(_00186_));
 DFFHQNx1_ASAP7_75t_R _34421_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02624_),
    .QN(_00189_));
 DFFHQNx1_ASAP7_75t_R _34422_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02625_),
    .QN(_00193_));
 DFFHQNx1_ASAP7_75t_R _34423_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02626_),
    .QN(_00196_));
 DFFHQNx1_ASAP7_75t_R _34424_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02627_),
    .QN(_00199_));
 DFFHQNx1_ASAP7_75t_R _34425_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02628_),
    .QN(_00201_));
 DFFHQNx1_ASAP7_75t_R _34426_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02629_),
    .QN(_00204_));
 DFFHQNx1_ASAP7_75t_R _34427_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02630_),
    .QN(_00206_));
 DFFHQNx1_ASAP7_75t_R _34428_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02631_),
    .QN(_00208_));
 DFFHQNx1_ASAP7_75t_R _34429_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02632_),
    .QN(_00209_));
 DFFHQNx1_ASAP7_75t_R _34430_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02633_),
    .QN(_00211_));
 DFFHQNx1_ASAP7_75t_R _34431_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02634_),
    .QN(_00212_));
 DFFHQNx1_ASAP7_75t_R _34432_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02635_),
    .QN(_00214_));
 DFFHQNx1_ASAP7_75t_R _34433_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_02636_),
    .QN(_00215_));
 DFFHQNx1_ASAP7_75t_R _34434_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02637_),
    .QN(_00217_));
 DFFHQNx1_ASAP7_75t_R _34435_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_02638_),
    .QN(_00218_));
 DFFHQNx1_ASAP7_75t_R _34436_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_02639_),
    .QN(_00220_));
 DFFHQNx1_ASAP7_75t_R _34437_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_02640_),
    .QN(_00221_));
 DFFHQNx1_ASAP7_75t_R _34438_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02641_),
    .QN(_00223_));
 DFFHQNx1_ASAP7_75t_R _34439_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_02642_),
    .QN(_00224_));
 DFFHQNx1_ASAP7_75t_R _34440_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02643_),
    .QN(_00226_));
 DFFHQNx1_ASAP7_75t_R _34441_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02644_),
    .QN(_00227_));
 DFFHQNx1_ASAP7_75t_R _34442_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02645_),
    .QN(_00229_));
 DFFHQNx1_ASAP7_75t_R _34443_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02646_),
    .QN(_00230_));
 DFFASRHQNx1_ASAP7_75t_R _34444_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.instr_valid_id_d ),
    .QN(_01317_),
    .RESETN(net456),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _34445_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(\id_stage_i.controller_i.illegal_insn_d ),
    .QN(_01312_),
    .RESETN(net457),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _34446_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(\id_stage_i.controller_i.exc_req_d ),
    .QN(_01724_),
    .RESETN(net458),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _34447_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(\id_stage_i.controller_i.store_err_d ),
    .QN(_01725_),
    .RESETN(net459),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34448_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(\id_stage_i.controller_i.load_err_d ),
    .QN(_01719_),
    .RESETN(net460),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34449_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_02647_),
    .QN(_01718_),
    .RESETN(net461),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34450_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02648_),
    .QN(_01717_),
    .RESETN(net462),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _34451_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02649_),
    .QN(_01716_),
    .RESETN(net463),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _34452_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02650_),
    .QN(_01715_),
    .RESETN(net464),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _34453_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02651_),
    .QN(_01714_),
    .RESETN(net465),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _34454_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02652_),
    .QN(_01713_),
    .RESETN(net466),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34455_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02653_),
    .QN(_01712_),
    .RESETN(net467),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _34456_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02654_),
    .QN(_01711_),
    .RESETN(net468),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _34457_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02655_),
    .QN(_01726_),
    .RESETN(net469),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34458_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(\id_stage_i.branch_set_d ),
    .QN(_01710_),
    .RESETN(net470),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34459_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_02656_),
    .QN(_01709_),
    .RESETN(net471),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34460_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_02657_),
    .QN(_01708_),
    .RESETN(net472),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34461_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_02658_),
    .QN(_01707_),
    .RESETN(net473),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _34462_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_02659_),
    .QN(_01706_),
    .RESETN(net474),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34463_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_02660_),
    .QN(_01705_),
    .RESETN(net475),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34464_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_02661_),
    .QN(_01704_),
    .RESETN(net476),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _34465_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_02662_),
    .QN(_01703_),
    .RESETN(net477),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34466_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_02663_),
    .QN(_01702_),
    .RESETN(net478),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34467_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_02664_),
    .QN(_01701_),
    .RESETN(net479),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _34468_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_02665_),
    .QN(_01700_),
    .RESETN(net480),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34469_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_02666_),
    .QN(_01699_),
    .RESETN(net481),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34470_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_02667_),
    .QN(_01698_),
    .RESETN(net482),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34471_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_02668_),
    .QN(_01697_),
    .RESETN(net483),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34472_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_02669_),
    .QN(_01696_),
    .RESETN(net484),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34473_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_02670_),
    .QN(_01695_),
    .RESETN(net485),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34474_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_02671_),
    .QN(_01694_),
    .RESETN(net486),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34475_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_02672_),
    .QN(_01693_),
    .RESETN(net487),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34476_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_02673_),
    .QN(_01692_),
    .RESETN(net488),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34477_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_02674_),
    .QN(_01691_),
    .RESETN(net489),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34478_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_02675_),
    .QN(_01690_),
    .RESETN(net490),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34479_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_02676_),
    .QN(_01689_),
    .RESETN(net491),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34480_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_02677_),
    .QN(_01688_),
    .RESETN(net492),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34481_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_02678_),
    .QN(_01687_),
    .RESETN(net493),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34482_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_02679_),
    .QN(_01686_),
    .RESETN(net494),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34483_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_02680_),
    .QN(_01685_),
    .RESETN(net495),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34484_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_02681_),
    .QN(_01684_),
    .RESETN(net496),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34485_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_02682_),
    .QN(_01683_),
    .RESETN(net497),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34486_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_02683_),
    .QN(_01682_),
    .RESETN(net498),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34487_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_02684_),
    .QN(_01681_),
    .RESETN(net499),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34488_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02685_),
    .QN(_01680_),
    .RESETN(net500),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34489_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_02686_),
    .QN(_01679_),
    .RESETN(net501),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34490_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_02687_),
    .QN(_01678_),
    .RESETN(net502),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34491_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02688_),
    .QN(_00324_),
    .RESETN(net503),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34492_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02689_),
    .QN(_00291_),
    .RESETN(net504),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34493_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02690_),
    .QN(_00663_),
    .RESETN(net505),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34494_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02691_),
    .QN(_00665_),
    .RESETN(net506),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34495_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02692_),
    .QN(_00668_),
    .RESETN(net507),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34496_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02693_),
    .QN(_00670_),
    .RESETN(net508),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34497_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02694_),
    .QN(_00672_),
    .RESETN(net509),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34498_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02695_),
    .QN(_00674_),
    .RESETN(net510),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34499_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02696_),
    .QN(_00677_),
    .RESETN(net511),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34500_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02697_),
    .QN(_00680_),
    .RESETN(net512),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34501_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02698_),
    .QN(_00682_),
    .RESETN(net513),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34502_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02699_),
    .QN(_00684_),
    .RESETN(net514),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34503_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02700_),
    .QN(_00686_),
    .RESETN(net515),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34504_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02701_),
    .QN(_00718_),
    .RESETN(net516),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34505_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02702_),
    .QN(_00750_),
    .RESETN(net517),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34506_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02703_),
    .QN(_00783_),
    .RESETN(net518),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34507_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02704_),
    .QN(_00816_),
    .RESETN(net519),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34508_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02705_),
    .QN(_00849_),
    .RESETN(net520),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34509_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02706_),
    .QN(_00881_),
    .RESETN(net521),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34510_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02707_),
    .QN(_00914_),
    .RESETN(net522),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34511_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02708_),
    .QN(_00946_),
    .RESETN(net523),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34512_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02709_),
    .QN(_00979_),
    .RESETN(net524),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34513_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02710_),
    .QN(_01011_),
    .RESETN(net525),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34514_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02711_),
    .QN(_01045_),
    .RESETN(net526),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34515_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02712_),
    .QN(_01077_),
    .RESETN(net527),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34516_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02713_),
    .QN(_01110_),
    .RESETN(net528),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34517_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02714_),
    .QN(_01142_),
    .RESETN(net529),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34518_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02715_),
    .QN(_01176_),
    .RESETN(net530),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34519_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02716_),
    .QN(_01208_),
    .RESETN(net531),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34520_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02717_),
    .QN(_01242_),
    .RESETN(net532),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34521_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02718_),
    .QN(_01274_),
    .RESETN(net533),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34522_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02719_),
    .QN(_01308_),
    .RESETN(net534),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34523_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02720_),
    .QN(_01677_),
    .RESETN(net535),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34524_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02721_),
    .QN(_00034_),
    .RESETN(net536),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34525_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_00002_),
    .QN(_01727_),
    .RESETN(net537),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34526_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_00003_),
    .QN(_01728_),
    .RESETN(net538),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34527_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_00004_),
    .QN(_00284_),
    .RESETN(net539),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34528_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_00005_),
    .QN(_01357_),
    .RESETN(net540),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34529_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02722_),
    .QN(_01676_),
    .RESETN(net541),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _34530_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02723_),
    .QN(_01675_),
    .RESETN(net542),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34531_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02724_),
    .QN(_01674_),
    .RESETN(net543),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _34532_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02725_),
    .QN(_01673_),
    .RESETN(net544),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _34533_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02726_),
    .QN(_01672_),
    .RESETN(net545),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34534_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02727_),
    .QN(_01671_),
    .RESETN(net546),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34535_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02728_),
    .QN(_01670_),
    .RESETN(net547),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34536_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02729_),
    .QN(_01669_),
    .RESETN(net548),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34537_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02730_),
    .QN(_01668_),
    .RESETN(net549),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34538_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02731_),
    .QN(_01667_),
    .RESETN(net550),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34539_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02732_),
    .QN(_01666_),
    .RESETN(net551),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34540_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02733_),
    .QN(_01665_),
    .RESETN(net552),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34541_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02734_),
    .QN(_01664_),
    .RESETN(net553),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34542_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02735_),
    .QN(_01663_),
    .RESETN(net554),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34543_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02736_),
    .QN(_01662_),
    .RESETN(net555),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34544_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02737_),
    .QN(_01661_),
    .RESETN(net556),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34545_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02738_),
    .QN(_01660_),
    .RESETN(net557),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34546_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02739_),
    .QN(_01659_),
    .RESETN(net558),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _34547_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02740_),
    .QN(_01658_),
    .RESETN(net559),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34548_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02741_),
    .QN(_01657_),
    .RESETN(net560),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34549_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02742_),
    .QN(_01656_),
    .RESETN(net561),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34550_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02743_),
    .QN(_01655_),
    .RESETN(net562),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34551_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02744_),
    .QN(_01654_),
    .RESETN(net563),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34552_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02745_),
    .QN(_01653_),
    .RESETN(net564),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34553_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02746_),
    .QN(_01652_),
    .RESETN(net565),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34554_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02747_),
    .QN(_01651_),
    .RESETN(net566),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34555_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02748_),
    .QN(_01650_),
    .RESETN(net567),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34556_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02749_),
    .QN(_01649_),
    .RESETN(net568),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34557_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02750_),
    .QN(_01648_),
    .RESETN(net569),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34558_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02751_),
    .QN(_01647_),
    .RESETN(net570),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34559_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02752_),
    .QN(_01646_),
    .RESETN(net571),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34560_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02753_),
    .QN(_01645_),
    .RESETN(net572),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34561_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02754_),
    .QN(_01323_),
    .RESETN(net573),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34562_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02755_),
    .QN(_01324_),
    .RESETN(net574),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34563_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02756_),
    .QN(_01325_),
    .RESETN(net575),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34564_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02757_),
    .QN(_01327_),
    .RESETN(net576),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34565_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02758_),
    .QN(_01328_),
    .RESETN(net577),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34566_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02759_),
    .QN(_01329_),
    .RESETN(net578),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34567_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02760_),
    .QN(_01330_),
    .RESETN(net579),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34568_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02761_),
    .QN(_01331_),
    .RESETN(net580),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34569_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02762_),
    .QN(_01332_),
    .RESETN(net581),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34570_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02763_),
    .QN(_01333_),
    .RESETN(net582),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34571_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02764_),
    .QN(_01334_),
    .RESETN(net583),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34572_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02765_),
    .QN(_01335_),
    .RESETN(net584),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34573_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02766_),
    .QN(_01336_),
    .RESETN(net585),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34574_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02767_),
    .QN(_01337_),
    .RESETN(net586),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34575_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02768_),
    .QN(_01338_),
    .RESETN(net587),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34576_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02769_),
    .QN(_01339_),
    .RESETN(net588),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34577_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02770_),
    .QN(_01340_),
    .RESETN(net589),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34578_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02771_),
    .QN(_01341_),
    .RESETN(net590),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34579_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02772_),
    .QN(_01342_),
    .RESETN(net591),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34580_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02773_),
    .QN(_01343_),
    .RESETN(net592),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34581_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02774_),
    .QN(_01344_),
    .RESETN(net593),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34582_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02775_),
    .QN(_01345_),
    .RESETN(net594),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34583_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02776_),
    .QN(_01346_),
    .RESETN(net595),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34584_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02777_),
    .QN(_01347_),
    .RESETN(net596),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34585_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02778_),
    .QN(_01348_),
    .RESETN(net597),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34586_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02779_),
    .QN(_01349_),
    .RESETN(net598),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34587_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02780_),
    .QN(_01350_),
    .RESETN(net599),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34588_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02781_),
    .QN(_01351_),
    .RESETN(net600),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34589_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_02782_),
    .QN(_01352_),
    .RESETN(net601),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34590_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02783_),
    .QN(_01353_),
    .RESETN(net602),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34591_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02784_),
    .QN(_01354_),
    .RESETN(net603),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34592_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02785_),
    .QN(_01355_),
    .RESETN(net604),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34593_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02786_),
    .QN(_17600_),
    .RESETN(net605),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34594_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02787_),
    .QN(_17601_),
    .RESETN(net606),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34595_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02788_),
    .QN(_17607_),
    .RESETN(net607),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34596_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02789_),
    .QN(_01322_),
    .RESETN(net608),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34597_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_02790_),
    .QN(_01318_),
    .RESETN(net609),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34598_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02791_),
    .QN(_01316_),
    .RESETN(net610),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34599_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02792_),
    .QN(_01644_),
    .RESETN(net611),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34600_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02793_),
    .QN(_01643_),
    .RESETN(net612),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34601_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02794_),
    .QN(_01642_),
    .RESETN(net613),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34602_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02795_),
    .QN(_01641_),
    .RESETN(net614),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34603_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02796_),
    .QN(_01640_),
    .RESETN(net615),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34604_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02797_),
    .QN(_01639_),
    .RESETN(net616),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34605_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02798_),
    .QN(_01638_),
    .RESETN(net617),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34606_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02799_),
    .QN(_01637_),
    .RESETN(net618),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34607_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02800_),
    .QN(_01636_),
    .RESETN(net619),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34608_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02801_),
    .QN(_01635_),
    .RESETN(net620),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34609_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02802_),
    .QN(_01634_),
    .RESETN(net621),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _34610_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02803_),
    .QN(_01633_),
    .RESETN(net622),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _34611_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02804_),
    .QN(_01632_),
    .RESETN(net623),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34612_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02805_),
    .QN(_01631_),
    .RESETN(net624),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _34613_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02806_),
    .QN(_01630_),
    .RESETN(net625),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _34614_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02807_),
    .QN(_01629_),
    .RESETN(net626),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34615_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02808_),
    .QN(_01628_),
    .RESETN(net627),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34616_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02809_),
    .QN(_01627_),
    .RESETN(net628),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34617_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02810_),
    .QN(_01626_),
    .RESETN(net629),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _34618_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02811_),
    .QN(_01625_),
    .RESETN(net630),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _34619_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02812_),
    .QN(_01624_),
    .RESETN(net631),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34620_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02813_),
    .QN(_01623_),
    .RESETN(net632),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34621_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02814_),
    .QN(_01622_),
    .RESETN(net633),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34622_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02815_),
    .QN(_01621_),
    .RESETN(net634),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34623_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02816_),
    .QN(_01620_),
    .RESETN(net635),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34624_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02817_),
    .QN(_01619_),
    .RESETN(net636),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _34625_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02818_),
    .QN(_01618_),
    .RESETN(net637),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34626_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02819_),
    .QN(_01617_),
    .RESETN(net638),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34627_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02820_),
    .QN(_01616_),
    .RESETN(net639),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _34628_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02821_),
    .QN(_01615_),
    .RESETN(net640),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34629_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02822_),
    .QN(_01614_),
    .RESETN(net641),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _34630_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02823_),
    .QN(_01613_),
    .RESETN(net642),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _34631_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02824_),
    .QN(_01612_),
    .RESETN(net643),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34632_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02825_),
    .QN(_01611_),
    .RESETN(net644),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34633_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02826_),
    .QN(_01610_),
    .RESETN(net645),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34634_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02827_),
    .QN(_01609_),
    .RESETN(net646),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34635_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02828_),
    .QN(_01608_),
    .RESETN(net647),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34636_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02829_),
    .QN(_00277_),
    .RESETN(net648),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34637_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02830_),
    .QN(_01607_),
    .RESETN(net649),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34638_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02831_),
    .QN(_18336_),
    .RESETN(net650),
    .SETN(net433));
 DFFHQNx1_ASAP7_75t_R _34639_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02832_),
    .QN(_00662_));
 DFFHQNx1_ASAP7_75t_R _34640_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02833_),
    .QN(_17536_));
 DFFHQNx1_ASAP7_75t_R _34641_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02834_),
    .QN(_01606_));
 DFFHQNx1_ASAP7_75t_R _34642_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02835_),
    .QN(_01605_));
 DFFHQNx1_ASAP7_75t_R _34643_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02836_),
    .QN(_01604_));
 DFFHQNx1_ASAP7_75t_R _34644_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02837_),
    .QN(_01603_));
 DFFHQNx1_ASAP7_75t_R _34645_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02838_),
    .QN(_01602_));
 DFFHQNx1_ASAP7_75t_R _34646_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02839_),
    .QN(_01601_));
 DFFHQNx1_ASAP7_75t_R _34647_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02840_),
    .QN(_01600_));
 DFFHQNx1_ASAP7_75t_R _34648_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02841_),
    .QN(_01599_));
 DFFHQNx1_ASAP7_75t_R _34649_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02842_),
    .QN(_01598_));
 DFFHQNx1_ASAP7_75t_R _34650_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02843_),
    .QN(_01597_));
 DFFHQNx1_ASAP7_75t_R _34651_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02844_),
    .QN(_01596_));
 DFFHQNx1_ASAP7_75t_R _34652_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02845_),
    .QN(_01595_));
 DFFHQNx1_ASAP7_75t_R _34653_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02846_),
    .QN(_01594_));
 DFFHQNx1_ASAP7_75t_R _34654_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02847_),
    .QN(_01593_));
 DFFHQNx1_ASAP7_75t_R _34655_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02848_),
    .QN(_01592_));
 DFFHQNx1_ASAP7_75t_R _34656_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02849_),
    .QN(_01591_));
 DFFHQNx1_ASAP7_75t_R _34657_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02850_),
    .QN(_01590_));
 DFFHQNx1_ASAP7_75t_R _34658_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02851_),
    .QN(_01589_));
 DFFHQNx1_ASAP7_75t_R _34659_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02852_),
    .QN(_01588_));
 DFFHQNx1_ASAP7_75t_R _34660_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02853_),
    .QN(_01587_));
 DFFHQNx1_ASAP7_75t_R _34661_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02854_),
    .QN(_01586_));
 DFFHQNx1_ASAP7_75t_R _34662_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02855_),
    .QN(_01585_));
 DFFHQNx1_ASAP7_75t_R _34663_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02856_),
    .QN(_01584_));
 DFFHQNx1_ASAP7_75t_R _34664_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02857_),
    .QN(_01583_));
 DFFHQNx1_ASAP7_75t_R _34665_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02858_),
    .QN(_01582_));
 DFFHQNx1_ASAP7_75t_R _34666_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02859_),
    .QN(_01581_));
 DFFHQNx1_ASAP7_75t_R _34667_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02860_),
    .QN(_01580_));
 DFFHQNx1_ASAP7_75t_R _34668_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02861_),
    .QN(_01579_));
 DFFHQNx1_ASAP7_75t_R _34669_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02862_),
    .QN(_01578_));
 DFFASRHQNx1_ASAP7_75t_R _34670_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_02863_),
    .QN(_01577_),
    .RESETN(net449),
    .SETN(net651));
 DFFASRHQNx1_ASAP7_75t_R _34671_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_02864_),
    .QN(_01576_),
    .RESETN(net449),
    .SETN(net652));
 DFFASRHQNx1_ASAP7_75t_R _34672_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02865_),
    .QN(_00658_),
    .RESETN(net653),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34673_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02866_),
    .QN(_01575_),
    .RESETN(net654),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34674_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02867_),
    .QN(_00081_),
    .RESETN(net655),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34675_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_02868_),
    .QN(_00084_),
    .RESETN(net656),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34676_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_02869_),
    .QN(_00087_),
    .RESETN(net657),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34677_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02870_),
    .QN(_00090_),
    .RESETN(net658),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _34678_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02871_),
    .QN(_01574_),
    .RESETN(net659),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _34679_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02872_),
    .QN(_01573_),
    .RESETN(net660),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _34680_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02873_),
    .QN(_01572_),
    .RESETN(net661),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _34681_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02874_),
    .QN(_01571_),
    .RESETN(net662),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _34682_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02875_),
    .QN(_01570_),
    .RESETN(net663),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34683_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02876_),
    .QN(_01569_),
    .RESETN(net664),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _34684_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_02877_),
    .QN(_01568_),
    .RESETN(net665),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _34685_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02878_),
    .QN(_01567_),
    .RESETN(net666),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34686_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02879_),
    .QN(_01566_),
    .RESETN(net667),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34687_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02880_),
    .QN(_01565_),
    .RESETN(net668),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _34688_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_02881_),
    .QN(_01564_),
    .RESETN(net669),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _34689_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02882_),
    .QN(_01563_),
    .RESETN(net670),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _34690_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02883_),
    .QN(_01562_),
    .RESETN(net671),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34691_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02884_),
    .QN(_01561_),
    .RESETN(net672),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _34692_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_02885_),
    .QN(_01560_),
    .RESETN(net673),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34693_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02886_),
    .QN(_01559_),
    .RESETN(net674),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _34694_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_02887_),
    .QN(_01558_),
    .RESETN(net675),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _34695_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_02888_),
    .QN(_01557_),
    .RESETN(net676),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _34696_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_02889_),
    .QN(_01556_),
    .RESETN(net677),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34697_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02890_),
    .QN(_01555_),
    .RESETN(net678),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34698_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_02891_),
    .QN(_01554_),
    .RESETN(net679),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34699_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02892_),
    .QN(_01553_),
    .RESETN(net680),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _34700_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_02893_),
    .QN(_01552_),
    .RESETN(net681),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _34701_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02894_),
    .QN(_01551_),
    .RESETN(net682),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _34702_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02895_),
    .QN(_01550_),
    .RESETN(net683),
    .SETN(net434));
 DFFHQNx1_ASAP7_75t_R _34703_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_02896_),
    .QN(_01549_));
 DFFHQNx1_ASAP7_75t_R _34704_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_02897_),
    .QN(_01548_));
 DFFHQNx1_ASAP7_75t_R _34705_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02898_),
    .QN(_01547_));
 DFFHQNx1_ASAP7_75t_R _34706_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_02899_),
    .QN(_01546_));
 DFFHQNx1_ASAP7_75t_R _34707_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_02900_),
    .QN(_01545_));
 DFFHQNx1_ASAP7_75t_R _34708_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02901_),
    .QN(_01544_));
 DFFHQNx1_ASAP7_75t_R _34709_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02902_),
    .QN(_01543_));
 DFFHQNx1_ASAP7_75t_R _34710_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02903_),
    .QN(_01542_));
 DFFHQNx1_ASAP7_75t_R _34711_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02904_),
    .QN(_01541_));
 DFFHQNx1_ASAP7_75t_R _34712_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02905_),
    .QN(_01540_));
 DFFHQNx1_ASAP7_75t_R _34713_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02906_),
    .QN(_01539_));
 DFFHQNx1_ASAP7_75t_R _34714_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02907_),
    .QN(_01538_));
 DFFHQNx1_ASAP7_75t_R _34715_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02908_),
    .QN(_01537_));
 DFFHQNx1_ASAP7_75t_R _34716_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02909_),
    .QN(_01536_));
 DFFHQNx1_ASAP7_75t_R _34717_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02910_),
    .QN(_01535_));
 DFFHQNx1_ASAP7_75t_R _34718_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02911_),
    .QN(_01534_));
 DFFHQNx1_ASAP7_75t_R _34719_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02912_),
    .QN(_01533_));
 DFFHQNx1_ASAP7_75t_R _34720_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02913_),
    .QN(_01532_));
 DFFHQNx1_ASAP7_75t_R _34721_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02914_),
    .QN(_01531_));
 DFFHQNx1_ASAP7_75t_R _34722_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02915_),
    .QN(_01530_));
 DFFHQNx1_ASAP7_75t_R _34723_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02916_),
    .QN(_01529_));
 DFFHQNx1_ASAP7_75t_R _34724_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02917_),
    .QN(_01528_));
 DFFHQNx1_ASAP7_75t_R _34725_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02918_),
    .QN(_01527_));
 DFFHQNx1_ASAP7_75t_R _34726_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02919_),
    .QN(_01526_));
 DFFHQNx1_ASAP7_75t_R _34727_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02920_),
    .QN(_01525_));
 DFFHQNx1_ASAP7_75t_R _34728_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02921_),
    .QN(_01524_));
 DFFHQNx1_ASAP7_75t_R _34729_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02922_),
    .QN(_01523_));
 DFFHQNx1_ASAP7_75t_R _34730_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02923_),
    .QN(_01522_));
 DFFHQNx1_ASAP7_75t_R _34731_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02924_),
    .QN(_01521_));
 DFFHQNx1_ASAP7_75t_R _34732_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02925_),
    .QN(_01520_));
 DFFASRHQNx1_ASAP7_75t_R _34733_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_02926_),
    .QN(_00293_),
    .RESETN(net684),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34734_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_02927_),
    .QN(_00247_),
    .RESETN(net685),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34735_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_02928_),
    .QN(_00355_),
    .RESETN(net686),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _34736_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_02929_),
    .QN(_00386_),
    .RESETN(net687),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34737_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_02930_),
    .QN(_00416_),
    .RESETN(net688),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34738_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_02931_),
    .QN(_00446_),
    .RESETN(net689),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _34739_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_02932_),
    .QN(_00476_),
    .RESETN(net690),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34740_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_02933_),
    .QN(_00506_),
    .RESETN(net691),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34741_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_02934_),
    .QN(_00536_),
    .RESETN(net692),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _34742_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_02935_),
    .QN(_00566_),
    .RESETN(net693),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _34743_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_02936_),
    .QN(_00596_),
    .RESETN(net694),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34744_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_02937_),
    .QN(_00626_),
    .RESETN(net695),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _34745_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_02938_),
    .QN(_00325_),
    .RESETN(net696),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34746_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_02939_),
    .QN(_00688_),
    .RESETN(net697),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34747_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_02940_),
    .QN(_00720_),
    .RESETN(net698),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _34748_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_02941_),
    .QN(_00753_),
    .RESETN(net699),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34749_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02942_),
    .QN(_00786_),
    .RESETN(net700),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34750_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_02943_),
    .QN(_00819_),
    .RESETN(net701),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34751_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_02944_),
    .QN(_00851_),
    .RESETN(net702),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34752_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_02945_),
    .QN(_00884_),
    .RESETN(net703),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34753_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_02946_),
    .QN(_00916_),
    .RESETN(net704),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34754_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_02947_),
    .QN(_00949_),
    .RESETN(net705),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _34755_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_02948_),
    .QN(_00981_),
    .RESETN(net706),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _34756_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_02949_),
    .QN(_01015_),
    .RESETN(net707),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34757_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02950_),
    .QN(_01047_),
    .RESETN(net708),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34758_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_02951_),
    .QN(_01080_),
    .RESETN(net709),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34759_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_02952_),
    .QN(_01112_),
    .RESETN(net710),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34760_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02953_),
    .QN(_01146_),
    .RESETN(net711),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34761_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_02954_),
    .QN(_01178_),
    .RESETN(net712),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _34762_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02955_),
    .QN(_01212_),
    .RESETN(net713),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34763_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_02956_),
    .QN(_01244_),
    .RESETN(net714),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34764_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_02957_),
    .QN(_01278_),
    .RESETN(net715),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34765_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_02958_),
    .QN(_00294_),
    .RESETN(net716),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34766_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_02959_),
    .QN(_00248_),
    .RESETN(net717),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34767_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_02960_),
    .QN(_00356_),
    .RESETN(net718),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _34768_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_02961_),
    .QN(_00387_),
    .RESETN(net719),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34769_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_02962_),
    .QN(_00417_),
    .RESETN(net720),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _34770_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_02963_),
    .QN(_00447_),
    .RESETN(net721),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34771_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_02964_),
    .QN(_00477_),
    .RESETN(net722),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34772_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_02965_),
    .QN(_00507_),
    .RESETN(net723),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34773_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_02966_),
    .QN(_00537_),
    .RESETN(net724),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34774_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_02967_),
    .QN(_00567_),
    .RESETN(net725),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34775_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_02968_),
    .QN(_00597_),
    .RESETN(net726),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34776_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_02969_),
    .QN(_00627_),
    .RESETN(net727),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34777_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_02970_),
    .QN(_00326_),
    .RESETN(net728),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34778_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_02971_),
    .QN(_00689_),
    .RESETN(net729),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34779_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_02972_),
    .QN(_00721_),
    .RESETN(net730),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _34780_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_02973_),
    .QN(_00754_),
    .RESETN(net731),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34781_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_02974_),
    .QN(_00787_),
    .RESETN(net732),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34782_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_02975_),
    .QN(_00820_),
    .RESETN(net733),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34783_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_02976_),
    .QN(_00852_),
    .RESETN(net734),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34784_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_02977_),
    .QN(_00885_),
    .RESETN(net735),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34785_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_02978_),
    .QN(_00917_),
    .RESETN(net736),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34786_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_02979_),
    .QN(_00950_),
    .RESETN(net737),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34787_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_02980_),
    .QN(_00982_),
    .RESETN(net738),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34788_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_02981_),
    .QN(_01016_),
    .RESETN(net739),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34789_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_02982_),
    .QN(_01048_),
    .RESETN(net740),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34790_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_02983_),
    .QN(_01081_),
    .RESETN(net741),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34791_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_02984_),
    .QN(_01113_),
    .RESETN(net742),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34792_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_02985_),
    .QN(_01147_),
    .RESETN(net743),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34793_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_02986_),
    .QN(_01179_),
    .RESETN(net744),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34794_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02987_),
    .QN(_01213_),
    .RESETN(net745),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34795_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_02988_),
    .QN(_01245_),
    .RESETN(net746),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34796_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_02989_),
    .QN(_01279_),
    .RESETN(net747),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34797_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_02990_),
    .QN(_00295_),
    .RESETN(net748),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34798_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_02991_),
    .QN(_00249_),
    .RESETN(net749),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34799_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_02992_),
    .QN(_00357_),
    .RESETN(net750),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34800_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_02993_),
    .QN(_00388_),
    .RESETN(net751),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34801_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_02994_),
    .QN(_00418_),
    .RESETN(net752),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34802_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_02995_),
    .QN(_00448_),
    .RESETN(net753),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34803_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_02996_),
    .QN(_00478_),
    .RESETN(net754),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34804_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_02997_),
    .QN(_00508_),
    .RESETN(net755),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34805_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_02998_),
    .QN(_00538_),
    .RESETN(net756),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _34806_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_02999_),
    .QN(_00568_),
    .RESETN(net757),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _34807_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03000_),
    .QN(_00598_),
    .RESETN(net758),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34808_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03001_),
    .QN(_00628_),
    .RESETN(net759),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34809_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03002_),
    .QN(_00327_),
    .RESETN(net760),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34810_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03003_),
    .QN(_00690_),
    .RESETN(net761),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34811_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03004_),
    .QN(_00722_),
    .RESETN(net762),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34812_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03005_),
    .QN(_00755_),
    .RESETN(net763),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34813_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03006_),
    .QN(_00788_),
    .RESETN(net764),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34814_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03007_),
    .QN(_00821_),
    .RESETN(net765),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34815_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03008_),
    .QN(_00853_),
    .RESETN(net766),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34816_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03009_),
    .QN(_00886_),
    .RESETN(net767),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _34817_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03010_),
    .QN(_00918_),
    .RESETN(net768),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34818_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03011_),
    .QN(_00951_),
    .RESETN(net769),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _34819_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03012_),
    .QN(_00983_),
    .RESETN(net770),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34820_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03013_),
    .QN(_01017_),
    .RESETN(net771),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34821_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03014_),
    .QN(_01049_),
    .RESETN(net772),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34822_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03015_),
    .QN(_01082_),
    .RESETN(net773),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34823_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03016_),
    .QN(_01114_),
    .RESETN(net774),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34824_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03017_),
    .QN(_01148_),
    .RESETN(net775),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34825_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03018_),
    .QN(_01180_),
    .RESETN(net776),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34826_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03019_),
    .QN(_01214_),
    .RESETN(net777),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34827_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03020_),
    .QN(_01246_),
    .RESETN(net778),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34828_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03021_),
    .QN(_01280_),
    .RESETN(net779),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34829_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03022_),
    .QN(_00296_),
    .RESETN(net780),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _34830_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03023_),
    .QN(_00250_),
    .RESETN(net781),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34831_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03024_),
    .QN(_00358_),
    .RESETN(net782),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34832_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03025_),
    .QN(_00389_),
    .RESETN(net783),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34833_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03026_),
    .QN(_00419_),
    .RESETN(net784),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34834_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03027_),
    .QN(_00449_),
    .RESETN(net785),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34835_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03028_),
    .QN(_00479_),
    .RESETN(net786),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34836_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03029_),
    .QN(_00509_),
    .RESETN(net787),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34837_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03030_),
    .QN(_00539_),
    .RESETN(net788),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _34838_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03031_),
    .QN(_00569_),
    .RESETN(net789),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _34839_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03032_),
    .QN(_00599_),
    .RESETN(net790),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34840_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03033_),
    .QN(_00629_),
    .RESETN(net791),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _34841_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03034_),
    .QN(_00328_),
    .RESETN(net792),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34842_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03035_),
    .QN(_00691_),
    .RESETN(net793),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34843_ (.CLK(clknet_level_3_1_34135_clk_i),
    .D(_03036_),
    .QN(_00723_),
    .RESETN(net794),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34844_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03037_),
    .QN(_00756_),
    .RESETN(net795),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34845_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03038_),
    .QN(_00789_),
    .RESETN(net796),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34846_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03039_),
    .QN(_00822_),
    .RESETN(net797),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34847_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03040_),
    .QN(_00854_),
    .RESETN(net798),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34848_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03041_),
    .QN(_00887_),
    .RESETN(net799),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34849_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03042_),
    .QN(_00919_),
    .RESETN(net800),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34850_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03043_),
    .QN(_00952_),
    .RESETN(net801),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _34851_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03044_),
    .QN(_00984_),
    .RESETN(net802),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34852_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03045_),
    .QN(_01018_),
    .RESETN(net803),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34853_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03046_),
    .QN(_01050_),
    .RESETN(net804),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34854_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03047_),
    .QN(_01083_),
    .RESETN(net805),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34855_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03048_),
    .QN(_01115_),
    .RESETN(net806),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34856_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03049_),
    .QN(_01149_),
    .RESETN(net807),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34857_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03050_),
    .QN(_01181_),
    .RESETN(net808),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34858_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03051_),
    .QN(_01215_),
    .RESETN(net809),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34859_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03052_),
    .QN(_01247_),
    .RESETN(net810),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34860_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03053_),
    .QN(_01281_),
    .RESETN(net811),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34861_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03054_),
    .QN(_00297_),
    .RESETN(net812),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34862_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03055_),
    .QN(_00251_),
    .RESETN(net813),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34863_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03056_),
    .QN(_00359_),
    .RESETN(net814),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34864_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03057_),
    .QN(_00390_),
    .RESETN(net815),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34865_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03058_),
    .QN(_00420_),
    .RESETN(net816),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34866_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03059_),
    .QN(_00450_),
    .RESETN(net817),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34867_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03060_),
    .QN(_00480_),
    .RESETN(net818),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34868_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03061_),
    .QN(_00510_),
    .RESETN(net819),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34869_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03062_),
    .QN(_00540_),
    .RESETN(net820),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _34870_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03063_),
    .QN(_00570_),
    .RESETN(net821),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34871_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03064_),
    .QN(_00600_),
    .RESETN(net822),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34872_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03065_),
    .QN(_00630_),
    .RESETN(net823),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34873_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03066_),
    .QN(_00329_),
    .RESETN(net824),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34874_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03067_),
    .QN(_00692_),
    .RESETN(net825),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34875_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03068_),
    .QN(_00724_),
    .RESETN(net826),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34876_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03069_),
    .QN(_00757_),
    .RESETN(net827),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34877_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03070_),
    .QN(_00790_),
    .RESETN(net828),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34878_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03071_),
    .QN(_00823_),
    .RESETN(net829),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34879_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03072_),
    .QN(_00855_),
    .RESETN(net830),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34880_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03073_),
    .QN(_00888_),
    .RESETN(net831),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34881_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03074_),
    .QN(_00920_),
    .RESETN(net832),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34882_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03075_),
    .QN(_00953_),
    .RESETN(net833),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _34883_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03076_),
    .QN(_00985_),
    .RESETN(net834),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34884_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03077_),
    .QN(_01019_),
    .RESETN(net835),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34885_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03078_),
    .QN(_01051_),
    .RESETN(net836),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34886_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03079_),
    .QN(_01084_),
    .RESETN(net837),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34887_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03080_),
    .QN(_01116_),
    .RESETN(net838),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34888_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03081_),
    .QN(_01150_),
    .RESETN(net839),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34889_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03082_),
    .QN(_01182_),
    .RESETN(net840),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34890_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03083_),
    .QN(_01216_),
    .RESETN(net841),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34891_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03084_),
    .QN(_01248_),
    .RESETN(net842),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34892_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03085_),
    .QN(_01282_),
    .RESETN(net843),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34893_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03086_),
    .QN(_00298_),
    .RESETN(net844),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34894_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03087_),
    .QN(_00252_),
    .RESETN(net845),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34895_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03088_),
    .QN(_00360_),
    .RESETN(net846),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _34896_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03089_),
    .QN(_00391_),
    .RESETN(net847),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34897_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03090_),
    .QN(_00421_),
    .RESETN(net848),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34898_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03091_),
    .QN(_00451_),
    .RESETN(net849),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34899_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03092_),
    .QN(_00481_),
    .RESETN(net850),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34900_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03093_),
    .QN(_00511_),
    .RESETN(net851),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34901_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03094_),
    .QN(_00541_),
    .RESETN(net852),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _34902_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03095_),
    .QN(_00571_),
    .RESETN(net853),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34903_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03096_),
    .QN(_00601_),
    .RESETN(net854),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34904_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03097_),
    .QN(_00631_),
    .RESETN(net855),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34905_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03098_),
    .QN(_00330_),
    .RESETN(net856),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34906_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03099_),
    .QN(_00693_),
    .RESETN(net857),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34907_ (.CLK(clknet_level_3_1_34135_clk_i),
    .D(_03100_),
    .QN(_00725_),
    .RESETN(net858),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34908_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03101_),
    .QN(_00758_),
    .RESETN(net859),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34909_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03102_),
    .QN(_00791_),
    .RESETN(net860),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34910_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03103_),
    .QN(_00824_),
    .RESETN(net861),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34911_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03104_),
    .QN(_00856_),
    .RESETN(net862),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34912_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03105_),
    .QN(_00889_),
    .RESETN(net863),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34913_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03106_),
    .QN(_00921_),
    .RESETN(net864),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34914_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03107_),
    .QN(_00954_),
    .RESETN(net865),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _34915_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03108_),
    .QN(_00986_),
    .RESETN(net866),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34916_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03109_),
    .QN(_01020_),
    .RESETN(net867),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34917_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03110_),
    .QN(_01052_),
    .RESETN(net868),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34918_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03111_),
    .QN(_01085_),
    .RESETN(net869),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34919_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03112_),
    .QN(_01117_),
    .RESETN(net870),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34920_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03113_),
    .QN(_01151_),
    .RESETN(net871),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34921_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03114_),
    .QN(_01183_),
    .RESETN(net872),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34922_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03115_),
    .QN(_01217_),
    .RESETN(net873),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34923_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03116_),
    .QN(_01249_),
    .RESETN(net874),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34924_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03117_),
    .QN(_01283_),
    .RESETN(net875),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34925_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03118_),
    .QN(_00299_),
    .RESETN(net876),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _34926_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03119_),
    .QN(_00253_),
    .RESETN(net877),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34927_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03120_),
    .QN(_00361_),
    .RESETN(net878),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _34928_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03121_),
    .QN(_00392_),
    .RESETN(net879),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34929_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03122_),
    .QN(_00422_),
    .RESETN(net880),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34930_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03123_),
    .QN(_00452_),
    .RESETN(net881),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _34931_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03124_),
    .QN(_00482_),
    .RESETN(net882),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34932_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03125_),
    .QN(_00512_),
    .RESETN(net883),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34933_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03126_),
    .QN(_00542_),
    .RESETN(net884),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34934_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03127_),
    .QN(_00572_),
    .RESETN(net885),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34935_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03128_),
    .QN(_00602_),
    .RESETN(net886),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34936_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03129_),
    .QN(_00632_),
    .RESETN(net887),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34937_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03130_),
    .QN(_00331_),
    .RESETN(net888),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34938_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03131_),
    .QN(_00694_),
    .RESETN(net889),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34939_ (.CLK(clknet_level_3_1_34135_clk_i),
    .D(_03132_),
    .QN(_00726_),
    .RESETN(net890),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34940_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03133_),
    .QN(_00759_),
    .RESETN(net891),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34941_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03134_),
    .QN(_00792_),
    .RESETN(net892),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34942_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03135_),
    .QN(_00825_),
    .RESETN(net893),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34943_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03136_),
    .QN(_00857_),
    .RESETN(net894),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34944_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03137_),
    .QN(_00890_),
    .RESETN(net895),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34945_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03138_),
    .QN(_00922_),
    .RESETN(net896),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34946_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03139_),
    .QN(_00955_),
    .RESETN(net897),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _34947_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03140_),
    .QN(_00987_),
    .RESETN(net898),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34948_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03141_),
    .QN(_01021_),
    .RESETN(net899),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34949_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03142_),
    .QN(_01053_),
    .RESETN(net900),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34950_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03143_),
    .QN(_01086_),
    .RESETN(net901),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34951_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03144_),
    .QN(_01118_),
    .RESETN(net902),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34952_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03145_),
    .QN(_01152_),
    .RESETN(net903),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34953_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03146_),
    .QN(_01184_),
    .RESETN(net904),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34954_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03147_),
    .QN(_01218_),
    .RESETN(net905),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34955_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03148_),
    .QN(_01250_),
    .RESETN(net906),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34956_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03149_),
    .QN(_01284_),
    .RESETN(net907),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34957_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03150_),
    .QN(_00300_),
    .RESETN(net908),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _34958_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03151_),
    .QN(_00254_),
    .RESETN(net909),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34959_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03152_),
    .QN(_00362_),
    .RESETN(net910),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _34960_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03153_),
    .QN(_00393_),
    .RESETN(net911),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34961_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03154_),
    .QN(_00423_),
    .RESETN(net912),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34962_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03155_),
    .QN(_00453_),
    .RESETN(net913),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _34963_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03156_),
    .QN(_00483_),
    .RESETN(net914),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _34964_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03157_),
    .QN(_00513_),
    .RESETN(net915),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34965_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03158_),
    .QN(_00543_),
    .RESETN(net916),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34966_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03159_),
    .QN(_00573_),
    .RESETN(net917),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34967_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03160_),
    .QN(_00603_),
    .RESETN(net918),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34968_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03161_),
    .QN(_00633_),
    .RESETN(net919),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34969_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03162_),
    .QN(_00332_),
    .RESETN(net920),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _34970_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03163_),
    .QN(_00695_),
    .RESETN(net921),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34971_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03164_),
    .QN(_00727_),
    .RESETN(net922),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _34972_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03165_),
    .QN(_00760_),
    .RESETN(net923),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34973_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03166_),
    .QN(_00793_),
    .RESETN(net924),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _34974_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03167_),
    .QN(_00826_),
    .RESETN(net925),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _34975_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03168_),
    .QN(_00858_),
    .RESETN(net926),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34976_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03169_),
    .QN(_00891_),
    .RESETN(net927),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _34977_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03170_),
    .QN(_00923_),
    .RESETN(net928),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34978_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03171_),
    .QN(_00956_),
    .RESETN(net929),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _34979_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03172_),
    .QN(_00988_),
    .RESETN(net930),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34980_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03173_),
    .QN(_01022_),
    .RESETN(net931),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34981_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03174_),
    .QN(_01054_),
    .RESETN(net932),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34982_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03175_),
    .QN(_01087_),
    .RESETN(net933),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34983_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03176_),
    .QN(_01119_),
    .RESETN(net934),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34984_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03177_),
    .QN(_01153_),
    .RESETN(net935),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34985_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03178_),
    .QN(_01185_),
    .RESETN(net936),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _34986_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03179_),
    .QN(_01219_),
    .RESETN(net937),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34987_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03180_),
    .QN(_01251_),
    .RESETN(net938),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _34988_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03181_),
    .QN(_01285_),
    .RESETN(net939),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34989_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03182_),
    .QN(_00301_),
    .RESETN(net940),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _34990_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03183_),
    .QN(_00255_),
    .RESETN(net941),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34991_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03184_),
    .QN(_00363_),
    .RESETN(net942),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _34992_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03185_),
    .QN(_00394_),
    .RESETN(net943),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _34993_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03186_),
    .QN(_00424_),
    .RESETN(net944),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34994_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03187_),
    .QN(_00454_),
    .RESETN(net945),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _34995_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03188_),
    .QN(_00484_),
    .RESETN(net946),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _34996_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03189_),
    .QN(_00514_),
    .RESETN(net947),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _34997_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03190_),
    .QN(_00544_),
    .RESETN(net948),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _34998_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03191_),
    .QN(_00574_),
    .RESETN(net949),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _34999_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03192_),
    .QN(_00604_),
    .RESETN(net950),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35000_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03193_),
    .QN(_00634_),
    .RESETN(net951),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35001_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03194_),
    .QN(_00333_),
    .RESETN(net952),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35002_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03195_),
    .QN(_00696_),
    .RESETN(net953),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35003_ (.CLK(clknet_level_3_1_34135_clk_i),
    .D(_03196_),
    .QN(_00728_),
    .RESETN(net954),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35004_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03197_),
    .QN(_00761_),
    .RESETN(net955),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35005_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03198_),
    .QN(_00794_),
    .RESETN(net956),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35006_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03199_),
    .QN(_00827_),
    .RESETN(net957),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35007_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03200_),
    .QN(_00859_),
    .RESETN(net958),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35008_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03201_),
    .QN(_00892_),
    .RESETN(net959),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35009_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03202_),
    .QN(_00924_),
    .RESETN(net960),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35010_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03203_),
    .QN(_00957_),
    .RESETN(net961),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35011_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03204_),
    .QN(_00989_),
    .RESETN(net962),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35012_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03205_),
    .QN(_01023_),
    .RESETN(net963),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35013_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03206_),
    .QN(_01055_),
    .RESETN(net964),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35014_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03207_),
    .QN(_01088_),
    .RESETN(net965),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35015_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03208_),
    .QN(_01120_),
    .RESETN(net966),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35016_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03209_),
    .QN(_01154_),
    .RESETN(net967),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35017_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03210_),
    .QN(_01186_),
    .RESETN(net968),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35018_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03211_),
    .QN(_01220_),
    .RESETN(net969),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35019_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03212_),
    .QN(_01252_),
    .RESETN(net970),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35020_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03213_),
    .QN(_01286_),
    .RESETN(net971),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35021_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03214_),
    .QN(_00302_),
    .RESETN(net972),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35022_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03215_),
    .QN(_00256_),
    .RESETN(net973),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35023_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03216_),
    .QN(_00364_),
    .RESETN(net974),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35024_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03217_),
    .QN(_00395_),
    .RESETN(net975),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35025_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03218_),
    .QN(_00425_),
    .RESETN(net976),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35026_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03219_),
    .QN(_00455_),
    .RESETN(net977),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35027_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03220_),
    .QN(_00485_),
    .RESETN(net978),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35028_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03221_),
    .QN(_00515_),
    .RESETN(net979),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35029_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03222_),
    .QN(_00545_),
    .RESETN(net980),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35030_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03223_),
    .QN(_00575_),
    .RESETN(net981),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35031_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03224_),
    .QN(_00605_),
    .RESETN(net982),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35032_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03225_),
    .QN(_00635_),
    .RESETN(net983),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35033_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03226_),
    .QN(_00334_),
    .RESETN(net984),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35034_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03227_),
    .QN(_00697_),
    .RESETN(net985),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35035_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03228_),
    .QN(_00729_),
    .RESETN(net986),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35036_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03229_),
    .QN(_00762_),
    .RESETN(net987),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35037_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03230_),
    .QN(_00795_),
    .RESETN(net988),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35038_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03231_),
    .QN(_00828_),
    .RESETN(net989),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35039_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03232_),
    .QN(_00860_),
    .RESETN(net990),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35040_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03233_),
    .QN(_00893_),
    .RESETN(net991),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35041_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03234_),
    .QN(_00925_),
    .RESETN(net992),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35042_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03235_),
    .QN(_00958_),
    .RESETN(net993),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35043_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03236_),
    .QN(_00990_),
    .RESETN(net994),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35044_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03237_),
    .QN(_01024_),
    .RESETN(net995),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35045_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03238_),
    .QN(_01056_),
    .RESETN(net996),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35046_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03239_),
    .QN(_01089_),
    .RESETN(net997),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35047_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03240_),
    .QN(_01121_),
    .RESETN(net998),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35048_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03241_),
    .QN(_01155_),
    .RESETN(net999),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35049_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03242_),
    .QN(_01187_),
    .RESETN(net1000),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35050_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03243_),
    .QN(_01221_),
    .RESETN(net1001),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35051_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03244_),
    .QN(_01253_),
    .RESETN(net1002),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35052_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03245_),
    .QN(_01287_),
    .RESETN(net1003),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35053_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03246_),
    .QN(_00303_),
    .RESETN(net1004),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35054_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03247_),
    .QN(_00257_),
    .RESETN(net1005),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35055_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03248_),
    .QN(_00365_),
    .RESETN(net1006),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35056_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03249_),
    .QN(_00396_),
    .RESETN(net1007),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35057_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03250_),
    .QN(_00426_),
    .RESETN(net1008),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35058_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03251_),
    .QN(_00456_),
    .RESETN(net1009),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35059_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03252_),
    .QN(_00486_),
    .RESETN(net1010),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35060_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03253_),
    .QN(_00516_),
    .RESETN(net1011),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35061_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03254_),
    .QN(_00546_),
    .RESETN(net1012),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35062_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03255_),
    .QN(_00576_),
    .RESETN(net1013),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35063_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03256_),
    .QN(_00606_),
    .RESETN(net1014),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35064_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03257_),
    .QN(_00636_),
    .RESETN(net1015),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35065_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03258_),
    .QN(_00335_),
    .RESETN(net1016),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35066_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03259_),
    .QN(_00698_),
    .RESETN(net1017),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35067_ (.CLK(clknet_level_3_1_34135_clk_i),
    .D(_03260_),
    .QN(_00730_),
    .RESETN(net1018),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35068_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03261_),
    .QN(_00763_),
    .RESETN(net1019),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35069_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03262_),
    .QN(_00796_),
    .RESETN(net1020),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35070_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03263_),
    .QN(_00829_),
    .RESETN(net1021),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35071_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03264_),
    .QN(_00861_),
    .RESETN(net1022),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35072_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03265_),
    .QN(_00894_),
    .RESETN(net1023),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35073_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03266_),
    .QN(_00926_),
    .RESETN(net1024),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35074_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03267_),
    .QN(_00959_),
    .RESETN(net1025),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35075_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03268_),
    .QN(_00991_),
    .RESETN(net1026),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35076_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03269_),
    .QN(_01025_),
    .RESETN(net1027),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35077_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03270_),
    .QN(_01057_),
    .RESETN(net1028),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35078_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03271_),
    .QN(_01090_),
    .RESETN(net1029),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35079_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03272_),
    .QN(_01122_),
    .RESETN(net1030),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35080_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03273_),
    .QN(_01156_),
    .RESETN(net1031),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35081_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03274_),
    .QN(_01188_),
    .RESETN(net1032),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35082_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03275_),
    .QN(_01222_),
    .RESETN(net1033),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35083_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03276_),
    .QN(_01254_),
    .RESETN(net1034),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35084_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03277_),
    .QN(_01288_),
    .RESETN(net1035),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35085_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03278_),
    .QN(_00304_),
    .RESETN(net1036),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35086_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03279_),
    .QN(_00258_),
    .RESETN(net1037),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35087_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03280_),
    .QN(_00366_),
    .RESETN(net1038),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35088_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03281_),
    .QN(_00397_),
    .RESETN(net1039),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35089_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03282_),
    .QN(_00427_),
    .RESETN(net1040),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35090_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03283_),
    .QN(_00457_),
    .RESETN(net1041),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35091_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03284_),
    .QN(_00487_),
    .RESETN(net1042),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35092_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03285_),
    .QN(_00517_),
    .RESETN(net1043),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35093_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03286_),
    .QN(_00547_),
    .RESETN(net1044),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35094_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03287_),
    .QN(_00577_),
    .RESETN(net1045),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35095_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03288_),
    .QN(_00607_),
    .RESETN(net1046),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35096_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03289_),
    .QN(_00637_),
    .RESETN(net1047),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35097_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03290_),
    .QN(_00336_),
    .RESETN(net1048),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35098_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03291_),
    .QN(_00699_),
    .RESETN(net1049),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35099_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03292_),
    .QN(_00731_),
    .RESETN(net1050),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35100_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03293_),
    .QN(_00764_),
    .RESETN(net1051),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35101_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03294_),
    .QN(_00797_),
    .RESETN(net1052),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35102_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03295_),
    .QN(_00830_),
    .RESETN(net1053),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35103_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03296_),
    .QN(_00862_),
    .RESETN(net1054),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35104_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03297_),
    .QN(_00895_),
    .RESETN(net1055),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35105_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03298_),
    .QN(_00927_),
    .RESETN(net1056),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35106_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03299_),
    .QN(_00960_),
    .RESETN(net1057),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35107_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03300_),
    .QN(_00992_),
    .RESETN(net1058),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35108_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03301_),
    .QN(_01026_),
    .RESETN(net1059),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35109_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03302_),
    .QN(_01058_),
    .RESETN(net1060),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35110_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03303_),
    .QN(_01091_),
    .RESETN(net1061),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35111_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03304_),
    .QN(_01123_),
    .RESETN(net1062),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35112_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03305_),
    .QN(_01157_),
    .RESETN(net1063),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35113_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03306_),
    .QN(_01189_),
    .RESETN(net1064),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35114_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03307_),
    .QN(_01223_),
    .RESETN(net1065),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35115_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03308_),
    .QN(_01255_),
    .RESETN(net1066),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35116_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03309_),
    .QN(_01289_),
    .RESETN(net1067),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35117_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03310_),
    .QN(_00305_),
    .RESETN(net1068),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35118_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03311_),
    .QN(_00259_),
    .RESETN(net1069),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35119_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03312_),
    .QN(_00367_),
    .RESETN(net1070),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35120_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03313_),
    .QN(_00398_),
    .RESETN(net1071),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35121_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03314_),
    .QN(_00428_),
    .RESETN(net1072),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35122_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03315_),
    .QN(_00458_),
    .RESETN(net1073),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35123_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03316_),
    .QN(_00488_),
    .RESETN(net1074),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35124_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03317_),
    .QN(_00518_),
    .RESETN(net1075),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35125_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03318_),
    .QN(_00548_),
    .RESETN(net1076),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35126_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03319_),
    .QN(_00578_),
    .RESETN(net1077),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35127_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03320_),
    .QN(_00608_),
    .RESETN(net1078),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35128_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03321_),
    .QN(_00638_),
    .RESETN(net1079),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35129_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03322_),
    .QN(_00337_),
    .RESETN(net1080),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35130_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03323_),
    .QN(_00700_),
    .RESETN(net1081),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35131_ (.CLK(clknet_level_3_1_34135_clk_i),
    .D(_03324_),
    .QN(_00732_),
    .RESETN(net1082),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35132_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03325_),
    .QN(_00765_),
    .RESETN(net1083),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35133_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03326_),
    .QN(_00798_),
    .RESETN(net1084),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35134_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03327_),
    .QN(_00831_),
    .RESETN(net1085),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35135_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03328_),
    .QN(_00863_),
    .RESETN(net1086),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35136_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03329_),
    .QN(_00896_),
    .RESETN(net1087),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35137_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03330_),
    .QN(_00928_),
    .RESETN(net1088),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35138_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03331_),
    .QN(_00961_),
    .RESETN(net1089),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35139_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03332_),
    .QN(_00993_),
    .RESETN(net1090),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35140_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03333_),
    .QN(_01027_),
    .RESETN(net1091),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35141_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03334_),
    .QN(_01059_),
    .RESETN(net1092),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35142_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03335_),
    .QN(_01092_),
    .RESETN(net1093),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35143_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03336_),
    .QN(_01124_),
    .RESETN(net1094),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35144_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03337_),
    .QN(_01158_),
    .RESETN(net1095),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35145_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03338_),
    .QN(_01190_),
    .RESETN(net1096),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35146_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03339_),
    .QN(_01224_),
    .RESETN(net1097),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35147_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03340_),
    .QN(_01256_),
    .RESETN(net1098),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35148_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03341_),
    .QN(_01290_),
    .RESETN(net1099),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35149_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03342_),
    .QN(_00306_),
    .RESETN(net1100),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35150_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03343_),
    .QN(_00260_),
    .RESETN(net1101),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35151_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03344_),
    .QN(_00368_),
    .RESETN(net1102),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35152_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03345_),
    .QN(_00399_),
    .RESETN(net1103),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35153_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03346_),
    .QN(_00429_),
    .RESETN(net1104),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35154_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03347_),
    .QN(_00459_),
    .RESETN(net1105),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35155_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03348_),
    .QN(_00489_),
    .RESETN(net1106),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35156_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03349_),
    .QN(_00519_),
    .RESETN(net1107),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35157_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03350_),
    .QN(_00549_),
    .RESETN(net1108),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35158_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03351_),
    .QN(_00579_),
    .RESETN(net1109),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35159_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03352_),
    .QN(_00609_),
    .RESETN(net1110),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35160_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03353_),
    .QN(_00639_),
    .RESETN(net1111),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35161_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03354_),
    .QN(_00338_),
    .RESETN(net1112),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35162_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03355_),
    .QN(_00701_),
    .RESETN(net1113),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35163_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03356_),
    .QN(_00733_),
    .RESETN(net1114),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35164_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03357_),
    .QN(_00766_),
    .RESETN(net1115),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35165_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03358_),
    .QN(_00799_),
    .RESETN(net1116),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35166_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03359_),
    .QN(_00832_),
    .RESETN(net1117),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35167_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03360_),
    .QN(_00864_),
    .RESETN(net1118),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35168_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03361_),
    .QN(_00897_),
    .RESETN(net1119),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35169_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03362_),
    .QN(_00929_),
    .RESETN(net1120),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35170_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03363_),
    .QN(_00962_),
    .RESETN(net1121),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35171_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03364_),
    .QN(_00994_),
    .RESETN(net1122),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35172_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03365_),
    .QN(_01028_),
    .RESETN(net1123),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35173_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03366_),
    .QN(_01060_),
    .RESETN(net1124),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35174_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03367_),
    .QN(_01093_),
    .RESETN(net1125),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35175_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03368_),
    .QN(_01125_),
    .RESETN(net1126),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35176_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03369_),
    .QN(_01159_),
    .RESETN(net1127),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35177_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03370_),
    .QN(_01191_),
    .RESETN(net1128),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35178_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03371_),
    .QN(_01225_),
    .RESETN(net1129),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35179_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03372_),
    .QN(_01257_),
    .RESETN(net1130),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35180_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03373_),
    .QN(_01291_),
    .RESETN(net1131),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35181_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03374_),
    .QN(_00307_),
    .RESETN(net1132),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35182_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03375_),
    .QN(_00261_),
    .RESETN(net1133),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35183_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03376_),
    .QN(_00369_),
    .RESETN(net1134),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35184_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03377_),
    .QN(_00400_),
    .RESETN(net1135),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35185_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03378_),
    .QN(_00430_),
    .RESETN(net1136),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35186_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03379_),
    .QN(_00460_),
    .RESETN(net1137),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35187_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03380_),
    .QN(_00490_),
    .RESETN(net1138),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35188_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03381_),
    .QN(_00520_),
    .RESETN(net1139),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35189_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03382_),
    .QN(_00550_),
    .RESETN(net1140),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35190_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03383_),
    .QN(_00580_),
    .RESETN(net1141),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35191_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03384_),
    .QN(_00610_),
    .RESETN(net1142),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35192_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03385_),
    .QN(_00640_),
    .RESETN(net1143),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35193_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03386_),
    .QN(_00339_),
    .RESETN(net1144),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35194_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03387_),
    .QN(_00702_),
    .RESETN(net1145),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35195_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03388_),
    .QN(_00734_),
    .RESETN(net1146),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35196_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03389_),
    .QN(_00767_),
    .RESETN(net1147),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35197_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03390_),
    .QN(_00800_),
    .RESETN(net1148),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35198_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03391_),
    .QN(_00833_),
    .RESETN(net1149),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35199_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03392_),
    .QN(_00865_),
    .RESETN(net1150),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35200_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03393_),
    .QN(_00898_),
    .RESETN(net1151),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35201_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03394_),
    .QN(_00930_),
    .RESETN(net1152),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35202_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03395_),
    .QN(_00963_),
    .RESETN(net1153),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35203_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03396_),
    .QN(_00995_),
    .RESETN(net1154),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35204_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03397_),
    .QN(_01029_),
    .RESETN(net1155),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35205_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03398_),
    .QN(_01061_),
    .RESETN(net1156),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35206_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03399_),
    .QN(_01094_),
    .RESETN(net1157),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35207_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03400_),
    .QN(_01126_),
    .RESETN(net1158),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35208_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03401_),
    .QN(_01160_),
    .RESETN(net1159),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35209_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03402_),
    .QN(_01192_),
    .RESETN(net1160),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35210_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03403_),
    .QN(_01226_),
    .RESETN(net1161),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35211_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03404_),
    .QN(_01258_),
    .RESETN(net1162),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35212_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03405_),
    .QN(_01292_),
    .RESETN(net1163),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35213_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03406_),
    .QN(_00308_),
    .RESETN(net1164),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35214_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03407_),
    .QN(_00262_),
    .RESETN(net1165),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35215_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03408_),
    .QN(_00370_),
    .RESETN(net1166),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35216_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03409_),
    .QN(_00401_),
    .RESETN(net1167),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35217_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03410_),
    .QN(_00431_),
    .RESETN(net1168),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35218_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03411_),
    .QN(_00461_),
    .RESETN(net1169),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35219_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03412_),
    .QN(_00491_),
    .RESETN(net1170),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35220_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03413_),
    .QN(_00521_),
    .RESETN(net1171),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35221_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03414_),
    .QN(_00551_),
    .RESETN(net1172),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35222_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03415_),
    .QN(_00581_),
    .RESETN(net1173),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35223_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03416_),
    .QN(_00611_),
    .RESETN(net1174),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35224_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03417_),
    .QN(_00641_),
    .RESETN(net1175),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35225_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03418_),
    .QN(_00340_),
    .RESETN(net1176),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35226_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03419_),
    .QN(_00703_),
    .RESETN(net1177),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35227_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03420_),
    .QN(_00735_),
    .RESETN(net1178),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35228_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03421_),
    .QN(_00768_),
    .RESETN(net1179),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35229_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03422_),
    .QN(_00801_),
    .RESETN(net1180),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35230_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03423_),
    .QN(_00834_),
    .RESETN(net1181),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35231_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03424_),
    .QN(_00866_),
    .RESETN(net1182),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35232_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03425_),
    .QN(_00899_),
    .RESETN(net1183),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35233_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03426_),
    .QN(_00931_),
    .RESETN(net1184),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35234_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03427_),
    .QN(_00964_),
    .RESETN(net1185),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35235_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03428_),
    .QN(_00996_),
    .RESETN(net1186),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35236_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03429_),
    .QN(_01030_),
    .RESETN(net1187),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35237_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03430_),
    .QN(_01062_),
    .RESETN(net1188),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35238_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03431_),
    .QN(_01095_),
    .RESETN(net1189),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35239_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03432_),
    .QN(_01127_),
    .RESETN(net1190),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35240_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03433_),
    .QN(_01161_),
    .RESETN(net1191),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35241_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03434_),
    .QN(_01193_),
    .RESETN(net1192),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35242_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03435_),
    .QN(_01227_),
    .RESETN(net1193),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35243_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03436_),
    .QN(_01259_),
    .RESETN(net1194),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35244_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03437_),
    .QN(_01293_),
    .RESETN(net1195),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35245_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03438_),
    .QN(_00309_),
    .RESETN(net1196),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35246_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03439_),
    .QN(_00263_),
    .RESETN(net1197),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35247_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03440_),
    .QN(_00371_),
    .RESETN(net1198),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35248_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03441_),
    .QN(_00402_),
    .RESETN(net1199),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35249_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03442_),
    .QN(_00432_),
    .RESETN(net1200),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35250_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03443_),
    .QN(_00462_),
    .RESETN(net1201),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35251_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03444_),
    .QN(_00492_),
    .RESETN(net1202),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35252_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03445_),
    .QN(_00522_),
    .RESETN(net1203),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35253_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03446_),
    .QN(_00552_),
    .RESETN(net1204),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35254_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03447_),
    .QN(_00582_),
    .RESETN(net1205),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35255_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03448_),
    .QN(_00612_),
    .RESETN(net1206),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35256_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03449_),
    .QN(_00642_),
    .RESETN(net1207),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35257_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03450_),
    .QN(_00341_),
    .RESETN(net1208),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35258_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03451_),
    .QN(_00704_),
    .RESETN(net1209),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35259_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03452_),
    .QN(_00736_),
    .RESETN(net1210),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35260_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03453_),
    .QN(_00769_),
    .RESETN(net1211),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35261_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03454_),
    .QN(_00802_),
    .RESETN(net1212),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35262_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03455_),
    .QN(_00835_),
    .RESETN(net1213),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35263_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03456_),
    .QN(_00867_),
    .RESETN(net1214),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35264_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03457_),
    .QN(_00900_),
    .RESETN(net1215),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35265_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03458_),
    .QN(_00932_),
    .RESETN(net1216),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35266_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03459_),
    .QN(_00965_),
    .RESETN(net1217),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35267_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03460_),
    .QN(_00997_),
    .RESETN(net1218),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35268_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03461_),
    .QN(_01031_),
    .RESETN(net1219),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35269_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03462_),
    .QN(_01063_),
    .RESETN(net1220),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35270_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03463_),
    .QN(_01096_),
    .RESETN(net1221),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35271_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03464_),
    .QN(_01128_),
    .RESETN(net1222),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35272_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03465_),
    .QN(_01162_),
    .RESETN(net1223),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35273_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03466_),
    .QN(_01194_),
    .RESETN(net1224),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35274_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03467_),
    .QN(_01228_),
    .RESETN(net1225),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35275_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03468_),
    .QN(_01260_),
    .RESETN(net1226),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35276_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03469_),
    .QN(_01294_),
    .RESETN(net1227),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35277_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03470_),
    .QN(_00310_),
    .RESETN(net1228),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35278_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03471_),
    .QN(_00264_),
    .RESETN(net1229),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35279_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03472_),
    .QN(_00372_),
    .RESETN(net1230),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35280_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03473_),
    .QN(_00403_),
    .RESETN(net1231),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35281_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03474_),
    .QN(_00433_),
    .RESETN(net1232),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35282_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03475_),
    .QN(_00463_),
    .RESETN(net1233),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35283_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03476_),
    .QN(_00493_),
    .RESETN(net1234),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35284_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03477_),
    .QN(_00523_),
    .RESETN(net1235),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35285_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03478_),
    .QN(_00553_),
    .RESETN(net1236),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35286_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03479_),
    .QN(_00583_),
    .RESETN(net1237),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35287_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03480_),
    .QN(_00613_),
    .RESETN(net1238),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35288_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03481_),
    .QN(_00643_),
    .RESETN(net1239),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35289_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03482_),
    .QN(_00342_),
    .RESETN(net1240),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35290_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03483_),
    .QN(_00705_),
    .RESETN(net1241),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35291_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03484_),
    .QN(_00737_),
    .RESETN(net1242),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35292_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03485_),
    .QN(_00770_),
    .RESETN(net1243),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35293_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03486_),
    .QN(_00803_),
    .RESETN(net1244),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35294_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03487_),
    .QN(_00836_),
    .RESETN(net1245),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35295_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03488_),
    .QN(_00868_),
    .RESETN(net1246),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35296_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03489_),
    .QN(_00901_),
    .RESETN(net1247),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35297_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03490_),
    .QN(_00933_),
    .RESETN(net1248),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35298_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03491_),
    .QN(_00966_),
    .RESETN(net1249),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35299_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03492_),
    .QN(_00998_),
    .RESETN(net1250),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35300_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03493_),
    .QN(_01032_),
    .RESETN(net1251),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35301_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03494_),
    .QN(_01064_),
    .RESETN(net1252),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35302_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03495_),
    .QN(_01097_),
    .RESETN(net1253),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35303_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03496_),
    .QN(_01129_),
    .RESETN(net1254),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35304_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03497_),
    .QN(_01163_),
    .RESETN(net1255),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35305_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03498_),
    .QN(_01195_),
    .RESETN(net1256),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35306_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03499_),
    .QN(_01229_),
    .RESETN(net1257),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35307_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03500_),
    .QN(_01261_),
    .RESETN(net1258),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35308_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03501_),
    .QN(_01295_),
    .RESETN(net1259),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35309_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03502_),
    .QN(_00311_),
    .RESETN(net1260),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35310_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03503_),
    .QN(_00265_),
    .RESETN(net1261),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35311_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03504_),
    .QN(_00373_),
    .RESETN(net1262),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35312_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03505_),
    .QN(_00404_),
    .RESETN(net1263),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35313_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03506_),
    .QN(_00434_),
    .RESETN(net1264),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35314_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03507_),
    .QN(_00464_),
    .RESETN(net1265),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35315_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03508_),
    .QN(_00494_),
    .RESETN(net1266),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35316_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03509_),
    .QN(_00524_),
    .RESETN(net1267),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35317_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03510_),
    .QN(_00554_),
    .RESETN(net1268),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35318_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03511_),
    .QN(_00584_),
    .RESETN(net1269),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35319_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03512_),
    .QN(_00614_),
    .RESETN(net1270),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35320_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03513_),
    .QN(_00644_),
    .RESETN(net1271),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35321_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03514_),
    .QN(_00343_),
    .RESETN(net1272),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35322_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03515_),
    .QN(_00706_),
    .RESETN(net1273),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35323_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03516_),
    .QN(_00738_),
    .RESETN(net1274),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35324_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03517_),
    .QN(_00771_),
    .RESETN(net1275),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35325_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03518_),
    .QN(_00804_),
    .RESETN(net1276),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35326_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03519_),
    .QN(_00837_),
    .RESETN(net1277),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35327_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03520_),
    .QN(_00869_),
    .RESETN(net1278),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35328_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03521_),
    .QN(_00902_),
    .RESETN(net1279),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35329_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03522_),
    .QN(_00934_),
    .RESETN(net1280),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35330_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03523_),
    .QN(_00967_),
    .RESETN(net1281),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35331_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03524_),
    .QN(_00999_),
    .RESETN(net1282),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35332_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03525_),
    .QN(_01033_),
    .RESETN(net1283),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35333_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03526_),
    .QN(_01065_),
    .RESETN(net1284),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35334_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03527_),
    .QN(_01098_),
    .RESETN(net1285),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35335_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03528_),
    .QN(_01130_),
    .RESETN(net1286),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35336_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03529_),
    .QN(_01164_),
    .RESETN(net1287),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35337_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03530_),
    .QN(_01196_),
    .RESETN(net1288),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35338_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03531_),
    .QN(_01230_),
    .RESETN(net1289),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35339_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03532_),
    .QN(_01262_),
    .RESETN(net1290),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35340_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03533_),
    .QN(_01296_),
    .RESETN(net1291),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35341_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03534_),
    .QN(_00312_),
    .RESETN(net1292),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35342_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03535_),
    .QN(_00266_),
    .RESETN(net1293),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35343_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03536_),
    .QN(_00374_),
    .RESETN(net1294),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35344_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03537_),
    .QN(_00405_),
    .RESETN(net1295),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35345_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03538_),
    .QN(_00435_),
    .RESETN(net1296),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35346_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03539_),
    .QN(_00465_),
    .RESETN(net1297),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35347_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03540_),
    .QN(_00495_),
    .RESETN(net1298),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35348_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03541_),
    .QN(_00525_),
    .RESETN(net1299),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35349_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03542_),
    .QN(_00555_),
    .RESETN(net1300),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35350_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03543_),
    .QN(_00585_),
    .RESETN(net1301),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35351_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03544_),
    .QN(_00615_),
    .RESETN(net1302),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35352_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03545_),
    .QN(_00645_),
    .RESETN(net1303),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35353_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03546_),
    .QN(_00344_),
    .RESETN(net1304),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35354_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03547_),
    .QN(_00707_),
    .RESETN(net1305),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35355_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03548_),
    .QN(_00739_),
    .RESETN(net1306),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35356_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03549_),
    .QN(_00772_),
    .RESETN(net1307),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35357_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03550_),
    .QN(_00805_),
    .RESETN(net1308),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35358_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03551_),
    .QN(_00838_),
    .RESETN(net1309),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35359_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03552_),
    .QN(_00870_),
    .RESETN(net1310),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35360_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03553_),
    .QN(_00903_),
    .RESETN(net1311),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35361_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03554_),
    .QN(_00935_),
    .RESETN(net1312),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35362_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03555_),
    .QN(_00968_),
    .RESETN(net1313),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35363_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03556_),
    .QN(_01000_),
    .RESETN(net1314),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35364_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03557_),
    .QN(_01034_),
    .RESETN(net1315),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35365_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03558_),
    .QN(_01066_),
    .RESETN(net1316),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35366_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03559_),
    .QN(_01099_),
    .RESETN(net1317),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35367_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03560_),
    .QN(_01131_),
    .RESETN(net1318),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35368_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03561_),
    .QN(_01165_),
    .RESETN(net1319),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35369_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03562_),
    .QN(_01197_),
    .RESETN(net1320),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35370_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03563_),
    .QN(_01231_),
    .RESETN(net1321),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35371_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03564_),
    .QN(_01263_),
    .RESETN(net1322),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35372_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03565_),
    .QN(_01297_),
    .RESETN(net1323),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35373_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03566_),
    .QN(_00313_),
    .RESETN(net1324),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35374_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03567_),
    .QN(_00267_),
    .RESETN(net1325),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35375_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03568_),
    .QN(_00375_),
    .RESETN(net1326),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35376_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03569_),
    .QN(_00406_),
    .RESETN(net1327),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35377_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03570_),
    .QN(_00436_),
    .RESETN(net1328),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35378_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03571_),
    .QN(_00466_),
    .RESETN(net1329),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35379_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03572_),
    .QN(_00496_),
    .RESETN(net1330),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35380_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03573_),
    .QN(_00526_),
    .RESETN(net1331),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35381_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03574_),
    .QN(_00556_),
    .RESETN(net1332),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35382_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03575_),
    .QN(_00586_),
    .RESETN(net1333),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35383_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03576_),
    .QN(_00616_),
    .RESETN(net1334),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35384_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03577_),
    .QN(_00646_),
    .RESETN(net1335),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35385_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03578_),
    .QN(_00345_),
    .RESETN(net1336),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35386_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03579_),
    .QN(_00708_),
    .RESETN(net1337),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35387_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03580_),
    .QN(_00740_),
    .RESETN(net1338),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35388_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03581_),
    .QN(_00773_),
    .RESETN(net1339),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35389_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03582_),
    .QN(_00806_),
    .RESETN(net1340),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35390_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03583_),
    .QN(_00839_),
    .RESETN(net1341),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35391_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03584_),
    .QN(_00871_),
    .RESETN(net1342),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35392_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03585_),
    .QN(_00904_),
    .RESETN(net1343),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35393_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03586_),
    .QN(_00936_),
    .RESETN(net1344),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35394_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03587_),
    .QN(_00969_),
    .RESETN(net1345),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35395_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03588_),
    .QN(_01001_),
    .RESETN(net1346),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35396_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03589_),
    .QN(_01035_),
    .RESETN(net1347),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35397_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03590_),
    .QN(_01067_),
    .RESETN(net1348),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35398_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03591_),
    .QN(_01100_),
    .RESETN(net1349),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35399_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03592_),
    .QN(_01132_),
    .RESETN(net1350),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35400_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03593_),
    .QN(_01166_),
    .RESETN(net1351),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35401_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03594_),
    .QN(_01198_),
    .RESETN(net1352),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35402_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03595_),
    .QN(_01232_),
    .RESETN(net1353),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35403_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03596_),
    .QN(_01264_),
    .RESETN(net1354),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35404_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03597_),
    .QN(_01298_),
    .RESETN(net1355),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35405_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03598_),
    .QN(_00314_),
    .RESETN(net1356),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35406_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03599_),
    .QN(_00268_),
    .RESETN(net1357),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35407_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03600_),
    .QN(_00376_),
    .RESETN(net1358),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35408_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03601_),
    .QN(_00407_),
    .RESETN(net1359),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35409_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03602_),
    .QN(_00437_),
    .RESETN(net1360),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35410_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03603_),
    .QN(_00467_),
    .RESETN(net1361),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35411_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03604_),
    .QN(_00497_),
    .RESETN(net1362),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35412_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03605_),
    .QN(_00527_),
    .RESETN(net1363),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35413_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03606_),
    .QN(_00557_),
    .RESETN(net1364),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35414_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03607_),
    .QN(_00587_),
    .RESETN(net1365),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35415_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03608_),
    .QN(_00617_),
    .RESETN(net1366),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35416_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03609_),
    .QN(_00647_),
    .RESETN(net1367),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35417_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03610_),
    .QN(_00346_),
    .RESETN(net1368),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35418_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03611_),
    .QN(_00709_),
    .RESETN(net1369),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35419_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03612_),
    .QN(_00741_),
    .RESETN(net1370),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35420_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03613_),
    .QN(_00774_),
    .RESETN(net1371),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35421_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03614_),
    .QN(_00807_),
    .RESETN(net1372),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35422_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03615_),
    .QN(_00840_),
    .RESETN(net1373),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35423_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03616_),
    .QN(_00872_),
    .RESETN(net1374),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35424_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03617_),
    .QN(_00905_),
    .RESETN(net1375),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35425_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03618_),
    .QN(_00937_),
    .RESETN(net1376),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35426_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03619_),
    .QN(_00970_),
    .RESETN(net1377),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35427_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03620_),
    .QN(_01002_),
    .RESETN(net1378),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35428_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03621_),
    .QN(_01036_),
    .RESETN(net1379),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35429_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03622_),
    .QN(_01068_),
    .RESETN(net1380),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35430_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03623_),
    .QN(_01101_),
    .RESETN(net1381),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35431_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03624_),
    .QN(_01133_),
    .RESETN(net1382),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35432_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03625_),
    .QN(_01167_),
    .RESETN(net1383),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35433_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03626_),
    .QN(_01199_),
    .RESETN(net1384),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35434_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03627_),
    .QN(_01233_),
    .RESETN(net1385),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35435_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03628_),
    .QN(_01265_),
    .RESETN(net1386),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35436_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03629_),
    .QN(_01299_),
    .RESETN(net1387),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35437_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03630_),
    .QN(_00315_),
    .RESETN(net1388),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35438_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03631_),
    .QN(_00269_),
    .RESETN(net1389),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35439_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03632_),
    .QN(_00377_),
    .RESETN(net1390),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35440_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03633_),
    .QN(_00408_),
    .RESETN(net1391),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35441_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03634_),
    .QN(_00438_),
    .RESETN(net1392),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35442_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03635_),
    .QN(_00468_),
    .RESETN(net1393),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35443_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03636_),
    .QN(_00498_),
    .RESETN(net1394),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35444_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03637_),
    .QN(_00528_),
    .RESETN(net1395),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35445_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03638_),
    .QN(_00558_),
    .RESETN(net1396),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35446_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03639_),
    .QN(_00588_),
    .RESETN(net1397),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35447_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03640_),
    .QN(_00618_),
    .RESETN(net1398),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35448_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03641_),
    .QN(_00648_),
    .RESETN(net1399),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35449_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03642_),
    .QN(_00347_),
    .RESETN(net1400),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35450_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03643_),
    .QN(_00710_),
    .RESETN(net1401),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35451_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03644_),
    .QN(_00742_),
    .RESETN(net1402),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35452_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03645_),
    .QN(_00775_),
    .RESETN(net1403),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35453_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03646_),
    .QN(_00808_),
    .RESETN(net1404),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35454_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03647_),
    .QN(_00841_),
    .RESETN(net1405),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35455_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03648_),
    .QN(_00873_),
    .RESETN(net1406),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35456_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03649_),
    .QN(_00906_),
    .RESETN(net1407),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35457_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03650_),
    .QN(_00938_),
    .RESETN(net1408),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35458_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03651_),
    .QN(_00971_),
    .RESETN(net1409),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35459_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03652_),
    .QN(_01003_),
    .RESETN(net1410),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35460_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03653_),
    .QN(_01037_),
    .RESETN(net1411),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35461_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03654_),
    .QN(_01069_),
    .RESETN(net1412),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35462_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03655_),
    .QN(_01102_),
    .RESETN(net1413),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35463_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03656_),
    .QN(_01134_),
    .RESETN(net1414),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35464_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03657_),
    .QN(_01168_),
    .RESETN(net1415),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35465_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03658_),
    .QN(_01200_),
    .RESETN(net1416),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35466_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03659_),
    .QN(_01234_),
    .RESETN(net1417),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35467_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03660_),
    .QN(_01266_),
    .RESETN(net1418),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35468_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03661_),
    .QN(_01300_),
    .RESETN(net1419),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35469_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03662_),
    .QN(_00316_),
    .RESETN(net1420),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35470_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03663_),
    .QN(_00270_),
    .RESETN(net1421),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35471_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03664_),
    .QN(_00378_),
    .RESETN(net1422),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35472_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03665_),
    .QN(_00409_),
    .RESETN(net1423),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35473_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03666_),
    .QN(_00439_),
    .RESETN(net1424),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35474_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03667_),
    .QN(_00469_),
    .RESETN(net1425),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35475_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03668_),
    .QN(_00499_),
    .RESETN(net1426),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35476_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03669_),
    .QN(_00529_),
    .RESETN(net1427),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35477_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03670_),
    .QN(_00559_),
    .RESETN(net1428),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35478_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03671_),
    .QN(_00589_),
    .RESETN(net1429),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35479_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03672_),
    .QN(_00619_),
    .RESETN(net1430),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35480_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03673_),
    .QN(_00649_),
    .RESETN(net1431),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35481_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03674_),
    .QN(_00348_),
    .RESETN(net1432),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35482_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03675_),
    .QN(_00711_),
    .RESETN(net1433),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35483_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03676_),
    .QN(_00743_),
    .RESETN(net1434),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35484_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03677_),
    .QN(_00776_),
    .RESETN(net1435),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35485_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03678_),
    .QN(_00809_),
    .RESETN(net1436),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35486_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03679_),
    .QN(_00842_),
    .RESETN(net1437),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35487_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03680_),
    .QN(_00874_),
    .RESETN(net1438),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35488_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03681_),
    .QN(_00907_),
    .RESETN(net1439),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35489_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03682_),
    .QN(_00939_),
    .RESETN(net1440),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35490_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03683_),
    .QN(_00972_),
    .RESETN(net1441),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35491_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03684_),
    .QN(_01004_),
    .RESETN(net1442),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35492_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03685_),
    .QN(_01038_),
    .RESETN(net1443),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35493_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03686_),
    .QN(_01070_),
    .RESETN(net1444),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35494_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03687_),
    .QN(_01103_),
    .RESETN(net1445),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35495_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03688_),
    .QN(_01135_),
    .RESETN(net1446),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35496_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03689_),
    .QN(_01169_),
    .RESETN(net1447),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35497_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03690_),
    .QN(_01201_),
    .RESETN(net1448),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35498_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03691_),
    .QN(_01235_),
    .RESETN(net1449),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35499_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03692_),
    .QN(_01267_),
    .RESETN(net1450),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35500_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03693_),
    .QN(_01301_),
    .RESETN(net1451),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35501_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03694_),
    .QN(_00317_),
    .RESETN(net1452),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35502_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03695_),
    .QN(_00271_),
    .RESETN(net1453),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35503_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03696_),
    .QN(_00379_),
    .RESETN(net1454),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35504_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03697_),
    .QN(_00410_),
    .RESETN(net1455),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35505_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03698_),
    .QN(_00440_),
    .RESETN(net1456),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35506_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03699_),
    .QN(_00470_),
    .RESETN(net1457),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35507_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03700_),
    .QN(_00500_),
    .RESETN(net1458),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35508_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03701_),
    .QN(_00530_),
    .RESETN(net1459),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35509_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03702_),
    .QN(_00560_),
    .RESETN(net1460),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35510_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03703_),
    .QN(_00590_),
    .RESETN(net1461),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35511_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03704_),
    .QN(_00620_),
    .RESETN(net1462),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35512_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03705_),
    .QN(_00650_),
    .RESETN(net1463),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35513_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03706_),
    .QN(_00349_),
    .RESETN(net1464),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35514_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03707_),
    .QN(_00712_),
    .RESETN(net1465),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35515_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03708_),
    .QN(_00744_),
    .RESETN(net1466),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35516_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03709_),
    .QN(_00777_),
    .RESETN(net1467),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35517_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03710_),
    .QN(_00810_),
    .RESETN(net1468),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35518_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03711_),
    .QN(_00843_),
    .RESETN(net1469),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35519_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03712_),
    .QN(_00875_),
    .RESETN(net1470),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35520_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03713_),
    .QN(_00908_),
    .RESETN(net1471),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35521_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03714_),
    .QN(_00940_),
    .RESETN(net1472),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35522_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03715_),
    .QN(_00973_),
    .RESETN(net1473),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35523_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03716_),
    .QN(_01005_),
    .RESETN(net1474),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35524_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03717_),
    .QN(_01039_),
    .RESETN(net1475),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35525_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03718_),
    .QN(_01071_),
    .RESETN(net1476),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35526_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03719_),
    .QN(_01104_),
    .RESETN(net1477),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35527_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03720_),
    .QN(_01136_),
    .RESETN(net1478),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35528_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03721_),
    .QN(_01170_),
    .RESETN(net1479),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35529_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03722_),
    .QN(_01202_),
    .RESETN(net1480),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35530_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03723_),
    .QN(_01236_),
    .RESETN(net1481),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35531_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03724_),
    .QN(_01268_),
    .RESETN(net1482),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35532_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03725_),
    .QN(_01302_),
    .RESETN(net1483),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35533_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03726_),
    .QN(_00318_),
    .RESETN(net1484),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35534_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03727_),
    .QN(_00272_),
    .RESETN(net1485),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35535_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03728_),
    .QN(_00380_),
    .RESETN(net1486),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35536_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03729_),
    .QN(_00411_),
    .RESETN(net1487),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35537_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03730_),
    .QN(_00441_),
    .RESETN(net1488),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35538_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03731_),
    .QN(_00471_),
    .RESETN(net1489),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35539_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03732_),
    .QN(_00501_),
    .RESETN(net1490),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35540_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03733_),
    .QN(_00531_),
    .RESETN(net1491),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35541_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03734_),
    .QN(_00561_),
    .RESETN(net1492),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35542_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03735_),
    .QN(_00591_),
    .RESETN(net1493),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35543_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03736_),
    .QN(_00621_),
    .RESETN(net1494),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35544_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03737_),
    .QN(_00651_),
    .RESETN(net1495),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35545_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03738_),
    .QN(_00350_),
    .RESETN(net1496),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35546_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03739_),
    .QN(_00713_),
    .RESETN(net1497),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35547_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03740_),
    .QN(_00745_),
    .RESETN(net1498),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35548_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03741_),
    .QN(_00778_),
    .RESETN(net1499),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35549_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03742_),
    .QN(_00811_),
    .RESETN(net1500),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35550_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03743_),
    .QN(_00844_),
    .RESETN(net1501),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35551_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03744_),
    .QN(_00876_),
    .RESETN(net1502),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35552_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03745_),
    .QN(_00909_),
    .RESETN(net1503),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35553_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03746_),
    .QN(_00941_),
    .RESETN(net1504),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35554_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03747_),
    .QN(_00974_),
    .RESETN(net1505),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35555_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03748_),
    .QN(_01006_),
    .RESETN(net1506),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35556_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03749_),
    .QN(_01040_),
    .RESETN(net1507),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35557_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03750_),
    .QN(_01072_),
    .RESETN(net1508),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35558_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03751_),
    .QN(_01105_),
    .RESETN(net1509),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35559_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03752_),
    .QN(_01137_),
    .RESETN(net1510),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35560_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03753_),
    .QN(_01171_),
    .RESETN(net1511),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35561_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03754_),
    .QN(_01203_),
    .RESETN(net1512),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35562_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03755_),
    .QN(_01237_),
    .RESETN(net1513),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35563_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03756_),
    .QN(_01269_),
    .RESETN(net1514),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35564_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03757_),
    .QN(_01303_),
    .RESETN(net1515),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35565_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03758_),
    .QN(_00319_),
    .RESETN(net1516),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35566_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03759_),
    .QN(_00273_),
    .RESETN(net1517),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35567_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03760_),
    .QN(_00381_),
    .RESETN(net1518),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35568_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03761_),
    .QN(_00412_),
    .RESETN(net1519),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35569_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03762_),
    .QN(_00442_),
    .RESETN(net1520),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35570_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03763_),
    .QN(_00472_),
    .RESETN(net1521),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35571_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03764_),
    .QN(_00502_),
    .RESETN(net1522),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35572_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03765_),
    .QN(_00532_),
    .RESETN(net1523),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35573_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03766_),
    .QN(_00562_),
    .RESETN(net1524),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35574_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03767_),
    .QN(_00592_),
    .RESETN(net1525),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35575_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03768_),
    .QN(_00622_),
    .RESETN(net1526),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35576_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03769_),
    .QN(_00652_),
    .RESETN(net1527),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35577_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03770_),
    .QN(_00351_),
    .RESETN(net1528),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35578_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03771_),
    .QN(_00714_),
    .RESETN(net1529),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35579_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03772_),
    .QN(_00746_),
    .RESETN(net1530),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35580_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03773_),
    .QN(_00779_),
    .RESETN(net1531),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35581_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03774_),
    .QN(_00812_),
    .RESETN(net1532),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35582_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03775_),
    .QN(_00845_),
    .RESETN(net1533),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35583_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03776_),
    .QN(_00877_),
    .RESETN(net1534),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35584_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03777_),
    .QN(_00910_),
    .RESETN(net1535),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35585_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03778_),
    .QN(_00942_),
    .RESETN(net1536),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35586_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03779_),
    .QN(_00975_),
    .RESETN(net1537),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35587_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03780_),
    .QN(_01007_),
    .RESETN(net1538),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35588_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03781_),
    .QN(_01041_),
    .RESETN(net1539),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35589_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03782_),
    .QN(_01073_),
    .RESETN(net1540),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35590_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03783_),
    .QN(_01106_),
    .RESETN(net1541),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35591_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03784_),
    .QN(_01138_),
    .RESETN(net1542),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35592_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03785_),
    .QN(_01172_),
    .RESETN(net1543),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35593_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03786_),
    .QN(_01204_),
    .RESETN(net1544),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35594_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03787_),
    .QN(_01238_),
    .RESETN(net1545),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35595_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03788_),
    .QN(_01270_),
    .RESETN(net1546),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35596_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03789_),
    .QN(_01304_),
    .RESETN(net1547),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35597_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03790_),
    .QN(_00320_),
    .RESETN(net1548),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35598_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03791_),
    .QN(_00274_),
    .RESETN(net1549),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35599_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03792_),
    .QN(_00382_),
    .RESETN(net1550),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35600_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03793_),
    .QN(_00413_),
    .RESETN(net1551),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35601_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03794_),
    .QN(_00443_),
    .RESETN(net1552),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35602_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03795_),
    .QN(_00473_),
    .RESETN(net1553),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35603_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03796_),
    .QN(_00503_),
    .RESETN(net1554),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35604_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03797_),
    .QN(_00533_),
    .RESETN(net1555),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35605_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03798_),
    .QN(_00563_),
    .RESETN(net1556),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35606_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03799_),
    .QN(_00593_),
    .RESETN(net1557),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35607_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03800_),
    .QN(_00623_),
    .RESETN(net1558),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35608_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03801_),
    .QN(_00653_),
    .RESETN(net1559),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35609_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03802_),
    .QN(_00352_),
    .RESETN(net1560),
    .SETN(net425));
 DFFASRHQNx1_ASAP7_75t_R _35610_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03803_),
    .QN(_00715_),
    .RESETN(net1561),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35611_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03804_),
    .QN(_00747_),
    .RESETN(net1562),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35612_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03805_),
    .QN(_00780_),
    .RESETN(net1563),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35613_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03806_),
    .QN(_00813_),
    .RESETN(net1564),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35614_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03807_),
    .QN(_00846_),
    .RESETN(net1565),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35615_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03808_),
    .QN(_00878_),
    .RESETN(net1566),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35616_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03809_),
    .QN(_00911_),
    .RESETN(net1567),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35617_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03810_),
    .QN(_00943_),
    .RESETN(net1568),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35618_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03811_),
    .QN(_00976_),
    .RESETN(net1569),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35619_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03812_),
    .QN(_01008_),
    .RESETN(net1570),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35620_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03813_),
    .QN(_01042_),
    .RESETN(net1571),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35621_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03814_),
    .QN(_01074_),
    .RESETN(net1572),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35622_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03815_),
    .QN(_01107_),
    .RESETN(net1573),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35623_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03816_),
    .QN(_01139_),
    .RESETN(net1574),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35624_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03817_),
    .QN(_01173_),
    .RESETN(net1575),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35625_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03818_),
    .QN(_01205_),
    .RESETN(net1576),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35626_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03819_),
    .QN(_01239_),
    .RESETN(net1577),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35627_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03820_),
    .QN(_01271_),
    .RESETN(net1578),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35628_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03821_),
    .QN(_01305_),
    .RESETN(net1579),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35629_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03822_),
    .QN(_00321_),
    .RESETN(net1580),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35630_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03823_),
    .QN(_00275_),
    .RESETN(net1581),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35631_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03824_),
    .QN(_00383_),
    .RESETN(net1582),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35632_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03825_),
    .QN(_00414_),
    .RESETN(net1583),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35633_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03826_),
    .QN(_00444_),
    .RESETN(net1584),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35634_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03827_),
    .QN(_00474_),
    .RESETN(net1585),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35635_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03828_),
    .QN(_00504_),
    .RESETN(net1586),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35636_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03829_),
    .QN(_00534_),
    .RESETN(net1587),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35637_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03830_),
    .QN(_00564_),
    .RESETN(net1588),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35638_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03831_),
    .QN(_00594_),
    .RESETN(net1589),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35639_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03832_),
    .QN(_00624_),
    .RESETN(net1590),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35640_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03833_),
    .QN(_00654_),
    .RESETN(net1591),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35641_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03834_),
    .QN(_00353_),
    .RESETN(net1592),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35642_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03835_),
    .QN(_00716_),
    .RESETN(net1593),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35643_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03836_),
    .QN(_00748_),
    .RESETN(net1594),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35644_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03837_),
    .QN(_00781_),
    .RESETN(net1595),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35645_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03838_),
    .QN(_00814_),
    .RESETN(net1596),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35646_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03839_),
    .QN(_00847_),
    .RESETN(net1597),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35647_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03840_),
    .QN(_00879_),
    .RESETN(net1598),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35648_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03841_),
    .QN(_00912_),
    .RESETN(net1599),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35649_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03842_),
    .QN(_00944_),
    .RESETN(net1600),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35650_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03843_),
    .QN(_00977_),
    .RESETN(net1601),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35651_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03844_),
    .QN(_01009_),
    .RESETN(net1602),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35652_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03845_),
    .QN(_01043_),
    .RESETN(net1603),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35653_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03846_),
    .QN(_01075_),
    .RESETN(net1604),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35654_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03847_),
    .QN(_01108_),
    .RESETN(net1605),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35655_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03848_),
    .QN(_01140_),
    .RESETN(net1606),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35656_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03849_),
    .QN(_01174_),
    .RESETN(net1607),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35657_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03850_),
    .QN(_01206_),
    .RESETN(net1608),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35658_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03851_),
    .QN(_01240_),
    .RESETN(net1609),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35659_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03852_),
    .QN(_01272_),
    .RESETN(net1610),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35660_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03853_),
    .QN(_01306_),
    .RESETN(net1611),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35661_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03854_),
    .QN(_00322_),
    .RESETN(net1612),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35662_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03855_),
    .QN(_00276_),
    .RESETN(net1613),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35663_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03856_),
    .QN(_00384_),
    .RESETN(net1614),
    .SETN(net429));
 DFFASRHQNx1_ASAP7_75t_R _35664_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03857_),
    .QN(_00415_),
    .RESETN(net1615),
    .SETN(net422));
 DFFASRHQNx1_ASAP7_75t_R _35665_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03858_),
    .QN(_00445_),
    .RESETN(net1616),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35666_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03859_),
    .QN(_00475_),
    .RESETN(net1617),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35667_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03860_),
    .QN(_00505_),
    .RESETN(net1618),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35668_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03861_),
    .QN(_00535_),
    .RESETN(net1619),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35669_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03862_),
    .QN(_00565_),
    .RESETN(net1620),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35670_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03863_),
    .QN(_00595_),
    .RESETN(net1621),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35671_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03864_),
    .QN(_00625_),
    .RESETN(net1622),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35672_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03865_),
    .QN(_00655_),
    .RESETN(net1623),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35673_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03866_),
    .QN(_00354_),
    .RESETN(net1624),
    .SETN(net428));
 DFFASRHQNx1_ASAP7_75t_R _35674_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03867_),
    .QN(_00717_),
    .RESETN(net1625),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35675_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03868_),
    .QN(_00749_),
    .RESETN(net1626),
    .SETN(net427));
 DFFASRHQNx1_ASAP7_75t_R _35676_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03869_),
    .QN(_00782_),
    .RESETN(net1627),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35677_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03870_),
    .QN(_00815_),
    .RESETN(net1628),
    .SETN(net431));
 DFFASRHQNx1_ASAP7_75t_R _35678_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03871_),
    .QN(_00848_),
    .RESETN(net1629),
    .SETN(net423));
 DFFASRHQNx1_ASAP7_75t_R _35679_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03872_),
    .QN(_00880_),
    .RESETN(net1630),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35680_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03873_),
    .QN(_00913_),
    .RESETN(net1631),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35681_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03874_),
    .QN(_00945_),
    .RESETN(net1632),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35682_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03875_),
    .QN(_00978_),
    .RESETN(net1633),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35683_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03876_),
    .QN(_01010_),
    .RESETN(net1634),
    .SETN(net426));
 DFFASRHQNx1_ASAP7_75t_R _35684_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03877_),
    .QN(_01044_),
    .RESETN(net1635),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _35685_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03878_),
    .QN(_01076_),
    .RESETN(net1636),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35686_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03879_),
    .QN(_01109_),
    .RESETN(net1637),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35687_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03880_),
    .QN(_01141_),
    .RESETN(net1638),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35688_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03881_),
    .QN(_01175_),
    .RESETN(net1639),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35689_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03882_),
    .QN(_01207_),
    .RESETN(net1640),
    .SETN(net430));
 DFFASRHQNx1_ASAP7_75t_R _35690_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03883_),
    .QN(_01241_),
    .RESETN(net1641),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35691_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03884_),
    .QN(_01273_),
    .RESETN(net1642),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35692_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03885_),
    .QN(_01307_),
    .RESETN(net1643),
    .SETN(net424));
 DFFASRHQNx1_ASAP7_75t_R _35693_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03886_),
    .QN(_01519_),
    .RESETN(net1644),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35694_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_03887_),
    .QN(_00659_),
    .RESETN(net1645),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35695_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_03888_),
    .QN(_01518_),
    .RESETN(net1646),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35696_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_03889_),
    .QN(_01517_),
    .RESETN(net1647),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35697_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_03890_),
    .QN(_01516_),
    .RESETN(net1648),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35698_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_03891_),
    .QN(_01515_),
    .RESETN(net1649),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35699_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_03892_),
    .QN(_01514_),
    .RESETN(net1650),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35700_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_03893_),
    .QN(_01513_),
    .RESETN(net1651),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35701_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_03894_),
    .QN(_01512_),
    .RESETN(net1652),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35702_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03895_),
    .QN(_01511_),
    .RESETN(net1653),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35703_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_03896_),
    .QN(_01510_),
    .RESETN(net1654),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35704_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03897_),
    .QN(_01509_),
    .RESETN(net1655),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35705_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03898_),
    .QN(_01508_),
    .RESETN(net1656),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35706_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03899_),
    .QN(_01507_),
    .RESETN(net1657),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35707_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03900_),
    .QN(_01506_),
    .RESETN(net1658),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35708_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03901_),
    .QN(_01505_),
    .RESETN(net1659),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35709_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03902_),
    .QN(_01504_),
    .RESETN(net1660),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35710_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03903_),
    .QN(_01503_),
    .RESETN(net1661),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35711_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03904_),
    .QN(_01502_),
    .RESETN(net1662),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35712_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03905_),
    .QN(_01501_),
    .RESETN(net1663),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35713_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03906_),
    .QN(_01500_),
    .RESETN(net1664),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35714_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03907_),
    .QN(_01499_),
    .RESETN(net1665),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35715_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03908_),
    .QN(_01498_),
    .RESETN(net1666),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35716_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03909_),
    .QN(_01497_),
    .RESETN(net1667),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35717_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03910_),
    .QN(_01496_),
    .RESETN(net1668),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35718_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03911_),
    .QN(_01495_),
    .RESETN(net1669),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35719_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03912_),
    .QN(_01494_),
    .RESETN(net1670),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35720_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03913_),
    .QN(_01493_),
    .RESETN(net1671),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35721_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03914_),
    .QN(_01492_),
    .RESETN(net1672),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35722_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_03915_),
    .QN(_01491_),
    .RESETN(net1673),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35723_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03916_),
    .QN(_01490_),
    .RESETN(net1674),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35724_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_03917_),
    .QN(_01489_),
    .RESETN(net1675),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35725_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_03918_),
    .QN(_01488_),
    .RESETN(net1676),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35726_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_03919_),
    .QN(_00660_),
    .RESETN(net1677),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35727_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_03920_),
    .QN(_01487_),
    .RESETN(net1678),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35728_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_03921_),
    .QN(_01486_),
    .RESETN(net1679),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35729_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_03922_),
    .QN(_01485_),
    .RESETN(net1680),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35730_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_03923_),
    .QN(_01484_),
    .RESETN(net1681),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35731_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_03924_),
    .QN(_01483_),
    .RESETN(net1682),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35732_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_03925_),
    .QN(_01482_),
    .RESETN(net1683),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35733_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_03926_),
    .QN(_01481_),
    .RESETN(net1684),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35734_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_03927_),
    .QN(_01480_),
    .RESETN(net1685),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35735_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_03928_),
    .QN(_01479_),
    .RESETN(net1686),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35736_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03929_),
    .QN(_01478_),
    .RESETN(net1687),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35737_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03930_),
    .QN(_01477_),
    .RESETN(net1688),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35738_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03931_),
    .QN(_01476_),
    .RESETN(net1689),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35739_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03932_),
    .QN(_01475_),
    .RESETN(net1690),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35740_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03933_),
    .QN(_01474_),
    .RESETN(net1691),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35741_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03934_),
    .QN(_01473_),
    .RESETN(net1692),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35742_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03935_),
    .QN(_01472_),
    .RESETN(net1693),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35743_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03936_),
    .QN(_01471_),
    .RESETN(net1694),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35744_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03937_),
    .QN(_01470_),
    .RESETN(net1695),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35745_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03938_),
    .QN(_01469_),
    .RESETN(net1696),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35746_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03939_),
    .QN(_01468_),
    .RESETN(net1697),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35747_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03940_),
    .QN(_01467_),
    .RESETN(net1698),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35748_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03941_),
    .QN(_01466_),
    .RESETN(net1699),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35749_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03942_),
    .QN(_01465_),
    .RESETN(net1700),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35750_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03943_),
    .QN(_01464_),
    .RESETN(net1701),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35751_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_03944_),
    .QN(_01463_),
    .RESETN(net1702),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35752_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03945_),
    .QN(_01462_),
    .RESETN(net1703),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35753_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03946_),
    .QN(_01461_),
    .RESETN(net1704),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35754_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_03947_),
    .QN(_01460_),
    .RESETN(net1705),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35755_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_03948_),
    .QN(_01459_),
    .RESETN(net1706),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35756_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_03949_),
    .QN(_01458_),
    .RESETN(net1707),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35757_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_03950_),
    .QN(_01457_),
    .RESETN(net1708),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35758_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_03951_),
    .QN(_01456_),
    .RESETN(net1709),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35759_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_03952_),
    .QN(_01455_),
    .RESETN(net1710),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35760_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_03953_),
    .QN(_01454_),
    .RESETN(net449),
    .SETN(net1711));
 DFFASRHQNx1_ASAP7_75t_R _35761_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_03954_),
    .QN(_01453_),
    .RESETN(net1712),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35762_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03955_),
    .QN(_01452_),
    .RESETN(net1713),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35763_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03956_),
    .QN(_01451_),
    .RESETN(net1714),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35764_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_03957_),
    .QN(_01450_),
    .RESETN(net1715),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35765_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03958_),
    .QN(_01449_),
    .RESETN(net1716),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35766_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03959_),
    .QN(_01448_),
    .RESETN(net1717),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35767_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_03960_),
    .QN(_01447_),
    .RESETN(net1718),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35768_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_03961_),
    .QN(_01446_),
    .RESETN(net1719),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35769_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_03962_),
    .QN(_01445_),
    .RESETN(net1720),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35770_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_03963_),
    .QN(_01444_),
    .RESETN(net1721),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35771_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03964_),
    .QN(_01443_),
    .RESETN(net1722),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35772_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_03965_),
    .QN(_01442_),
    .RESETN(net1723),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35773_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_03966_),
    .QN(_01441_),
    .RESETN(net1724),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35774_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_03967_),
    .QN(_02221_),
    .RESETN(net1725),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35775_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_03968_),
    .QN(_02220_),
    .RESETN(net1726),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35776_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03969_),
    .QN(_02219_),
    .RESETN(net1727),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35777_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_03970_),
    .QN(_02218_),
    .RESETN(net1728),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35778_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03971_),
    .QN(_02217_),
    .RESETN(net1729),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35779_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03972_),
    .QN(_02216_),
    .RESETN(net1730),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35780_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_03973_),
    .QN(_02215_),
    .RESETN(net1731),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35781_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_03974_),
    .QN(_02214_),
    .RESETN(net1732),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35782_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03975_),
    .QN(_02213_),
    .RESETN(net1733),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35783_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_03976_),
    .QN(_02212_),
    .RESETN(net1734),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35784_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_03977_),
    .QN(_02211_),
    .RESETN(net1735),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35785_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03978_),
    .QN(_02210_),
    .RESETN(net1736),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35786_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_03979_),
    .QN(_02209_),
    .RESETN(net1737),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35787_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03980_),
    .QN(_02208_),
    .RESETN(net1738),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35788_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_03981_),
    .QN(_02207_),
    .RESETN(net1739),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35789_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03982_),
    .QN(_02206_),
    .RESETN(net1740),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35790_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_03983_),
    .QN(_02205_),
    .RESETN(net1741),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35791_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03984_),
    .QN(_02204_),
    .RESETN(net1742),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35792_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03985_),
    .QN(_02203_),
    .RESETN(net1743),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35793_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_03986_),
    .QN(_02202_),
    .RESETN(net1744),
    .SETN(net443));
 DFFHQNx1_ASAP7_75t_R _35794_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_03987_),
    .QN(_02201_));
 DFFHQNx1_ASAP7_75t_R _35795_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_03988_),
    .QN(_02200_));
 DFFHQNx1_ASAP7_75t_R _35796_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_03989_),
    .QN(_02199_));
 DFFHQNx1_ASAP7_75t_R _35797_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_03990_),
    .QN(_02198_));
 DFFHQNx1_ASAP7_75t_R _35798_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_03991_),
    .QN(_02197_));
 DFFHQNx1_ASAP7_75t_R _35799_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_03992_),
    .QN(_02196_));
 DFFHQNx1_ASAP7_75t_R _35800_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_03993_),
    .QN(_02195_));
 DFFHQNx1_ASAP7_75t_R _35801_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_03994_),
    .QN(_02194_));
 DFFHQNx1_ASAP7_75t_R _35802_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_03995_),
    .QN(_02193_));
 DFFHQNx1_ASAP7_75t_R _35803_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_03996_),
    .QN(_02192_));
 DFFHQNx1_ASAP7_75t_R _35804_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_03997_),
    .QN(_02191_));
 DFFHQNx1_ASAP7_75t_R _35805_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_03998_),
    .QN(_02190_));
 DFFHQNx1_ASAP7_75t_R _35806_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_03999_),
    .QN(_02189_));
 DFFHQNx1_ASAP7_75t_R _35807_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_04000_),
    .QN(_02188_));
 DFFHQNx1_ASAP7_75t_R _35808_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_04001_),
    .QN(_02187_));
 DFFHQNx1_ASAP7_75t_R _35809_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04002_),
    .QN(_02186_));
 DFFHQNx1_ASAP7_75t_R _35810_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04003_),
    .QN(_02185_));
 DFFHQNx1_ASAP7_75t_R _35811_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04004_),
    .QN(_02184_));
 DFFHQNx1_ASAP7_75t_R _35812_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04005_),
    .QN(_02183_));
 DFFHQNx1_ASAP7_75t_R _35813_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04006_),
    .QN(_02182_));
 DFFHQNx1_ASAP7_75t_R _35814_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04007_),
    .QN(_02181_));
 DFFHQNx1_ASAP7_75t_R _35815_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04008_),
    .QN(_02180_));
 DFFHQNx1_ASAP7_75t_R _35816_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04009_),
    .QN(_02179_));
 DFFHQNx1_ASAP7_75t_R _35817_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04010_),
    .QN(_02178_));
 DFFHQNx1_ASAP7_75t_R _35818_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04011_),
    .QN(_02177_));
 DFFHQNx1_ASAP7_75t_R _35819_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04012_),
    .QN(_02176_));
 DFFHQNx1_ASAP7_75t_R _35820_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04013_),
    .QN(_02175_));
 DFFHQNx1_ASAP7_75t_R _35821_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04014_),
    .QN(_02174_));
 DFFHQNx1_ASAP7_75t_R _35822_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_04015_),
    .QN(_02173_));
 DFFHQNx1_ASAP7_75t_R _35823_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_04016_),
    .QN(_01729_));
 DFFASRHQNx1_ASAP7_75t_R _35824_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_00006_),
    .QN(_01730_),
    .RESETN(net1745),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35825_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_00007_),
    .QN(_01731_),
    .RESETN(net1746),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _35826_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_00000_),
    .QN(_01732_),
    .RESETN(net442),
    .SETN(net1747));
 DFFASRHQNx1_ASAP7_75t_R _35827_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_00001_),
    .QN(_01314_),
    .RESETN(net1748),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35828_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04017_),
    .QN(_02172_),
    .RESETN(net1749),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35829_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04018_),
    .QN(_02171_),
    .RESETN(net1750),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35830_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04019_),
    .QN(_02170_),
    .RESETN(net1751),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35831_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_04020_),
    .QN(_02169_),
    .RESETN(net1752),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35832_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04021_),
    .QN(_02168_),
    .RESETN(net1753),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35833_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04022_),
    .QN(_02167_),
    .RESETN(net1754),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35834_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04023_),
    .QN(_02166_),
    .RESETN(net1755),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35835_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04024_),
    .QN(_02165_),
    .RESETN(net1756),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35836_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04025_),
    .QN(_02164_),
    .RESETN(net1757),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35837_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04026_),
    .QN(_02163_),
    .RESETN(net1758),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35838_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04027_),
    .QN(_02162_),
    .RESETN(net1759),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35839_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04028_),
    .QN(_02161_),
    .RESETN(net1760),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35840_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04029_),
    .QN(_02160_),
    .RESETN(net1761),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35841_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04030_),
    .QN(_02159_),
    .RESETN(net1762),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35842_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04031_),
    .QN(_02158_),
    .RESETN(net1763),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35843_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04032_),
    .QN(_02157_),
    .RESETN(net1764),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35844_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04033_),
    .QN(_02156_),
    .RESETN(net1765),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35845_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04034_),
    .QN(_02155_),
    .RESETN(net1766),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35846_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04035_),
    .QN(_02154_),
    .RESETN(net1767),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35847_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04036_),
    .QN(_02153_),
    .RESETN(net1768),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35848_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04037_),
    .QN(_02152_),
    .RESETN(net1769),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35849_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04038_),
    .QN(_02151_),
    .RESETN(net1770),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35850_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04039_),
    .QN(_02150_),
    .RESETN(net1771),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35851_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04040_),
    .QN(_02149_),
    .RESETN(net1772),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35852_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04041_),
    .QN(_02148_),
    .RESETN(net1773),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35853_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04042_),
    .QN(_02147_),
    .RESETN(net1774),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35854_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04043_),
    .QN(_02146_),
    .RESETN(net1775),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35855_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04044_),
    .QN(_02145_),
    .RESETN(net1776),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35856_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04045_),
    .QN(_02144_),
    .RESETN(net1777),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35857_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04046_),
    .QN(_02143_),
    .RESETN(net1778),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35858_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04047_),
    .QN(_02142_),
    .RESETN(net1779),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35859_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_04048_),
    .QN(_02141_),
    .RESETN(net1780),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35860_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04049_),
    .QN(_02140_),
    .RESETN(net449),
    .SETN(net1781));
 DFFASRHQNx1_ASAP7_75t_R _35861_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04050_),
    .QN(_17592_),
    .RESETN(net449),
    .SETN(net1782));
 DFFASRHQNx1_ASAP7_75t_R _35862_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04051_),
    .QN(_02139_),
    .RESETN(net1783),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35863_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04052_),
    .QN(_02138_),
    .RESETN(net1784),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35864_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04053_),
    .QN(_02137_),
    .RESETN(net1785),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35865_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04054_),
    .QN(_02136_),
    .RESETN(net1786),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35866_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04055_),
    .QN(_02135_),
    .RESETN(net1787),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35867_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04056_),
    .QN(_02134_),
    .RESETN(net1788),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35868_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04057_),
    .QN(_02133_),
    .RESETN(net1789),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35869_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04058_),
    .QN(_02132_),
    .RESETN(net1790),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35870_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04059_),
    .QN(_02131_),
    .RESETN(net1791),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35871_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04060_),
    .QN(_02130_),
    .RESETN(net1792),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35872_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04061_),
    .QN(_02129_),
    .RESETN(net1793),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35873_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04062_),
    .QN(_02128_),
    .RESETN(net1794),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _35874_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04063_),
    .QN(_02127_),
    .RESETN(net1795),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35875_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04064_),
    .QN(_02126_),
    .RESETN(net1796),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35876_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04065_),
    .QN(_02125_),
    .RESETN(net1797),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _35877_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04066_),
    .QN(_02124_),
    .RESETN(net1798),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35878_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04067_),
    .QN(_02123_),
    .RESETN(net1799),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35879_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04068_),
    .QN(_02122_),
    .RESETN(net1800),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35880_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04069_),
    .QN(_02121_),
    .RESETN(net1801),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35881_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04070_),
    .QN(_02120_),
    .RESETN(net1802),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35882_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04071_),
    .QN(_02119_),
    .RESETN(net1803),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35883_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04072_),
    .QN(_02118_),
    .RESETN(net1804),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35884_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04073_),
    .QN(_02117_),
    .RESETN(net1805),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35885_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04074_),
    .QN(_02116_),
    .RESETN(net1806),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35886_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04075_),
    .QN(_02115_),
    .RESETN(net1807),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35887_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04076_),
    .QN(_02114_),
    .RESETN(net1808),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35888_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04077_),
    .QN(_02113_),
    .RESETN(net1809),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35889_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04078_),
    .QN(_02112_),
    .RESETN(net1810),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35890_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04079_),
    .QN(_02111_),
    .RESETN(net1811),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35891_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04080_),
    .QN(_02110_),
    .RESETN(net1812),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35892_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04081_),
    .QN(_02109_),
    .RESETN(net1813),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35893_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04082_),
    .QN(_02108_),
    .RESETN(net1814),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35894_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04083_),
    .QN(_02107_),
    .RESETN(net1815),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35895_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04084_),
    .QN(_02106_),
    .RESETN(net1816),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35896_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04085_),
    .QN(_02105_),
    .RESETN(net449),
    .SETN(net1817));
 DFFASRHQNx1_ASAP7_75t_R _35897_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04086_),
    .QN(_02104_),
    .RESETN(net1818),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35898_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04087_),
    .QN(_02103_),
    .RESETN(net1819),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _35899_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04088_),
    .QN(_02102_),
    .RESETN(net1820),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _35900_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04089_),
    .QN(_02101_),
    .RESETN(net1821),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35901_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04090_),
    .QN(_02100_),
    .RESETN(net1822),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35902_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04091_),
    .QN(_02099_),
    .RESETN(net1823),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35903_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04092_),
    .QN(_02098_),
    .RESETN(net1824),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35904_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04093_),
    .QN(_02097_),
    .RESETN(net1825),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35905_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04094_),
    .QN(_02096_),
    .RESETN(net1826),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35906_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04095_),
    .QN(_02095_),
    .RESETN(net1827),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35907_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04096_),
    .QN(_02094_),
    .RESETN(net1828),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35908_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04097_),
    .QN(_02093_),
    .RESETN(net1829),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35909_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04098_),
    .QN(_02092_),
    .RESETN(net1830),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35910_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04099_),
    .QN(_02091_),
    .RESETN(net1831),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _35911_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04100_),
    .QN(_02090_),
    .RESETN(net1832),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35912_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04101_),
    .QN(_02089_),
    .RESETN(net1833),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35913_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04102_),
    .QN(_02088_),
    .RESETN(net1834),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35914_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04103_),
    .QN(_02087_),
    .RESETN(net1835),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _35915_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04104_),
    .QN(_02086_),
    .RESETN(net1836),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35916_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04105_),
    .QN(_02085_),
    .RESETN(net1837),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35917_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04106_),
    .QN(_02084_),
    .RESETN(net1838),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35918_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04107_),
    .QN(_02083_),
    .RESETN(net1839),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35919_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04108_),
    .QN(_02082_),
    .RESETN(net1840),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35920_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04109_),
    .QN(_02081_),
    .RESETN(net1841),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35921_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04110_),
    .QN(_02080_),
    .RESETN(net1842),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _35922_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04111_),
    .QN(_02079_),
    .RESETN(net1843),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35923_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04112_),
    .QN(_02078_),
    .RESETN(net1844),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _35924_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04113_),
    .QN(_02077_),
    .RESETN(net1845),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35925_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04114_),
    .QN(_02076_),
    .RESETN(net1846),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35926_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04115_),
    .QN(_02075_),
    .RESETN(net1847),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35927_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04116_),
    .QN(_02074_),
    .RESETN(net1848),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35928_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04117_),
    .QN(_02073_),
    .RESETN(net1849),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35929_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04118_),
    .QN(_02072_),
    .RESETN(net1850),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _35930_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04119_),
    .QN(_02071_),
    .RESETN(net1851),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35931_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04120_),
    .QN(_02070_),
    .RESETN(net1852),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35932_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04121_),
    .QN(_02069_),
    .RESETN(net1853),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35933_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04122_),
    .QN(_02068_),
    .RESETN(net1854),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35934_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04123_),
    .QN(_02067_),
    .RESETN(net1855),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35935_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04124_),
    .QN(_00095_),
    .RESETN(net1856),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35936_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04125_),
    .QN(_00098_),
    .RESETN(net1857),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35937_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04126_),
    .QN(_00101_),
    .RESETN(net1858),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35938_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04127_),
    .QN(_00657_),
    .RESETN(net1859),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35939_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04128_),
    .QN(_00656_),
    .RESETN(net1860),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35940_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04129_),
    .QN(_00108_),
    .RESETN(net1861),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _35941_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04130_),
    .QN(_00111_),
    .RESETN(net1862),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35942_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04131_),
    .QN(_00114_),
    .RESETN(net1863),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35943_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04132_),
    .QN(_00117_),
    .RESETN(net1864),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35944_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04133_),
    .QN(_00120_),
    .RESETN(net1865),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _35945_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04134_),
    .QN(_00123_),
    .RESETN(net1866),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35946_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04135_),
    .QN(_00126_),
    .RESETN(net1867),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35947_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04136_),
    .QN(_00129_),
    .RESETN(net1868),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35948_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04137_),
    .QN(_00132_),
    .RESETN(net1869),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35949_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04138_),
    .QN(_00135_),
    .RESETN(net1870),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35950_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04139_),
    .QN(_00138_),
    .RESETN(net1871),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _35951_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04140_),
    .QN(_00141_),
    .RESETN(net1872),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35952_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04141_),
    .QN(_00144_),
    .RESETN(net1873),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35953_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04142_),
    .QN(_00147_),
    .RESETN(net1874),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35954_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04143_),
    .QN(_00150_),
    .RESETN(net1875),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _35955_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04144_),
    .QN(_00153_),
    .RESETN(net1876),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35956_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04145_),
    .QN(_00156_),
    .RESETN(net1877),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35957_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04146_),
    .QN(_00159_),
    .RESETN(net1878),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _35958_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04147_),
    .QN(_00161_),
    .RESETN(net1879),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _35959_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04148_),
    .QN(_02066_),
    .RESETN(net1880),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35960_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04149_),
    .QN(_02065_),
    .RESETN(net1881),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35961_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04150_),
    .QN(_02064_),
    .RESETN(net1882),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35962_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04151_),
    .QN(_02063_),
    .RESETN(net1883),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35963_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04152_),
    .QN(_02062_),
    .RESETN(net1884),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35964_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04153_),
    .QN(_02061_),
    .RESETN(net1885),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35965_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04154_),
    .QN(_02060_),
    .RESETN(net1886),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35966_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04155_),
    .QN(_02059_),
    .RESETN(net1887),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35967_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04156_),
    .QN(_02058_),
    .RESETN(net1888),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35968_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04157_),
    .QN(_02057_),
    .RESETN(net1889),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35969_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04158_),
    .QN(_02056_),
    .RESETN(net1890),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35970_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04159_),
    .QN(_02055_),
    .RESETN(net1891),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35971_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04160_),
    .QN(_02054_),
    .RESETN(net1892),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35972_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04161_),
    .QN(_02053_),
    .RESETN(net1893),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35973_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04162_),
    .QN(_02052_),
    .RESETN(net1894),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35974_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04163_),
    .QN(_02051_),
    .RESETN(net1895),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35975_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04164_),
    .QN(_02050_),
    .RESETN(net1896),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35976_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04165_),
    .QN(_02049_),
    .RESETN(net1897),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35977_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04166_),
    .QN(_02048_),
    .RESETN(net1898),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35978_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04167_),
    .QN(_02047_),
    .RESETN(net1899),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35979_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04168_),
    .QN(_02046_),
    .RESETN(net1900),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35980_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04169_),
    .QN(_02045_),
    .RESETN(net1901),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35981_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04170_),
    .QN(_02044_),
    .RESETN(net1902),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35982_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04171_),
    .QN(_02043_),
    .RESETN(net1903),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35983_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04172_),
    .QN(_02042_),
    .RESETN(net1904),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35984_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04173_),
    .QN(_02041_),
    .RESETN(net1905),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35985_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04174_),
    .QN(_02040_),
    .RESETN(net1906),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35986_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04175_),
    .QN(_02039_),
    .RESETN(net1907),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35987_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04176_),
    .QN(_02038_),
    .RESETN(net1908),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35988_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04177_),
    .QN(_02037_),
    .RESETN(net1909),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35989_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_04178_),
    .QN(_02036_),
    .RESETN(net1910),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35990_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_04179_),
    .QN(_02035_),
    .RESETN(net1911),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35991_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04180_),
    .QN(_02034_),
    .RESETN(net1912),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _35992_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04181_),
    .QN(_02033_),
    .RESETN(net1913),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _35993_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04182_),
    .QN(_02032_),
    .RESETN(net1914),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35994_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04183_),
    .QN(_02031_),
    .RESETN(net1915),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _35995_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04184_),
    .QN(_02030_),
    .RESETN(net1916),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _35996_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04185_),
    .QN(_02029_),
    .RESETN(net1917),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35997_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04186_),
    .QN(_02028_),
    .RESETN(net1918),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _35998_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04187_),
    .QN(_02027_),
    .RESETN(net1919),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35999_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04188_),
    .QN(_02026_),
    .RESETN(net1920),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36000_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04189_),
    .QN(_02025_),
    .RESETN(net1921),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36001_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04190_),
    .QN(_02024_),
    .RESETN(net1922),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36002_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04191_),
    .QN(_02023_),
    .RESETN(net1923),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36003_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04192_),
    .QN(_02022_),
    .RESETN(net1924),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36004_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04193_),
    .QN(_02021_),
    .RESETN(net1925),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36005_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04194_),
    .QN(_02020_),
    .RESETN(net1926),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36006_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04195_),
    .QN(_02019_),
    .RESETN(net1927),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36007_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04196_),
    .QN(_02018_),
    .RESETN(net1928),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36008_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04197_),
    .QN(_02017_),
    .RESETN(net1929),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36009_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04198_),
    .QN(_02016_),
    .RESETN(net1930),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36010_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04199_),
    .QN(_02015_),
    .RESETN(net1931),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36011_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04200_),
    .QN(_02014_),
    .RESETN(net1932),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36012_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04201_),
    .QN(_02013_),
    .RESETN(net1933),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36013_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04202_),
    .QN(_02012_),
    .RESETN(net1934),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36014_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04203_),
    .QN(_02011_),
    .RESETN(net1935),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36015_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04204_),
    .QN(_02010_),
    .RESETN(net1936),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36016_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04205_),
    .QN(_02009_),
    .RESETN(net1937),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36017_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04206_),
    .QN(_02008_),
    .RESETN(net1938),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36018_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04207_),
    .QN(_02007_),
    .RESETN(net1939),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36019_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04208_),
    .QN(_02006_),
    .RESETN(net1940),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36020_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04209_),
    .QN(_02005_),
    .RESETN(net1941),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36021_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04210_),
    .QN(_02004_),
    .RESETN(net1942),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36022_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04211_),
    .QN(_02003_),
    .RESETN(net1943),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36023_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04212_),
    .QN(_02002_),
    .RESETN(net1944),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36024_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04213_),
    .QN(_02001_),
    .RESETN(net1945),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36025_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04214_),
    .QN(_02000_),
    .RESETN(net1946),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36026_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04215_),
    .QN(_01999_),
    .RESETN(net1947),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36027_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04216_),
    .QN(_01998_),
    .RESETN(net1948),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36028_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04217_),
    .QN(_01997_),
    .RESETN(net1949),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36029_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04218_),
    .QN(_01996_),
    .RESETN(net1950),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36030_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04219_),
    .QN(_01995_),
    .RESETN(net1951),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36031_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04220_),
    .QN(_01994_),
    .RESETN(net1952),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36032_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04221_),
    .QN(_01993_),
    .RESETN(net1953),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36033_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04222_),
    .QN(_01992_),
    .RESETN(net1954),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36034_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04223_),
    .QN(_01991_),
    .RESETN(net1955),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36035_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04224_),
    .QN(_01990_),
    .RESETN(net1956),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36036_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04225_),
    .QN(_01989_),
    .RESETN(net1957),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36037_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04226_),
    .QN(_01988_),
    .RESETN(net1958),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36038_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04227_),
    .QN(_01987_),
    .RESETN(net1959),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36039_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04228_),
    .QN(_01986_),
    .RESETN(net1960),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36040_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04229_),
    .QN(_01985_),
    .RESETN(net1961),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36041_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04230_),
    .QN(_01984_),
    .RESETN(net1962),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36042_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04231_),
    .QN(_01983_),
    .RESETN(net1963),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36043_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04232_),
    .QN(_01982_),
    .RESETN(net1964),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36044_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04233_),
    .QN(_01981_),
    .RESETN(net1965),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36045_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04234_),
    .QN(_01980_),
    .RESETN(net1966),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36046_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04235_),
    .QN(_01979_),
    .RESETN(net1967),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36047_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04236_),
    .QN(_01978_),
    .RESETN(net1968),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36048_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04237_),
    .QN(_01977_),
    .RESETN(net1969),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36049_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04238_),
    .QN(_01976_),
    .RESETN(net1970),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36050_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04239_),
    .QN(_01975_),
    .RESETN(net1971),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36051_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04240_),
    .QN(_01974_),
    .RESETN(net1972),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36052_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04241_),
    .QN(_01973_),
    .RESETN(net1973),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36053_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04242_),
    .QN(_01972_),
    .RESETN(net1974),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36054_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04243_),
    .QN(_01971_),
    .RESETN(net1975),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36055_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04244_),
    .QN(_01970_),
    .RESETN(net1976),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36056_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04245_),
    .QN(_01969_),
    .RESETN(net1977),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36057_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04246_),
    .QN(_01968_),
    .RESETN(net1978),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36058_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04247_),
    .QN(_01967_),
    .RESETN(net1979),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36059_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04248_),
    .QN(_01966_),
    .RESETN(net1980),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36060_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04249_),
    .QN(_01965_),
    .RESETN(net1981),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36061_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04250_),
    .QN(_01964_),
    .RESETN(net1982),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36062_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04251_),
    .QN(_01963_),
    .RESETN(net1983),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36063_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04252_),
    .QN(_01962_),
    .RESETN(net1984),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36064_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04253_),
    .QN(_01961_),
    .RESETN(net1985),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36065_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04254_),
    .QN(_01960_),
    .RESETN(net1986),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36066_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04255_),
    .QN(_01959_),
    .RESETN(net1987),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36067_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04256_),
    .QN(_01958_),
    .RESETN(net1988),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36068_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04257_),
    .QN(_01957_),
    .RESETN(net1989),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36069_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04258_),
    .QN(_01956_),
    .RESETN(net1990),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36070_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04259_),
    .QN(_01955_),
    .RESETN(net1991),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36071_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04260_),
    .QN(_01954_),
    .RESETN(net1992),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36072_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04261_),
    .QN(_01953_),
    .RESETN(net1993),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36073_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04262_),
    .QN(_01952_),
    .RESETN(net1994),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36074_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04263_),
    .QN(_01951_),
    .RESETN(net1995),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36075_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04264_),
    .QN(_01950_),
    .RESETN(net1996),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36076_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04265_),
    .QN(_01949_),
    .RESETN(net1997),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36077_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04266_),
    .QN(_01948_),
    .RESETN(net1998),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36078_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04267_),
    .QN(_01947_),
    .RESETN(net1999),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36079_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04268_),
    .QN(_01946_),
    .RESETN(net2000),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36080_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04269_),
    .QN(_01945_),
    .RESETN(net2001),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36081_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04270_),
    .QN(_01944_),
    .RESETN(net2002),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36082_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04271_),
    .QN(_01943_),
    .RESETN(net2003),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36083_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04272_),
    .QN(_01942_),
    .RESETN(net2004),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36084_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04273_),
    .QN(_01941_),
    .RESETN(net2005),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36085_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04274_),
    .QN(_01940_),
    .RESETN(net2006),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36086_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04275_),
    .QN(_01939_),
    .RESETN(net2007),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36087_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04276_),
    .QN(_01938_),
    .RESETN(net2008),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36088_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04277_),
    .QN(_01937_),
    .RESETN(net2009),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36089_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04278_),
    .QN(_01936_),
    .RESETN(net2010),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36090_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04279_),
    .QN(_01935_),
    .RESETN(net2011),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36091_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04280_),
    .QN(_01934_),
    .RESETN(net2012),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36092_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04281_),
    .QN(_01933_),
    .RESETN(net2013),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36093_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04282_),
    .QN(_01932_),
    .RESETN(net2014),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36094_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04283_),
    .QN(_01931_),
    .RESETN(net2015),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36095_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04284_),
    .QN(_01930_),
    .RESETN(net2016),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36096_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04285_),
    .QN(_01929_),
    .RESETN(net2017),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36097_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04286_),
    .QN(_01928_),
    .RESETN(net2018),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36098_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04287_),
    .QN(_01927_),
    .RESETN(net2019),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36099_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04288_),
    .QN(_01926_),
    .RESETN(net2020),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36100_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04289_),
    .QN(_01925_),
    .RESETN(net2021),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36101_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04290_),
    .QN(_01924_),
    .RESETN(net2022),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36102_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04291_),
    .QN(_01923_),
    .RESETN(net2023),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36103_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04292_),
    .QN(_01922_),
    .RESETN(net2024),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36104_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04293_),
    .QN(_01921_),
    .RESETN(net2025),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36105_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04294_),
    .QN(_01920_),
    .RESETN(net2026),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36106_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04295_),
    .QN(_01919_),
    .RESETN(net2027),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36107_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04296_),
    .QN(_01918_),
    .RESETN(net2028),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36108_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04297_),
    .QN(_01917_),
    .RESETN(net2029),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36109_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04298_),
    .QN(_01916_),
    .RESETN(net2030),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36110_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04299_),
    .QN(_01915_),
    .RESETN(net2031),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36111_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04300_),
    .QN(_01914_),
    .RESETN(net2032),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36112_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04301_),
    .QN(_01913_),
    .RESETN(net2033),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36113_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04302_),
    .QN(_01912_),
    .RESETN(net2034),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36114_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04303_),
    .QN(_01911_),
    .RESETN(net2035),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36115_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04304_),
    .QN(_01910_),
    .RESETN(net2036),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36116_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04305_),
    .QN(_01909_),
    .RESETN(net2037),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36117_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04306_),
    .QN(_01908_),
    .RESETN(net2038),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36118_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04307_),
    .QN(_01907_),
    .RESETN(net2039),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36119_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04308_),
    .QN(_01906_),
    .RESETN(net2040),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36120_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04309_),
    .QN(_01905_),
    .RESETN(net2041),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36121_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04310_),
    .QN(_01904_),
    .RESETN(net2042),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36122_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04311_),
    .QN(_01903_),
    .RESETN(net2043),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36123_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04312_),
    .QN(_01902_),
    .RESETN(net2044),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36124_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04313_),
    .QN(_01901_),
    .RESETN(net2045),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36125_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04314_),
    .QN(_01900_),
    .RESETN(net2046),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36126_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04315_),
    .QN(_01899_),
    .RESETN(net2047),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36127_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_04316_),
    .QN(_01898_),
    .RESETN(net2048),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36128_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_04317_),
    .QN(_01897_),
    .RESETN(net2049),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36129_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04318_),
    .QN(_01896_),
    .RESETN(net2050),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36130_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_04319_),
    .QN(_01895_),
    .RESETN(net2051),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36131_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04320_),
    .QN(_01894_),
    .RESETN(net2052),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36132_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04321_),
    .QN(_01893_),
    .RESETN(net2053),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36133_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04322_),
    .QN(_01892_),
    .RESETN(net2054),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36134_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04323_),
    .QN(_01891_),
    .RESETN(net2055),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36135_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04324_),
    .QN(_01890_),
    .RESETN(net2056),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36136_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04325_),
    .QN(_01889_),
    .RESETN(net2057),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36137_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04326_),
    .QN(_01888_),
    .RESETN(net2058),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36138_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04327_),
    .QN(_01887_),
    .RESETN(net2059),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36139_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04328_),
    .QN(_01886_),
    .RESETN(net2060),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36140_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04329_),
    .QN(_01885_),
    .RESETN(net2061),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36141_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04330_),
    .QN(_01884_),
    .RESETN(net2062),
    .SETN(net148));
 DFFASRHQNx1_ASAP7_75t_R _36142_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04331_),
    .QN(_01883_),
    .RESETN(net2063),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36143_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04332_),
    .QN(_01882_),
    .RESETN(net2064),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36144_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04333_),
    .QN(_01881_),
    .RESETN(net2065),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36145_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04334_),
    .QN(_01880_),
    .RESETN(net2066),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36146_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04335_),
    .QN(_01879_),
    .RESETN(net2067),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36147_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04336_),
    .QN(_01878_),
    .RESETN(net2068),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36148_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04337_),
    .QN(_01877_),
    .RESETN(net2069),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36149_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04338_),
    .QN(_01876_),
    .RESETN(net2070),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36150_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04339_),
    .QN(_00661_),
    .RESETN(net2071),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36151_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04340_),
    .QN(_01315_),
    .RESETN(net2072),
    .SETN(net434));
 DFFASRHQNx1_ASAP7_75t_R _36152_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_04341_),
    .QN(_01875_),
    .RESETN(net2073),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _36153_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_04342_),
    .QN(_01874_),
    .RESETN(net2074),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _36154_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_04343_),
    .QN(_00285_),
    .RESETN(net2075),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _36155_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_04344_),
    .QN(_01873_),
    .RESETN(net2076),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _36156_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_04345_),
    .QN(_01872_),
    .RESETN(net443),
    .SETN(net2077));
 DFFASRHQNx1_ASAP7_75t_R _36157_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04346_),
    .QN(_01871_),
    .RESETN(net2078),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36158_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04347_),
    .QN(_01870_),
    .RESETN(net2079),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36159_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04348_),
    .QN(_01869_),
    .RESETN(net2080),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36160_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04349_),
    .QN(_01868_),
    .RESETN(net2081),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36161_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04350_),
    .QN(_01867_),
    .RESETN(net2082),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36162_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04351_),
    .QN(_01866_),
    .RESETN(net2083),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36163_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04352_),
    .QN(_01865_),
    .RESETN(net2084),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36164_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04353_),
    .QN(_01864_),
    .RESETN(net2085),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36165_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04354_),
    .QN(_01863_),
    .RESETN(net2086),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36166_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04355_),
    .QN(_01862_),
    .RESETN(net2087),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _36167_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04356_),
    .QN(_01861_),
    .RESETN(net2088),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36168_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04357_),
    .QN(_01860_),
    .RESETN(net2089),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36169_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04358_),
    .QN(_01859_),
    .RESETN(net2090),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36170_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04359_),
    .QN(_01858_),
    .RESETN(net2091),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36171_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04360_),
    .QN(_01857_),
    .RESETN(net2092),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36172_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04361_),
    .QN(_01856_),
    .RESETN(net2093),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36173_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04362_),
    .QN(_01855_),
    .RESETN(net2094),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36174_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04363_),
    .QN(_01854_),
    .RESETN(net2095),
    .SETN(net433));
 DFFASRHQNx1_ASAP7_75t_R _36175_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04364_),
    .QN(_01853_),
    .RESETN(net2096),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36176_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04365_),
    .QN(_01852_),
    .RESETN(net2097),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36177_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04366_),
    .QN(_01851_),
    .RESETN(net2098),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36178_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04367_),
    .QN(_01850_),
    .RESETN(net2099),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36179_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04368_),
    .QN(_01849_),
    .RESETN(net2100),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36180_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04369_),
    .QN(_01733_),
    .RESETN(net2101),
    .SETN(net432));
 DFFASRHQNx1_ASAP7_75t_R _36181_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(core_busy_d),
    .QN(_01734_),
    .RESETN(net2102),
    .SETN(net437));
 DLLx1_ASAP7_75t_R _36182_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_00008_),
    .Q(\core_clock_gate_i.en_latch ));
 DFFASRHQNx1_ASAP7_75t_R _36183_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ),
    .QN(_00237_),
    .RESETN(net2103),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36184_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .QN(_01735_),
    .RESETN(net2104),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36185_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ),
    .QN(_01736_),
    .RESETN(net2105),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36186_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ),
    .QN(_00238_),
    .RESETN(net2106),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36187_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ),
    .QN(_01737_),
    .RESETN(net2107),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36188_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ),
    .QN(_01848_),
    .RESETN(net2108),
    .SETN(net437));
 DFFHQNx1_ASAP7_75t_R _36189_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04370_),
    .QN(_01847_));
 DFFHQNx1_ASAP7_75t_R _36190_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04371_),
    .QN(_01846_));
 DFFHQNx1_ASAP7_75t_R _36191_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04372_),
    .QN(_01845_));
 DFFHQNx1_ASAP7_75t_R _36192_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04373_),
    .QN(_01844_));
 DFFHQNx1_ASAP7_75t_R _36193_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04374_),
    .QN(_01843_));
 DFFHQNx1_ASAP7_75t_R _36194_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04375_),
    .QN(_01842_));
 DFFHQNx1_ASAP7_75t_R _36195_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04376_),
    .QN(_01841_));
 DFFHQNx1_ASAP7_75t_R _36196_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04377_),
    .QN(_01840_));
 DFFHQNx1_ASAP7_75t_R _36197_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04378_),
    .QN(_01839_));
 DFFHQNx1_ASAP7_75t_R _36198_ (.CLK(\clknet_leaf_31_core_clock_gate_i.clk_o ),
    .D(_04379_),
    .QN(_01838_));
 DFFHQNx1_ASAP7_75t_R _36199_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04380_),
    .QN(_01837_));
 DFFHQNx1_ASAP7_75t_R _36200_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04381_),
    .QN(_01836_));
 DFFHQNx1_ASAP7_75t_R _36201_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04382_),
    .QN(_01835_));
 DFFHQNx1_ASAP7_75t_R _36202_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04383_),
    .QN(_01834_));
 DFFHQNx1_ASAP7_75t_R _36203_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04384_),
    .QN(_01833_));
 DFFHQNx1_ASAP7_75t_R _36204_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04385_),
    .QN(_01832_));
 DFFHQNx1_ASAP7_75t_R _36205_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04386_),
    .QN(_01831_));
 DFFHQNx1_ASAP7_75t_R _36206_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04387_),
    .QN(_01830_));
 DFFHQNx1_ASAP7_75t_R _36207_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04388_),
    .QN(_01829_));
 DFFHQNx1_ASAP7_75t_R _36208_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04389_),
    .QN(_01828_));
 DFFHQNx1_ASAP7_75t_R _36209_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04390_),
    .QN(_01827_));
 DFFHQNx1_ASAP7_75t_R _36210_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04391_),
    .QN(_01826_));
 DFFHQNx1_ASAP7_75t_R _36211_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04392_),
    .QN(_01825_));
 DFFHQNx1_ASAP7_75t_R _36212_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04393_),
    .QN(_01824_));
 DFFHQNx1_ASAP7_75t_R _36213_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04394_),
    .QN(_01823_));
 DFFHQNx1_ASAP7_75t_R _36214_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04395_),
    .QN(_01822_));
 DFFHQNx1_ASAP7_75t_R _36215_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04396_),
    .QN(_01821_));
 DFFHQNx1_ASAP7_75t_R _36216_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04397_),
    .QN(_01820_));
 DFFHQNx1_ASAP7_75t_R _36217_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04398_),
    .QN(_01819_));
 DFFHQNx1_ASAP7_75t_R _36218_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04399_),
    .QN(_01818_));
 DFFHQNx1_ASAP7_75t_R _36219_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04400_),
    .QN(_01817_));
 DFFHQNx1_ASAP7_75t_R _36220_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04401_),
    .QN(_01816_));
 DFFHQNx1_ASAP7_75t_R _36221_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04402_),
    .QN(_01738_));
 DFFASRHQNx1_ASAP7_75t_R _36222_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ),
    .QN(_00240_),
    .RESETN(net2109),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36223_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ),
    .QN(_00239_),
    .RESETN(net2110),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36224_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ),
    .QN(_01815_),
    .RESETN(net2111),
    .SETN(net437));
 DFFHQNx1_ASAP7_75t_R _36225_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04403_),
    .QN(_01814_));
 DFFHQNx1_ASAP7_75t_R _36226_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04404_),
    .QN(_01813_));
 DFFHQNx1_ASAP7_75t_R _36227_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04405_),
    .QN(_01812_));
 DFFHQNx1_ASAP7_75t_R _36228_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04406_),
    .QN(_01811_));
 DFFHQNx1_ASAP7_75t_R _36229_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04407_),
    .QN(_01810_));
 DFFHQNx1_ASAP7_75t_R _36230_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04408_),
    .QN(_01809_));
 DFFHQNx1_ASAP7_75t_R _36231_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04409_),
    .QN(_01808_));
 DFFHQNx1_ASAP7_75t_R _36232_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04410_),
    .QN(_01807_));
 DFFHQNx1_ASAP7_75t_R _36233_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04411_),
    .QN(_01806_));
 DFFHQNx1_ASAP7_75t_R _36234_ (.CLK(\clknet_leaf_31_core_clock_gate_i.clk_o ),
    .D(_04412_),
    .QN(_01805_));
 DFFHQNx1_ASAP7_75t_R _36235_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04413_),
    .QN(_01804_));
 DFFHQNx1_ASAP7_75t_R _36236_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04414_),
    .QN(_01803_));
 DFFHQNx1_ASAP7_75t_R _36237_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04415_),
    .QN(_01802_));
 DFFHQNx1_ASAP7_75t_R _36238_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04416_),
    .QN(_01801_));
 DFFHQNx1_ASAP7_75t_R _36239_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04417_),
    .QN(_01800_));
 DFFHQNx1_ASAP7_75t_R _36240_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04418_),
    .QN(_01799_));
 DFFHQNx1_ASAP7_75t_R _36241_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04419_),
    .QN(_01798_));
 DFFHQNx1_ASAP7_75t_R _36242_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04420_),
    .QN(_01797_));
 DFFHQNx1_ASAP7_75t_R _36243_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04421_),
    .QN(_01796_));
 DFFHQNx1_ASAP7_75t_R _36244_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04422_),
    .QN(_01795_));
 DFFHQNx1_ASAP7_75t_R _36245_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04423_),
    .QN(_01794_));
 DFFHQNx1_ASAP7_75t_R _36246_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04424_),
    .QN(_01793_));
 DFFHQNx1_ASAP7_75t_R _36247_ (.CLK(\clknet_leaf_31_core_clock_gate_i.clk_o ),
    .D(_04425_),
    .QN(_01792_));
 DFFHQNx1_ASAP7_75t_R _36248_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04426_),
    .QN(_01791_));
 DFFHQNx1_ASAP7_75t_R _36249_ (.CLK(\clknet_leaf_31_core_clock_gate_i.clk_o ),
    .D(_04427_),
    .QN(_01790_));
 DFFHQNx1_ASAP7_75t_R _36250_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04428_),
    .QN(_01789_));
 DFFHQNx1_ASAP7_75t_R _36251_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04429_),
    .QN(_01788_));
 DFFHQNx1_ASAP7_75t_R _36252_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04430_),
    .QN(_01787_));
 DFFHQNx1_ASAP7_75t_R _36253_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04431_),
    .QN(_01786_));
 DFFHQNx1_ASAP7_75t_R _36254_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04432_),
    .QN(_01785_));
 DFFHQNx1_ASAP7_75t_R _36255_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04433_),
    .QN(_01784_));
 DFFHQNx1_ASAP7_75t_R _36256_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04434_),
    .QN(_01783_));
 DFFHQNx1_ASAP7_75t_R _36257_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04435_),
    .QN(_01782_));
 DFFHQNx1_ASAP7_75t_R _36258_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04436_),
    .QN(_01781_));
 DFFHQNx1_ASAP7_75t_R _36259_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04437_),
    .QN(_01780_));
 DFFHQNx1_ASAP7_75t_R _36260_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04438_),
    .QN(_01779_));
 DFFHQNx1_ASAP7_75t_R _36261_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04439_),
    .QN(_01778_));
 DFFHQNx1_ASAP7_75t_R _36262_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04440_),
    .QN(_01777_));
 DFFHQNx1_ASAP7_75t_R _36263_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04441_),
    .QN(_01776_));
 DFFHQNx1_ASAP7_75t_R _36264_ (.CLK(\clknet_leaf_31_core_clock_gate_i.clk_o ),
    .D(_04442_),
    .QN(_01775_));
 DFFHQNx1_ASAP7_75t_R _36265_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04443_),
    .QN(_01774_));
 DFFHQNx1_ASAP7_75t_R _36266_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04444_),
    .QN(_01773_));
 DFFHQNx1_ASAP7_75t_R _36267_ (.CLK(\clknet_leaf_31_core_clock_gate_i.clk_o ),
    .D(_04445_),
    .QN(_01772_));
 DFFHQNx1_ASAP7_75t_R _36268_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04446_),
    .QN(_01771_));
 DFFHQNx1_ASAP7_75t_R _36269_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04447_),
    .QN(_01770_));
 DFFHQNx1_ASAP7_75t_R _36270_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04448_),
    .QN(_01769_));
 DFFHQNx1_ASAP7_75t_R _36271_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04449_),
    .QN(_01768_));
 DFFHQNx1_ASAP7_75t_R _36272_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04450_),
    .QN(_01767_));
 DFFHQNx1_ASAP7_75t_R _36273_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04451_),
    .QN(_01766_));
 DFFHQNx1_ASAP7_75t_R _36274_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04452_),
    .QN(_01765_));
 DFFHQNx1_ASAP7_75t_R _36275_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04453_),
    .QN(_01764_));
 DFFHQNx1_ASAP7_75t_R _36276_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04454_),
    .QN(_01763_));
 DFFHQNx1_ASAP7_75t_R _36277_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04455_),
    .QN(_01762_));
 DFFHQNx1_ASAP7_75t_R _36278_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04456_),
    .QN(_01761_));
 DFFHQNx1_ASAP7_75t_R _36279_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04457_),
    .QN(_01760_));
 DFFHQNx1_ASAP7_75t_R _36280_ (.CLK(\clknet_leaf_31_core_clock_gate_i.clk_o ),
    .D(_04458_),
    .QN(_01759_));
 DFFHQNx1_ASAP7_75t_R _36281_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04459_),
    .QN(_01758_));
 DFFHQNx1_ASAP7_75t_R _36282_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04460_),
    .QN(_01757_));
 DFFHQNx1_ASAP7_75t_R _36283_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04461_),
    .QN(_01756_));
 DFFHQNx1_ASAP7_75t_R _36284_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04462_),
    .QN(_01755_));
 DFFHQNx1_ASAP7_75t_R _36285_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04463_),
    .QN(_01754_));
 DFFHQNx1_ASAP7_75t_R _36286_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04464_),
    .QN(_01753_));
 DFFHQNx1_ASAP7_75t_R _36287_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04465_),
    .QN(_01752_));
 DFFHQNx1_ASAP7_75t_R _36288_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04466_),
    .QN(_01751_));
 DFFHQNx1_ASAP7_75t_R _36289_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04467_),
    .QN(_01750_));
 DFFHQNx1_ASAP7_75t_R _36290_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04468_),
    .QN(_01749_));
 DFFHQNx1_ASAP7_75t_R _36291_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04469_),
    .QN(_01748_));
 DFFASRHQNx1_ASAP7_75t_R _36292_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_04470_),
    .QN(_01747_),
    .RESETN(net2112),
    .SETN(net437));
 DFFHQNx1_ASAP7_75t_R _36293_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04471_),
    .QN(_01746_));
 DFFHQNx1_ASAP7_75t_R _36294_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04472_),
    .QN(_00163_));
 DFFHQNx1_ASAP7_75t_R _36295_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04473_),
    .QN(_00165_));
 DFFHQNx1_ASAP7_75t_R _36296_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04474_),
    .QN(_00168_));
 DFFHQNx1_ASAP7_75t_R _36297_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04475_),
    .QN(_00172_));
 DFFHQNx1_ASAP7_75t_R _36298_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04476_),
    .QN(_00175_));
 DFFHQNx1_ASAP7_75t_R _36299_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04477_),
    .QN(_00278_));
 DFFHQNx1_ASAP7_75t_R _36300_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04478_),
    .QN(_00323_));
 DFFHQNx1_ASAP7_75t_R _36301_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04479_),
    .QN(_00184_));
 DFFHQNx1_ASAP7_75t_R _36302_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04480_),
    .QN(_00187_));
 DFFHQNx1_ASAP7_75t_R _36303_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04481_),
    .QN(_00191_));
 DFFHQNx1_ASAP7_75t_R _36304_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04482_),
    .QN(_00194_));
 DFFHQNx1_ASAP7_75t_R _36305_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04483_),
    .QN(_00281_));
 DFFHQNx1_ASAP7_75t_R _36306_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04484_),
    .QN(_00282_));
 DFFHQNx1_ASAP7_75t_R _36307_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04485_),
    .QN(_00279_));
 DFFHQNx1_ASAP7_75t_R _36308_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04486_),
    .QN(_00290_));
 DFFHQNx1_ASAP7_75t_R _36309_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04487_),
    .QN(_00289_));
 DFFHQNx1_ASAP7_75t_R _36310_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04488_),
    .QN(_00288_));
 DFFHQNx1_ASAP7_75t_R _36311_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04489_),
    .QN(_00287_));
 DFFHQNx1_ASAP7_75t_R _36312_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04490_),
    .QN(_00286_));
 DFFHQNx1_ASAP7_75t_R _36313_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04491_),
    .QN(_00246_));
 DFFHQNx1_ASAP7_75t_R _36314_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04492_),
    .QN(_01745_));
 DFFHQNx1_ASAP7_75t_R _36315_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04493_),
    .QN(_01744_));
 DFFHQNx1_ASAP7_75t_R _36316_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04494_),
    .QN(_00245_));
 DFFHQNx1_ASAP7_75t_R _36317_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04495_),
    .QN(_00244_));
 DFFHQNx1_ASAP7_75t_R _36318_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04496_),
    .QN(_01743_));
 DFFHQNx1_ASAP7_75t_R _36319_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04497_),
    .QN(_00283_));
 DFFHQNx1_ASAP7_75t_R _36320_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04498_),
    .QN(_01742_));
 DFFHQNx1_ASAP7_75t_R _36321_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04499_),
    .QN(_01741_));
 DFFHQNx1_ASAP7_75t_R _36322_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04500_),
    .QN(_01740_));
 DFFHQNx1_ASAP7_75t_R _36323_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04501_),
    .QN(_01739_));
 DFFHQNx1_ASAP7_75t_R _36324_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04502_),
    .QN(_00280_));
 DFFASRHQNx1_ASAP7_75t_R _36325_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04503_),
    .QN(_01311_),
    .RESETN(net2113),
    .SETN(net435));
 BUFx4_ASAP7_75t_R clkbuf_leaf_0_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_0_clk_i));
 TIEHIx1_ASAP7_75t_R _34444__456 (.H(net456));
 TAPCELL_ASAP7_75t_R PHY_30 ();
 BUFx2_ASAP7_75t_R _36329_ (.A(net451),
    .Y(alert_minor_o));
 BUFx2_ASAP7_75t_R _36330_ (.A(net452),
    .Y(data_addr_o[0]));
 BUFx2_ASAP7_75t_R _36331_ (.A(net453),
    .Y(data_addr_o[1]));
 TAPCELL_ASAP7_75t_R PHY_29 ();
 TAPCELL_ASAP7_75t_R PHY_28 ();
 TAPCELL_ASAP7_75t_R PHY_27 ();
 TAPCELL_ASAP7_75t_R PHY_26 ();
 TAPCELL_ASAP7_75t_R PHY_25 ();
 TAPCELL_ASAP7_75t_R PHY_24 ();
 TAPCELL_ASAP7_75t_R PHY_23 ();
 TAPCELL_ASAP7_75t_R PHY_22 ();
 TAPCELL_ASAP7_75t_R PHY_21 ();
 TAPCELL_ASAP7_75t_R PHY_20 ();
 TAPCELL_ASAP7_75t_R PHY_19 ();
 TAPCELL_ASAP7_75t_R PHY_18 ();
 TAPCELL_ASAP7_75t_R PHY_17 ();
 TAPCELL_ASAP7_75t_R PHY_16 ();
 TAPCELL_ASAP7_75t_R PHY_15 ();
 TAPCELL_ASAP7_75t_R PHY_14 ();
 TAPCELL_ASAP7_75t_R PHY_13 ();
 TAPCELL_ASAP7_75t_R PHY_12 ();
 TAPCELL_ASAP7_75t_R PHY_11 ();
 TAPCELL_ASAP7_75t_R PHY_10 ();
 TAPCELL_ASAP7_75t_R PHY_9 ();
 TAPCELL_ASAP7_75t_R PHY_8 ();
 TAPCELL_ASAP7_75t_R PHY_7 ();
 TAPCELL_ASAP7_75t_R PHY_6 ();
 TAPCELL_ASAP7_75t_R PHY_5 ();
 TAPCELL_ASAP7_75t_R PHY_4 ();
 TAPCELL_ASAP7_75t_R PHY_3 ();
 TAPCELL_ASAP7_75t_R PHY_2 ();
 TAPCELL_ASAP7_75t_R PHY_1 ();
 TAPCELL_ASAP7_75t_R PHY_0 ();
 BUFx2_ASAP7_75t_R _36362_ (.A(net454),
    .Y(instr_addr_o[0]));
 BUFx2_ASAP7_75t_R _36363_ (.A(net455),
    .Y(instr_addr_o[1]));
 TIEHIx1_ASAP7_75t_R _34857__808 (.H(net808));
 TIEHIx1_ASAP7_75t_R _34858__809 (.H(net809));
 TIEHIx1_ASAP7_75t_R _34859__810 (.H(net810));
 TIEHIx1_ASAP7_75t_R _34860__811 (.H(net811));
 TIEHIx1_ASAP7_75t_R _34861__812 (.H(net812));
 TIEHIx1_ASAP7_75t_R _34862__813 (.H(net813));
 TIEHIx1_ASAP7_75t_R _34863__814 (.H(net814));
 TIEHIx1_ASAP7_75t_R _34864__815 (.H(net815));
 TIEHIx1_ASAP7_75t_R _34865__816 (.H(net816));
 TIEHIx1_ASAP7_75t_R _34866__817 (.H(net817));
 TIEHIx1_ASAP7_75t_R _34867__818 (.H(net818));
 TIEHIx1_ASAP7_75t_R _34868__819 (.H(net819));
 TIEHIx1_ASAP7_75t_R _34869__820 (.H(net820));
 TIEHIx1_ASAP7_75t_R _34870__821 (.H(net821));
 TIEHIx1_ASAP7_75t_R _34871__822 (.H(net822));
 TIEHIx1_ASAP7_75t_R _34872__823 (.H(net823));
 TIEHIx1_ASAP7_75t_R _34873__824 (.H(net824));
 TIEHIx1_ASAP7_75t_R _34874__825 (.H(net825));
 TIEHIx1_ASAP7_75t_R _34875__826 (.H(net826));
 TIEHIx1_ASAP7_75t_R _34876__827 (.H(net827));
 TIEHIx1_ASAP7_75t_R _34877__828 (.H(net828));
 TIEHIx1_ASAP7_75t_R _34878__829 (.H(net829));
 TIEHIx1_ASAP7_75t_R _34879__830 (.H(net830));
 TIEHIx1_ASAP7_75t_R _34880__831 (.H(net831));
 TIEHIx1_ASAP7_75t_R _34881__832 (.H(net832));
 TIEHIx1_ASAP7_75t_R _34882__833 (.H(net833));
 TIEHIx1_ASAP7_75t_R _34883__834 (.H(net834));
 TIEHIx1_ASAP7_75t_R _34884__835 (.H(net835));
 TIEHIx1_ASAP7_75t_R _34885__836 (.H(net836));
 TIEHIx1_ASAP7_75t_R _34886__837 (.H(net837));
 TIEHIx1_ASAP7_75t_R _34887__838 (.H(net838));
 TIEHIx1_ASAP7_75t_R _34888__839 (.H(net839));
 TIEHIx1_ASAP7_75t_R _34889__840 (.H(net840));
 TIEHIx1_ASAP7_75t_R _34890__841 (.H(net841));
 TIEHIx1_ASAP7_75t_R _34891__842 (.H(net842));
 TIEHIx1_ASAP7_75t_R _34892__843 (.H(net843));
 TIEHIx1_ASAP7_75t_R _34893__844 (.H(net844));
 TIEHIx1_ASAP7_75t_R _34894__845 (.H(net845));
 TIEHIx1_ASAP7_75t_R _34895__846 (.H(net846));
 TIEHIx1_ASAP7_75t_R _34896__847 (.H(net847));
 TIEHIx1_ASAP7_75t_R _34897__848 (.H(net848));
 TIEHIx1_ASAP7_75t_R _34898__849 (.H(net849));
 TIEHIx1_ASAP7_75t_R _34899__850 (.H(net850));
 TIEHIx1_ASAP7_75t_R _34900__851 (.H(net851));
 TIEHIx1_ASAP7_75t_R _34901__852 (.H(net852));
 TIEHIx1_ASAP7_75t_R _34902__853 (.H(net853));
 TIEHIx1_ASAP7_75t_R _34903__854 (.H(net854));
 TIEHIx1_ASAP7_75t_R _34904__855 (.H(net855));
 TIEHIx1_ASAP7_75t_R _34905__856 (.H(net856));
 TIEHIx1_ASAP7_75t_R _34906__857 (.H(net857));
 TIEHIx1_ASAP7_75t_R _34907__858 (.H(net858));
 TIEHIx1_ASAP7_75t_R _34908__859 (.H(net859));
 TIEHIx1_ASAP7_75t_R _34909__860 (.H(net860));
 TIEHIx1_ASAP7_75t_R _34910__861 (.H(net861));
 TIEHIx1_ASAP7_75t_R _34911__862 (.H(net862));
 TIEHIx1_ASAP7_75t_R _34912__863 (.H(net863));
 TIEHIx1_ASAP7_75t_R _34913__864 (.H(net864));
 TIEHIx1_ASAP7_75t_R _34914__865 (.H(net865));
 TIEHIx1_ASAP7_75t_R _34915__866 (.H(net866));
 TIEHIx1_ASAP7_75t_R _34916__867 (.H(net867));
 TIEHIx1_ASAP7_75t_R _34917__868 (.H(net868));
 TIEHIx1_ASAP7_75t_R _34918__869 (.H(net869));
 TIEHIx1_ASAP7_75t_R _34919__870 (.H(net870));
 TIEHIx1_ASAP7_75t_R _34920__871 (.H(net871));
 TIEHIx1_ASAP7_75t_R _34921__872 (.H(net872));
 TIEHIx1_ASAP7_75t_R _34922__873 (.H(net873));
 TIEHIx1_ASAP7_75t_R _34923__874 (.H(net874));
 TIEHIx1_ASAP7_75t_R _34924__875 (.H(net875));
 TIEHIx1_ASAP7_75t_R _34925__876 (.H(net876));
 TIEHIx1_ASAP7_75t_R _34926__877 (.H(net877));
 TIEHIx1_ASAP7_75t_R _34927__878 (.H(net878));
 TIEHIx1_ASAP7_75t_R _34928__879 (.H(net879));
 TIEHIx1_ASAP7_75t_R _34929__880 (.H(net880));
 TIEHIx1_ASAP7_75t_R _34930__881 (.H(net881));
 TIEHIx1_ASAP7_75t_R _34931__882 (.H(net882));
 TIEHIx1_ASAP7_75t_R _34932__883 (.H(net883));
 TIEHIx1_ASAP7_75t_R _34933__884 (.H(net884));
 TIEHIx1_ASAP7_75t_R _34934__885 (.H(net885));
 TIEHIx1_ASAP7_75t_R _34935__886 (.H(net886));
 TIEHIx1_ASAP7_75t_R _34936__887 (.H(net887));
 TIEHIx1_ASAP7_75t_R _34937__888 (.H(net888));
 TIEHIx1_ASAP7_75t_R _34938__889 (.H(net889));
 TIEHIx1_ASAP7_75t_R _34939__890 (.H(net890));
 TIEHIx1_ASAP7_75t_R _34940__891 (.H(net891));
 TIEHIx1_ASAP7_75t_R _34941__892 (.H(net892));
 TIEHIx1_ASAP7_75t_R _34942__893 (.H(net893));
 TIEHIx1_ASAP7_75t_R _34943__894 (.H(net894));
 TIEHIx1_ASAP7_75t_R _34944__895 (.H(net895));
 TIEHIx1_ASAP7_75t_R _34945__896 (.H(net896));
 TIEHIx1_ASAP7_75t_R _34946__897 (.H(net897));
 TIEHIx1_ASAP7_75t_R _34947__898 (.H(net898));
 TIEHIx1_ASAP7_75t_R _34948__899 (.H(net899));
 TIEHIx1_ASAP7_75t_R _34949__900 (.H(net900));
 TIEHIx1_ASAP7_75t_R _34950__901 (.H(net901));
 TIEHIx1_ASAP7_75t_R _34951__902 (.H(net902));
 TIEHIx1_ASAP7_75t_R _34952__903 (.H(net903));
 TIEHIx1_ASAP7_75t_R _34953__904 (.H(net904));
 TIEHIx1_ASAP7_75t_R _34954__905 (.H(net905));
 TIEHIx1_ASAP7_75t_R _34955__906 (.H(net906));
 TIEHIx1_ASAP7_75t_R _34956__907 (.H(net907));
 TIEHIx1_ASAP7_75t_R _34957__908 (.H(net908));
 TIEHIx1_ASAP7_75t_R _34958__909 (.H(net909));
 TIEHIx1_ASAP7_75t_R _34959__910 (.H(net910));
 TIEHIx1_ASAP7_75t_R _34960__911 (.H(net911));
 TIEHIx1_ASAP7_75t_R _34961__912 (.H(net912));
 TIEHIx1_ASAP7_75t_R _34962__913 (.H(net913));
 TIEHIx1_ASAP7_75t_R _34963__914 (.H(net914));
 TIEHIx1_ASAP7_75t_R _34964__915 (.H(net915));
 TIEHIx1_ASAP7_75t_R _34965__916 (.H(net916));
 TIEHIx1_ASAP7_75t_R _34966__917 (.H(net917));
 TIEHIx1_ASAP7_75t_R _34967__918 (.H(net918));
 TIEHIx1_ASAP7_75t_R _34968__919 (.H(net919));
 TIEHIx1_ASAP7_75t_R _34969__920 (.H(net920));
 TIEHIx1_ASAP7_75t_R _34970__921 (.H(net921));
 TIEHIx1_ASAP7_75t_R _34971__922 (.H(net922));
 TIEHIx1_ASAP7_75t_R _34972__923 (.H(net923));
 TIEHIx1_ASAP7_75t_R _34973__924 (.H(net924));
 TIEHIx1_ASAP7_75t_R _34974__925 (.H(net925));
 TIEHIx1_ASAP7_75t_R _34975__926 (.H(net926));
 TIEHIx1_ASAP7_75t_R _34976__927 (.H(net927));
 TIEHIx1_ASAP7_75t_R _34977__928 (.H(net928));
 TIEHIx1_ASAP7_75t_R _34978__929 (.H(net929));
 TIEHIx1_ASAP7_75t_R _34979__930 (.H(net930));
 TIEHIx1_ASAP7_75t_R _34980__931 (.H(net931));
 TIEHIx1_ASAP7_75t_R _34981__932 (.H(net932));
 TIEHIx1_ASAP7_75t_R _34982__933 (.H(net933));
 TIEHIx1_ASAP7_75t_R _34983__934 (.H(net934));
 TIEHIx1_ASAP7_75t_R _34984__935 (.H(net935));
 TIEHIx1_ASAP7_75t_R _34985__936 (.H(net936));
 TIEHIx1_ASAP7_75t_R _34986__937 (.H(net937));
 TIEHIx1_ASAP7_75t_R _34987__938 (.H(net938));
 TIEHIx1_ASAP7_75t_R _34988__939 (.H(net939));
 TIEHIx1_ASAP7_75t_R _34989__940 (.H(net940));
 TIEHIx1_ASAP7_75t_R _34990__941 (.H(net941));
 TIEHIx1_ASAP7_75t_R _34991__942 (.H(net942));
 TIEHIx1_ASAP7_75t_R _34992__943 (.H(net943));
 TIEHIx1_ASAP7_75t_R _34993__944 (.H(net944));
 TIEHIx1_ASAP7_75t_R _34994__945 (.H(net945));
 TIEHIx1_ASAP7_75t_R _34995__946 (.H(net946));
 TIEHIx1_ASAP7_75t_R _34996__947 (.H(net947));
 TIEHIx1_ASAP7_75t_R _34997__948 (.H(net948));
 TIEHIx1_ASAP7_75t_R _34998__949 (.H(net949));
 TIEHIx1_ASAP7_75t_R _34999__950 (.H(net950));
 TIEHIx1_ASAP7_75t_R _35000__951 (.H(net951));
 TIEHIx1_ASAP7_75t_R _35001__952 (.H(net952));
 TIEHIx1_ASAP7_75t_R _35002__953 (.H(net953));
 TIEHIx1_ASAP7_75t_R _35003__954 (.H(net954));
 TIEHIx1_ASAP7_75t_R _35004__955 (.H(net955));
 TIEHIx1_ASAP7_75t_R _35005__956 (.H(net956));
 TIEHIx1_ASAP7_75t_R _35006__957 (.H(net957));
 TIEHIx1_ASAP7_75t_R _35007__958 (.H(net958));
 TIEHIx1_ASAP7_75t_R _35008__959 (.H(net959));
 TIEHIx1_ASAP7_75t_R _35009__960 (.H(net960));
 TIEHIx1_ASAP7_75t_R _35010__961 (.H(net961));
 TIEHIx1_ASAP7_75t_R _35011__962 (.H(net962));
 TIEHIx1_ASAP7_75t_R _35012__963 (.H(net963));
 TIEHIx1_ASAP7_75t_R _35013__964 (.H(net964));
 TIEHIx1_ASAP7_75t_R _35014__965 (.H(net965));
 TIEHIx1_ASAP7_75t_R _35015__966 (.H(net966));
 TIEHIx1_ASAP7_75t_R _35016__967 (.H(net967));
 TIEHIx1_ASAP7_75t_R _35017__968 (.H(net968));
 TIEHIx1_ASAP7_75t_R _35018__969 (.H(net969));
 TIEHIx1_ASAP7_75t_R _35019__970 (.H(net970));
 TIEHIx1_ASAP7_75t_R _35020__971 (.H(net971));
 TIEHIx1_ASAP7_75t_R _35021__972 (.H(net972));
 TIEHIx1_ASAP7_75t_R _35022__973 (.H(net973));
 TIEHIx1_ASAP7_75t_R _35023__974 (.H(net974));
 TIEHIx1_ASAP7_75t_R _35024__975 (.H(net975));
 TIEHIx1_ASAP7_75t_R _35025__976 (.H(net976));
 TIEHIx1_ASAP7_75t_R _35026__977 (.H(net977));
 TIEHIx1_ASAP7_75t_R _35027__978 (.H(net978));
 TIEHIx1_ASAP7_75t_R _35028__979 (.H(net979));
 TIEHIx1_ASAP7_75t_R _35029__980 (.H(net980));
 TIEHIx1_ASAP7_75t_R _35030__981 (.H(net981));
 TIEHIx1_ASAP7_75t_R _35031__982 (.H(net982));
 TIEHIx1_ASAP7_75t_R _35032__983 (.H(net983));
 TIEHIx1_ASAP7_75t_R _35033__984 (.H(net984));
 TIEHIx1_ASAP7_75t_R _35034__985 (.H(net985));
 TIEHIx1_ASAP7_75t_R _35035__986 (.H(net986));
 TIEHIx1_ASAP7_75t_R _35036__987 (.H(net987));
 TIEHIx1_ASAP7_75t_R _35037__988 (.H(net988));
 TIEHIx1_ASAP7_75t_R _35038__989 (.H(net989));
 TIEHIx1_ASAP7_75t_R _35039__990 (.H(net990));
 TIEHIx1_ASAP7_75t_R _35040__991 (.H(net991));
 TIEHIx1_ASAP7_75t_R _35041__992 (.H(net992));
 TIEHIx1_ASAP7_75t_R _35042__993 (.H(net993));
 TIEHIx1_ASAP7_75t_R _35043__994 (.H(net994));
 TIEHIx1_ASAP7_75t_R _35044__995 (.H(net995));
 TIEHIx1_ASAP7_75t_R _35045__996 (.H(net996));
 TIEHIx1_ASAP7_75t_R _35046__997 (.H(net997));
 TIEHIx1_ASAP7_75t_R _35047__998 (.H(net998));
 TIEHIx1_ASAP7_75t_R _35048__999 (.H(net999));
 TIEHIx1_ASAP7_75t_R _35049__1000 (.H(net1000));
 TIEHIx1_ASAP7_75t_R _35050__1001 (.H(net1001));
 TIEHIx1_ASAP7_75t_R _35051__1002 (.H(net1002));
 TIEHIx1_ASAP7_75t_R _35052__1003 (.H(net1003));
 TIEHIx1_ASAP7_75t_R _35053__1004 (.H(net1004));
 TIEHIx1_ASAP7_75t_R _35054__1005 (.H(net1005));
 TIEHIx1_ASAP7_75t_R _35055__1006 (.H(net1006));
 TIEHIx1_ASAP7_75t_R _35056__1007 (.H(net1007));
 TIEHIx1_ASAP7_75t_R _35057__1008 (.H(net1008));
 TIEHIx1_ASAP7_75t_R _35058__1009 (.H(net1009));
 TIEHIx1_ASAP7_75t_R _35059__1010 (.H(net1010));
 TIEHIx1_ASAP7_75t_R _35060__1011 (.H(net1011));
 TIEHIx1_ASAP7_75t_R _35061__1012 (.H(net1012));
 TIEHIx1_ASAP7_75t_R _35062__1013 (.H(net1013));
 TIEHIx1_ASAP7_75t_R _35063__1014 (.H(net1014));
 TIEHIx1_ASAP7_75t_R _35064__1015 (.H(net1015));
 TIEHIx1_ASAP7_75t_R _35065__1016 (.H(net1016));
 TIEHIx1_ASAP7_75t_R _35066__1017 (.H(net1017));
 TIEHIx1_ASAP7_75t_R _35067__1018 (.H(net1018));
 TIEHIx1_ASAP7_75t_R _35068__1019 (.H(net1019));
 TIEHIx1_ASAP7_75t_R _35069__1020 (.H(net1020));
 TIEHIx1_ASAP7_75t_R _35070__1021 (.H(net1021));
 TIEHIx1_ASAP7_75t_R _35071__1022 (.H(net1022));
 TIEHIx1_ASAP7_75t_R _35072__1023 (.H(net1023));
 TIEHIx1_ASAP7_75t_R _35073__1024 (.H(net1024));
 TIEHIx1_ASAP7_75t_R _35074__1025 (.H(net1025));
 TIEHIx1_ASAP7_75t_R _35075__1026 (.H(net1026));
 TIEHIx1_ASAP7_75t_R _35076__1027 (.H(net1027));
 TIEHIx1_ASAP7_75t_R _35077__1028 (.H(net1028));
 TIEHIx1_ASAP7_75t_R _35078__1029 (.H(net1029));
 TIEHIx1_ASAP7_75t_R _35079__1030 (.H(net1030));
 TIEHIx1_ASAP7_75t_R _35080__1031 (.H(net1031));
 TIEHIx1_ASAP7_75t_R _35081__1032 (.H(net1032));
 TIEHIx1_ASAP7_75t_R _35082__1033 (.H(net1033));
 TIEHIx1_ASAP7_75t_R _35083__1034 (.H(net1034));
 TIEHIx1_ASAP7_75t_R _35084__1035 (.H(net1035));
 TIEHIx1_ASAP7_75t_R _35085__1036 (.H(net1036));
 TIEHIx1_ASAP7_75t_R _35086__1037 (.H(net1037));
 TIEHIx1_ASAP7_75t_R _35087__1038 (.H(net1038));
 TIEHIx1_ASAP7_75t_R _35088__1039 (.H(net1039));
 TIEHIx1_ASAP7_75t_R _35089__1040 (.H(net1040));
 TIEHIx1_ASAP7_75t_R _35090__1041 (.H(net1041));
 TIEHIx1_ASAP7_75t_R _35091__1042 (.H(net1042));
 TIEHIx1_ASAP7_75t_R _35092__1043 (.H(net1043));
 TIEHIx1_ASAP7_75t_R _35093__1044 (.H(net1044));
 TIEHIx1_ASAP7_75t_R _35094__1045 (.H(net1045));
 TIEHIx1_ASAP7_75t_R _35095__1046 (.H(net1046));
 TIEHIx1_ASAP7_75t_R _35096__1047 (.H(net1047));
 TIEHIx1_ASAP7_75t_R _35097__1048 (.H(net1048));
 TIEHIx1_ASAP7_75t_R _35098__1049 (.H(net1049));
 TIEHIx1_ASAP7_75t_R _35099__1050 (.H(net1050));
 TIEHIx1_ASAP7_75t_R _35100__1051 (.H(net1051));
 TIEHIx1_ASAP7_75t_R _35101__1052 (.H(net1052));
 TIEHIx1_ASAP7_75t_R _35102__1053 (.H(net1053));
 TIEHIx1_ASAP7_75t_R _35103__1054 (.H(net1054));
 TIEHIx1_ASAP7_75t_R _35104__1055 (.H(net1055));
 TIEHIx1_ASAP7_75t_R _35105__1056 (.H(net1056));
 TIEHIx1_ASAP7_75t_R _35106__1057 (.H(net1057));
 TIEHIx1_ASAP7_75t_R _35107__1058 (.H(net1058));
 TIEHIx1_ASAP7_75t_R _35108__1059 (.H(net1059));
 TIEHIx1_ASAP7_75t_R _35109__1060 (.H(net1060));
 TIEHIx1_ASAP7_75t_R _35110__1061 (.H(net1061));
 TIEHIx1_ASAP7_75t_R _35111__1062 (.H(net1062));
 TIEHIx1_ASAP7_75t_R _35112__1063 (.H(net1063));
 TIEHIx1_ASAP7_75t_R _35113__1064 (.H(net1064));
 TIEHIx1_ASAP7_75t_R _35114__1065 (.H(net1065));
 TIEHIx1_ASAP7_75t_R _35115__1066 (.H(net1066));
 TIEHIx1_ASAP7_75t_R _35116__1067 (.H(net1067));
 TIEHIx1_ASAP7_75t_R _35117__1068 (.H(net1068));
 TIEHIx1_ASAP7_75t_R _35118__1069 (.H(net1069));
 TIEHIx1_ASAP7_75t_R _35119__1070 (.H(net1070));
 TIEHIx1_ASAP7_75t_R _35120__1071 (.H(net1071));
 TIEHIx1_ASAP7_75t_R _35121__1072 (.H(net1072));
 TIEHIx1_ASAP7_75t_R _35122__1073 (.H(net1073));
 TIEHIx1_ASAP7_75t_R _35123__1074 (.H(net1074));
 TIEHIx1_ASAP7_75t_R _35124__1075 (.H(net1075));
 TIEHIx1_ASAP7_75t_R _35125__1076 (.H(net1076));
 TIEHIx1_ASAP7_75t_R _35126__1077 (.H(net1077));
 TIEHIx1_ASAP7_75t_R _35127__1078 (.H(net1078));
 TIEHIx1_ASAP7_75t_R _35128__1079 (.H(net1079));
 TIEHIx1_ASAP7_75t_R _35129__1080 (.H(net1080));
 TIEHIx1_ASAP7_75t_R _35130__1081 (.H(net1081));
 TIEHIx1_ASAP7_75t_R _35131__1082 (.H(net1082));
 TIEHIx1_ASAP7_75t_R _35132__1083 (.H(net1083));
 TIEHIx1_ASAP7_75t_R _35133__1084 (.H(net1084));
 TIEHIx1_ASAP7_75t_R _35134__1085 (.H(net1085));
 TIEHIx1_ASAP7_75t_R _35135__1086 (.H(net1086));
 TIEHIx1_ASAP7_75t_R _35136__1087 (.H(net1087));
 TIEHIx1_ASAP7_75t_R _35137__1088 (.H(net1088));
 TIEHIx1_ASAP7_75t_R _35138__1089 (.H(net1089));
 TIEHIx1_ASAP7_75t_R _35139__1090 (.H(net1090));
 TIEHIx1_ASAP7_75t_R _35140__1091 (.H(net1091));
 TIEHIx1_ASAP7_75t_R _35141__1092 (.H(net1092));
 TIEHIx1_ASAP7_75t_R _35142__1093 (.H(net1093));
 TIEHIx1_ASAP7_75t_R _35143__1094 (.H(net1094));
 TIEHIx1_ASAP7_75t_R _35144__1095 (.H(net1095));
 TIEHIx1_ASAP7_75t_R _35145__1096 (.H(net1096));
 TIEHIx1_ASAP7_75t_R _35146__1097 (.H(net1097));
 TIEHIx1_ASAP7_75t_R _35147__1098 (.H(net1098));
 TIEHIx1_ASAP7_75t_R _35148__1099 (.H(net1099));
 TIEHIx1_ASAP7_75t_R _35149__1100 (.H(net1100));
 TIEHIx1_ASAP7_75t_R _35150__1101 (.H(net1101));
 TIEHIx1_ASAP7_75t_R _35151__1102 (.H(net1102));
 TIEHIx1_ASAP7_75t_R _35152__1103 (.H(net1103));
 TIEHIx1_ASAP7_75t_R _35153__1104 (.H(net1104));
 TIEHIx1_ASAP7_75t_R _35154__1105 (.H(net1105));
 TIEHIx1_ASAP7_75t_R _35155__1106 (.H(net1106));
 TIEHIx1_ASAP7_75t_R _35156__1107 (.H(net1107));
 TIEHIx1_ASAP7_75t_R _35157__1108 (.H(net1108));
 TIEHIx1_ASAP7_75t_R _35158__1109 (.H(net1109));
 TIEHIx1_ASAP7_75t_R _35159__1110 (.H(net1110));
 TIEHIx1_ASAP7_75t_R _35160__1111 (.H(net1111));
 TIEHIx1_ASAP7_75t_R _35161__1112 (.H(net1112));
 TIEHIx1_ASAP7_75t_R _35162__1113 (.H(net1113));
 TIEHIx1_ASAP7_75t_R _35163__1114 (.H(net1114));
 TIEHIx1_ASAP7_75t_R _35164__1115 (.H(net1115));
 TIEHIx1_ASAP7_75t_R _35165__1116 (.H(net1116));
 TIEHIx1_ASAP7_75t_R _35166__1117 (.H(net1117));
 TIEHIx1_ASAP7_75t_R _35167__1118 (.H(net1118));
 TIEHIx1_ASAP7_75t_R _35168__1119 (.H(net1119));
 TIEHIx1_ASAP7_75t_R _35169__1120 (.H(net1120));
 TIEHIx1_ASAP7_75t_R _35170__1121 (.H(net1121));
 TIEHIx1_ASAP7_75t_R _35171__1122 (.H(net1122));
 TIEHIx1_ASAP7_75t_R _35172__1123 (.H(net1123));
 TIEHIx1_ASAP7_75t_R _35173__1124 (.H(net1124));
 TIEHIx1_ASAP7_75t_R _35174__1125 (.H(net1125));
 TIEHIx1_ASAP7_75t_R _35175__1126 (.H(net1126));
 TIEHIx1_ASAP7_75t_R _35176__1127 (.H(net1127));
 TIEHIx1_ASAP7_75t_R _35177__1128 (.H(net1128));
 TIEHIx1_ASAP7_75t_R _35178__1129 (.H(net1129));
 TIEHIx1_ASAP7_75t_R _35179__1130 (.H(net1130));
 TIEHIx1_ASAP7_75t_R _35180__1131 (.H(net1131));
 TIEHIx1_ASAP7_75t_R _35181__1132 (.H(net1132));
 TIEHIx1_ASAP7_75t_R _35182__1133 (.H(net1133));
 TIEHIx1_ASAP7_75t_R _35183__1134 (.H(net1134));
 TIEHIx1_ASAP7_75t_R _35184__1135 (.H(net1135));
 TIEHIx1_ASAP7_75t_R _35185__1136 (.H(net1136));
 TIEHIx1_ASAP7_75t_R _35186__1137 (.H(net1137));
 TIEHIx1_ASAP7_75t_R _35187__1138 (.H(net1138));
 TIEHIx1_ASAP7_75t_R _35188__1139 (.H(net1139));
 TIEHIx1_ASAP7_75t_R _35189__1140 (.H(net1140));
 TIEHIx1_ASAP7_75t_R _35190__1141 (.H(net1141));
 TIEHIx1_ASAP7_75t_R _35191__1142 (.H(net1142));
 TIEHIx1_ASAP7_75t_R _35192__1143 (.H(net1143));
 TIEHIx1_ASAP7_75t_R _35193__1144 (.H(net1144));
 TIEHIx1_ASAP7_75t_R _35194__1145 (.H(net1145));
 TIEHIx1_ASAP7_75t_R _35195__1146 (.H(net1146));
 TIEHIx1_ASAP7_75t_R _35196__1147 (.H(net1147));
 TIEHIx1_ASAP7_75t_R _35197__1148 (.H(net1148));
 TIEHIx1_ASAP7_75t_R _35198__1149 (.H(net1149));
 TIEHIx1_ASAP7_75t_R _35199__1150 (.H(net1150));
 TIEHIx1_ASAP7_75t_R _35200__1151 (.H(net1151));
 TIEHIx1_ASAP7_75t_R _35201__1152 (.H(net1152));
 TIEHIx1_ASAP7_75t_R _35202__1153 (.H(net1153));
 TIEHIx1_ASAP7_75t_R _35203__1154 (.H(net1154));
 TIEHIx1_ASAP7_75t_R _35204__1155 (.H(net1155));
 TIEHIx1_ASAP7_75t_R _35205__1156 (.H(net1156));
 TIEHIx1_ASAP7_75t_R _35206__1157 (.H(net1157));
 TIEHIx1_ASAP7_75t_R _35207__1158 (.H(net1158));
 TIEHIx1_ASAP7_75t_R _35208__1159 (.H(net1159));
 TIEHIx1_ASAP7_75t_R _35209__1160 (.H(net1160));
 TIEHIx1_ASAP7_75t_R _35210__1161 (.H(net1161));
 TIEHIx1_ASAP7_75t_R _35211__1162 (.H(net1162));
 TIEHIx1_ASAP7_75t_R _35212__1163 (.H(net1163));
 TIEHIx1_ASAP7_75t_R _35213__1164 (.H(net1164));
 TIEHIx1_ASAP7_75t_R _35214__1165 (.H(net1165));
 TIEHIx1_ASAP7_75t_R _35215__1166 (.H(net1166));
 TIEHIx1_ASAP7_75t_R _35216__1167 (.H(net1167));
 TIEHIx1_ASAP7_75t_R _35217__1168 (.H(net1168));
 TIEHIx1_ASAP7_75t_R _35218__1169 (.H(net1169));
 TIEHIx1_ASAP7_75t_R _35219__1170 (.H(net1170));
 TIEHIx1_ASAP7_75t_R _35220__1171 (.H(net1171));
 TIEHIx1_ASAP7_75t_R _35221__1172 (.H(net1172));
 TIEHIx1_ASAP7_75t_R _35222__1173 (.H(net1173));
 TIEHIx1_ASAP7_75t_R _35223__1174 (.H(net1174));
 TIEHIx1_ASAP7_75t_R _35224__1175 (.H(net1175));
 TIEHIx1_ASAP7_75t_R _35225__1176 (.H(net1176));
 TIEHIx1_ASAP7_75t_R _35226__1177 (.H(net1177));
 TIEHIx1_ASAP7_75t_R _35227__1178 (.H(net1178));
 TIEHIx1_ASAP7_75t_R _35228__1179 (.H(net1179));
 TIEHIx1_ASAP7_75t_R _35229__1180 (.H(net1180));
 TIEHIx1_ASAP7_75t_R _35230__1181 (.H(net1181));
 TIEHIx1_ASAP7_75t_R _35231__1182 (.H(net1182));
 TIEHIx1_ASAP7_75t_R _35232__1183 (.H(net1183));
 TIEHIx1_ASAP7_75t_R _35233__1184 (.H(net1184));
 TIEHIx1_ASAP7_75t_R _35234__1185 (.H(net1185));
 TIEHIx1_ASAP7_75t_R _35235__1186 (.H(net1186));
 TIEHIx1_ASAP7_75t_R _35236__1187 (.H(net1187));
 TIEHIx1_ASAP7_75t_R _35237__1188 (.H(net1188));
 TIEHIx1_ASAP7_75t_R _35238__1189 (.H(net1189));
 TIEHIx1_ASAP7_75t_R _35239__1190 (.H(net1190));
 TIEHIx1_ASAP7_75t_R _35240__1191 (.H(net1191));
 TIEHIx1_ASAP7_75t_R _35241__1192 (.H(net1192));
 TIEHIx1_ASAP7_75t_R _35242__1193 (.H(net1193));
 TIEHIx1_ASAP7_75t_R _35243__1194 (.H(net1194));
 TIEHIx1_ASAP7_75t_R _35244__1195 (.H(net1195));
 TIEHIx1_ASAP7_75t_R _35245__1196 (.H(net1196));
 TIEHIx1_ASAP7_75t_R _35246__1197 (.H(net1197));
 TIEHIx1_ASAP7_75t_R _35247__1198 (.H(net1198));
 TIEHIx1_ASAP7_75t_R _35248__1199 (.H(net1199));
 TIEHIx1_ASAP7_75t_R _35249__1200 (.H(net1200));
 TIEHIx1_ASAP7_75t_R _35250__1201 (.H(net1201));
 TIEHIx1_ASAP7_75t_R _35251__1202 (.H(net1202));
 TIEHIx1_ASAP7_75t_R _35252__1203 (.H(net1203));
 TIEHIx1_ASAP7_75t_R _35253__1204 (.H(net1204));
 TIEHIx1_ASAP7_75t_R _35254__1205 (.H(net1205));
 TIEHIx1_ASAP7_75t_R _35255__1206 (.H(net1206));
 TIEHIx1_ASAP7_75t_R _35256__1207 (.H(net1207));
 TIEHIx1_ASAP7_75t_R _35257__1208 (.H(net1208));
 TIEHIx1_ASAP7_75t_R _35258__1209 (.H(net1209));
 TIEHIx1_ASAP7_75t_R _35259__1210 (.H(net1210));
 TIEHIx1_ASAP7_75t_R _35260__1211 (.H(net1211));
 TIEHIx1_ASAP7_75t_R _35261__1212 (.H(net1212));
 TIEHIx1_ASAP7_75t_R _35262__1213 (.H(net1213));
 TIEHIx1_ASAP7_75t_R _35263__1214 (.H(net1214));
 TIEHIx1_ASAP7_75t_R _35264__1215 (.H(net1215));
 TIEHIx1_ASAP7_75t_R _35265__1216 (.H(net1216));
 TIEHIx1_ASAP7_75t_R _35266__1217 (.H(net1217));
 TIEHIx1_ASAP7_75t_R _35267__1218 (.H(net1218));
 TIEHIx1_ASAP7_75t_R _35268__1219 (.H(net1219));
 TIEHIx1_ASAP7_75t_R _35269__1220 (.H(net1220));
 TIEHIx1_ASAP7_75t_R _35270__1221 (.H(net1221));
 TIEHIx1_ASAP7_75t_R _35271__1222 (.H(net1222));
 TIEHIx1_ASAP7_75t_R _35272__1223 (.H(net1223));
 TIEHIx1_ASAP7_75t_R _35273__1224 (.H(net1224));
 TIEHIx1_ASAP7_75t_R _35274__1225 (.H(net1225));
 TIEHIx1_ASAP7_75t_R _35275__1226 (.H(net1226));
 TIEHIx1_ASAP7_75t_R _35276__1227 (.H(net1227));
 TIEHIx1_ASAP7_75t_R _35277__1228 (.H(net1228));
 TIEHIx1_ASAP7_75t_R _35278__1229 (.H(net1229));
 TIEHIx1_ASAP7_75t_R _35279__1230 (.H(net1230));
 TIEHIx1_ASAP7_75t_R _35280__1231 (.H(net1231));
 TIEHIx1_ASAP7_75t_R _35281__1232 (.H(net1232));
 TIEHIx1_ASAP7_75t_R _35282__1233 (.H(net1233));
 TIEHIx1_ASAP7_75t_R _35283__1234 (.H(net1234));
 TIEHIx1_ASAP7_75t_R _35284__1235 (.H(net1235));
 TIEHIx1_ASAP7_75t_R _35285__1236 (.H(net1236));
 TIEHIx1_ASAP7_75t_R _35286__1237 (.H(net1237));
 TIEHIx1_ASAP7_75t_R _35287__1238 (.H(net1238));
 TIEHIx1_ASAP7_75t_R _35288__1239 (.H(net1239));
 TIEHIx1_ASAP7_75t_R _35289__1240 (.H(net1240));
 TIEHIx1_ASAP7_75t_R _35290__1241 (.H(net1241));
 TIEHIx1_ASAP7_75t_R _35291__1242 (.H(net1242));
 TIEHIx1_ASAP7_75t_R _35292__1243 (.H(net1243));
 TIEHIx1_ASAP7_75t_R _35293__1244 (.H(net1244));
 TIEHIx1_ASAP7_75t_R _35294__1245 (.H(net1245));
 TIEHIx1_ASAP7_75t_R _35295__1246 (.H(net1246));
 TIEHIx1_ASAP7_75t_R _35296__1247 (.H(net1247));
 TIEHIx1_ASAP7_75t_R _35297__1248 (.H(net1248));
 TIEHIx1_ASAP7_75t_R _35298__1249 (.H(net1249));
 TIEHIx1_ASAP7_75t_R _35299__1250 (.H(net1250));
 TIEHIx1_ASAP7_75t_R _35300__1251 (.H(net1251));
 TIEHIx1_ASAP7_75t_R _35301__1252 (.H(net1252));
 TIEHIx1_ASAP7_75t_R _35302__1253 (.H(net1253));
 TIEHIx1_ASAP7_75t_R _35303__1254 (.H(net1254));
 TIEHIx1_ASAP7_75t_R _35304__1255 (.H(net1255));
 TIEHIx1_ASAP7_75t_R _35305__1256 (.H(net1256));
 TIEHIx1_ASAP7_75t_R _35306__1257 (.H(net1257));
 TIEHIx1_ASAP7_75t_R _35307__1258 (.H(net1258));
 TIEHIx1_ASAP7_75t_R _35308__1259 (.H(net1259));
 TIEHIx1_ASAP7_75t_R _35309__1260 (.H(net1260));
 TIEHIx1_ASAP7_75t_R _35310__1261 (.H(net1261));
 TIEHIx1_ASAP7_75t_R _35311__1262 (.H(net1262));
 TIEHIx1_ASAP7_75t_R _35312__1263 (.H(net1263));
 TIEHIx1_ASAP7_75t_R _35313__1264 (.H(net1264));
 TIEHIx1_ASAP7_75t_R _35314__1265 (.H(net1265));
 TIEHIx1_ASAP7_75t_R _35315__1266 (.H(net1266));
 TIEHIx1_ASAP7_75t_R _35316__1267 (.H(net1267));
 TIEHIx1_ASAP7_75t_R _35317__1268 (.H(net1268));
 TIEHIx1_ASAP7_75t_R _35318__1269 (.H(net1269));
 TIEHIx1_ASAP7_75t_R _35319__1270 (.H(net1270));
 TIEHIx1_ASAP7_75t_R _35320__1271 (.H(net1271));
 TIEHIx1_ASAP7_75t_R _35321__1272 (.H(net1272));
 TIEHIx1_ASAP7_75t_R _35322__1273 (.H(net1273));
 TIEHIx1_ASAP7_75t_R _35323__1274 (.H(net1274));
 TIEHIx1_ASAP7_75t_R _35324__1275 (.H(net1275));
 TIEHIx1_ASAP7_75t_R _35325__1276 (.H(net1276));
 TIEHIx1_ASAP7_75t_R _35326__1277 (.H(net1277));
 TIEHIx1_ASAP7_75t_R _35327__1278 (.H(net1278));
 TIEHIx1_ASAP7_75t_R _35328__1279 (.H(net1279));
 TIEHIx1_ASAP7_75t_R _35329__1280 (.H(net1280));
 TIEHIx1_ASAP7_75t_R _35330__1281 (.H(net1281));
 TIEHIx1_ASAP7_75t_R _35331__1282 (.H(net1282));
 TIEHIx1_ASAP7_75t_R _35332__1283 (.H(net1283));
 TIEHIx1_ASAP7_75t_R _35333__1284 (.H(net1284));
 TIEHIx1_ASAP7_75t_R _35334__1285 (.H(net1285));
 TIEHIx1_ASAP7_75t_R _35335__1286 (.H(net1286));
 TIEHIx1_ASAP7_75t_R _35336__1287 (.H(net1287));
 TIEHIx1_ASAP7_75t_R _35337__1288 (.H(net1288));
 TIEHIx1_ASAP7_75t_R _35338__1289 (.H(net1289));
 TIEHIx1_ASAP7_75t_R _35339__1290 (.H(net1290));
 TIEHIx1_ASAP7_75t_R _35340__1291 (.H(net1291));
 TIEHIx1_ASAP7_75t_R _35341__1292 (.H(net1292));
 TIEHIx1_ASAP7_75t_R _35342__1293 (.H(net1293));
 TIEHIx1_ASAP7_75t_R _35343__1294 (.H(net1294));
 TIEHIx1_ASAP7_75t_R _35344__1295 (.H(net1295));
 TIEHIx1_ASAP7_75t_R _35345__1296 (.H(net1296));
 TIEHIx1_ASAP7_75t_R _35346__1297 (.H(net1297));
 TIEHIx1_ASAP7_75t_R _35347__1298 (.H(net1298));
 TIEHIx1_ASAP7_75t_R _35348__1299 (.H(net1299));
 TIEHIx1_ASAP7_75t_R _35349__1300 (.H(net1300));
 TIEHIx1_ASAP7_75t_R _35350__1301 (.H(net1301));
 TIEHIx1_ASAP7_75t_R _35351__1302 (.H(net1302));
 TIEHIx1_ASAP7_75t_R _35352__1303 (.H(net1303));
 TIEHIx1_ASAP7_75t_R _35353__1304 (.H(net1304));
 TIEHIx1_ASAP7_75t_R _35354__1305 (.H(net1305));
 TIEHIx1_ASAP7_75t_R _35355__1306 (.H(net1306));
 TIEHIx1_ASAP7_75t_R _35356__1307 (.H(net1307));
 TIEHIx1_ASAP7_75t_R _35357__1308 (.H(net1308));
 TIEHIx1_ASAP7_75t_R _35358__1309 (.H(net1309));
 TIEHIx1_ASAP7_75t_R _35359__1310 (.H(net1310));
 TIEHIx1_ASAP7_75t_R _35360__1311 (.H(net1311));
 TIEHIx1_ASAP7_75t_R _35361__1312 (.H(net1312));
 TIEHIx1_ASAP7_75t_R _35362__1313 (.H(net1313));
 TIEHIx1_ASAP7_75t_R _35363__1314 (.H(net1314));
 TIEHIx1_ASAP7_75t_R _35364__1315 (.H(net1315));
 TIEHIx1_ASAP7_75t_R _35365__1316 (.H(net1316));
 TIEHIx1_ASAP7_75t_R _35366__1317 (.H(net1317));
 TIEHIx1_ASAP7_75t_R _35367__1318 (.H(net1318));
 TIEHIx1_ASAP7_75t_R _35368__1319 (.H(net1319));
 TIEHIx1_ASAP7_75t_R _35369__1320 (.H(net1320));
 TIEHIx1_ASAP7_75t_R _35370__1321 (.H(net1321));
 TIEHIx1_ASAP7_75t_R _35371__1322 (.H(net1322));
 TIEHIx1_ASAP7_75t_R _35372__1323 (.H(net1323));
 TIEHIx1_ASAP7_75t_R _35373__1324 (.H(net1324));
 TIEHIx1_ASAP7_75t_R _35374__1325 (.H(net1325));
 TIEHIx1_ASAP7_75t_R _35375__1326 (.H(net1326));
 TIEHIx1_ASAP7_75t_R _35376__1327 (.H(net1327));
 TIEHIx1_ASAP7_75t_R _35377__1328 (.H(net1328));
 TIEHIx1_ASAP7_75t_R _35378__1329 (.H(net1329));
 TIEHIx1_ASAP7_75t_R _35379__1330 (.H(net1330));
 TIEHIx1_ASAP7_75t_R _35380__1331 (.H(net1331));
 TIEHIx1_ASAP7_75t_R _35381__1332 (.H(net1332));
 TIEHIx1_ASAP7_75t_R _35382__1333 (.H(net1333));
 TIEHIx1_ASAP7_75t_R _35383__1334 (.H(net1334));
 TIEHIx1_ASAP7_75t_R _35384__1335 (.H(net1335));
 TIEHIx1_ASAP7_75t_R _35385__1336 (.H(net1336));
 TIEHIx1_ASAP7_75t_R _35386__1337 (.H(net1337));
 TIEHIx1_ASAP7_75t_R _35387__1338 (.H(net1338));
 TIEHIx1_ASAP7_75t_R _35388__1339 (.H(net1339));
 TIEHIx1_ASAP7_75t_R _35389__1340 (.H(net1340));
 TIEHIx1_ASAP7_75t_R _35390__1341 (.H(net1341));
 TIEHIx1_ASAP7_75t_R _35391__1342 (.H(net1342));
 TIEHIx1_ASAP7_75t_R _35392__1343 (.H(net1343));
 TIEHIx1_ASAP7_75t_R _35393__1344 (.H(net1344));
 TIEHIx1_ASAP7_75t_R _35394__1345 (.H(net1345));
 TIEHIx1_ASAP7_75t_R _35395__1346 (.H(net1346));
 TIEHIx1_ASAP7_75t_R _35396__1347 (.H(net1347));
 TIEHIx1_ASAP7_75t_R _35397__1348 (.H(net1348));
 TIEHIx1_ASAP7_75t_R _35398__1349 (.H(net1349));
 TIEHIx1_ASAP7_75t_R _35399__1350 (.H(net1350));
 TIEHIx1_ASAP7_75t_R _35400__1351 (.H(net1351));
 TIEHIx1_ASAP7_75t_R _35401__1352 (.H(net1352));
 TIEHIx1_ASAP7_75t_R _35402__1353 (.H(net1353));
 TIEHIx1_ASAP7_75t_R _35403__1354 (.H(net1354));
 TIEHIx1_ASAP7_75t_R _35404__1355 (.H(net1355));
 TIEHIx1_ASAP7_75t_R _35405__1356 (.H(net1356));
 TIEHIx1_ASAP7_75t_R _35406__1357 (.H(net1357));
 TIEHIx1_ASAP7_75t_R _35407__1358 (.H(net1358));
 TIEHIx1_ASAP7_75t_R _35408__1359 (.H(net1359));
 TIEHIx1_ASAP7_75t_R _35409__1360 (.H(net1360));
 TIEHIx1_ASAP7_75t_R _35410__1361 (.H(net1361));
 TIEHIx1_ASAP7_75t_R _35411__1362 (.H(net1362));
 TIEHIx1_ASAP7_75t_R _35412__1363 (.H(net1363));
 TIEHIx1_ASAP7_75t_R _35413__1364 (.H(net1364));
 TIEHIx1_ASAP7_75t_R _35414__1365 (.H(net1365));
 TIEHIx1_ASAP7_75t_R _35415__1366 (.H(net1366));
 TIEHIx1_ASAP7_75t_R _35416__1367 (.H(net1367));
 TIEHIx1_ASAP7_75t_R _35417__1368 (.H(net1368));
 TIEHIx1_ASAP7_75t_R _35418__1369 (.H(net1369));
 TIEHIx1_ASAP7_75t_R _35419__1370 (.H(net1370));
 TIEHIx1_ASAP7_75t_R _35420__1371 (.H(net1371));
 TIEHIx1_ASAP7_75t_R _35421__1372 (.H(net1372));
 TIEHIx1_ASAP7_75t_R _35422__1373 (.H(net1373));
 TIEHIx1_ASAP7_75t_R _35423__1374 (.H(net1374));
 TIEHIx1_ASAP7_75t_R _35424__1375 (.H(net1375));
 TIEHIx1_ASAP7_75t_R _35425__1376 (.H(net1376));
 TIEHIx1_ASAP7_75t_R _35426__1377 (.H(net1377));
 TIEHIx1_ASAP7_75t_R _35427__1378 (.H(net1378));
 TIEHIx1_ASAP7_75t_R _35428__1379 (.H(net1379));
 TIEHIx1_ASAP7_75t_R _35429__1380 (.H(net1380));
 TIEHIx1_ASAP7_75t_R _35430__1381 (.H(net1381));
 TIEHIx1_ASAP7_75t_R _35431__1382 (.H(net1382));
 TIEHIx1_ASAP7_75t_R _35432__1383 (.H(net1383));
 TIEHIx1_ASAP7_75t_R _35433__1384 (.H(net1384));
 TIEHIx1_ASAP7_75t_R _35434__1385 (.H(net1385));
 TIEHIx1_ASAP7_75t_R _35435__1386 (.H(net1386));
 TIEHIx1_ASAP7_75t_R _35436__1387 (.H(net1387));
 TIEHIx1_ASAP7_75t_R _35437__1388 (.H(net1388));
 TIEHIx1_ASAP7_75t_R _35438__1389 (.H(net1389));
 TIEHIx1_ASAP7_75t_R _35439__1390 (.H(net1390));
 TIEHIx1_ASAP7_75t_R _35440__1391 (.H(net1391));
 TIEHIx1_ASAP7_75t_R _35441__1392 (.H(net1392));
 TIEHIx1_ASAP7_75t_R _35442__1393 (.H(net1393));
 TIEHIx1_ASAP7_75t_R _35443__1394 (.H(net1394));
 TIEHIx1_ASAP7_75t_R _35444__1395 (.H(net1395));
 TIEHIx1_ASAP7_75t_R _35445__1396 (.H(net1396));
 TIEHIx1_ASAP7_75t_R _35446__1397 (.H(net1397));
 TIEHIx1_ASAP7_75t_R _35447__1398 (.H(net1398));
 TIEHIx1_ASAP7_75t_R _35448__1399 (.H(net1399));
 TIEHIx1_ASAP7_75t_R _35449__1400 (.H(net1400));
 TIEHIx1_ASAP7_75t_R _35450__1401 (.H(net1401));
 TIEHIx1_ASAP7_75t_R _35451__1402 (.H(net1402));
 TIEHIx1_ASAP7_75t_R _35452__1403 (.H(net1403));
 TIEHIx1_ASAP7_75t_R _35453__1404 (.H(net1404));
 TIEHIx1_ASAP7_75t_R _35454__1405 (.H(net1405));
 TIEHIx1_ASAP7_75t_R _35455__1406 (.H(net1406));
 TIEHIx1_ASAP7_75t_R _35456__1407 (.H(net1407));
 TIEHIx1_ASAP7_75t_R _35457__1408 (.H(net1408));
 TIEHIx1_ASAP7_75t_R _35458__1409 (.H(net1409));
 TIEHIx1_ASAP7_75t_R _35459__1410 (.H(net1410));
 TIEHIx1_ASAP7_75t_R _35460__1411 (.H(net1411));
 TIEHIx1_ASAP7_75t_R _35461__1412 (.H(net1412));
 TIEHIx1_ASAP7_75t_R _35462__1413 (.H(net1413));
 TIEHIx1_ASAP7_75t_R _35463__1414 (.H(net1414));
 TIEHIx1_ASAP7_75t_R _35464__1415 (.H(net1415));
 TIEHIx1_ASAP7_75t_R _35465__1416 (.H(net1416));
 TIEHIx1_ASAP7_75t_R _35466__1417 (.H(net1417));
 TIEHIx1_ASAP7_75t_R _35467__1418 (.H(net1418));
 TIEHIx1_ASAP7_75t_R _35468__1419 (.H(net1419));
 TIEHIx1_ASAP7_75t_R _35469__1420 (.H(net1420));
 TIEHIx1_ASAP7_75t_R _35470__1421 (.H(net1421));
 TIEHIx1_ASAP7_75t_R _35471__1422 (.H(net1422));
 TIEHIx1_ASAP7_75t_R _35472__1423 (.H(net1423));
 TIEHIx1_ASAP7_75t_R _35473__1424 (.H(net1424));
 TIEHIx1_ASAP7_75t_R _35474__1425 (.H(net1425));
 TIEHIx1_ASAP7_75t_R _35475__1426 (.H(net1426));
 TIEHIx1_ASAP7_75t_R _35476__1427 (.H(net1427));
 TIEHIx1_ASAP7_75t_R _35477__1428 (.H(net1428));
 TIEHIx1_ASAP7_75t_R _35478__1429 (.H(net1429));
 TIEHIx1_ASAP7_75t_R _35479__1430 (.H(net1430));
 TIEHIx1_ASAP7_75t_R _35480__1431 (.H(net1431));
 TIEHIx1_ASAP7_75t_R _35481__1432 (.H(net1432));
 TIEHIx1_ASAP7_75t_R _35482__1433 (.H(net1433));
 TIEHIx1_ASAP7_75t_R _35483__1434 (.H(net1434));
 TIEHIx1_ASAP7_75t_R _35484__1435 (.H(net1435));
 TIEHIx1_ASAP7_75t_R _35485__1436 (.H(net1436));
 TIEHIx1_ASAP7_75t_R _35486__1437 (.H(net1437));
 TIEHIx1_ASAP7_75t_R _35487__1438 (.H(net1438));
 TIEHIx1_ASAP7_75t_R _35488__1439 (.H(net1439));
 TIEHIx1_ASAP7_75t_R _35489__1440 (.H(net1440));
 TIEHIx1_ASAP7_75t_R _35490__1441 (.H(net1441));
 TIEHIx1_ASAP7_75t_R _35491__1442 (.H(net1442));
 TIEHIx1_ASAP7_75t_R _35492__1443 (.H(net1443));
 TIEHIx1_ASAP7_75t_R _35493__1444 (.H(net1444));
 TIEHIx1_ASAP7_75t_R _35494__1445 (.H(net1445));
 TIEHIx1_ASAP7_75t_R _35495__1446 (.H(net1446));
 TIEHIx1_ASAP7_75t_R _35496__1447 (.H(net1447));
 TIEHIx1_ASAP7_75t_R _35497__1448 (.H(net1448));
 TIEHIx1_ASAP7_75t_R _35498__1449 (.H(net1449));
 TIEHIx1_ASAP7_75t_R _35499__1450 (.H(net1450));
 TIEHIx1_ASAP7_75t_R _35500__1451 (.H(net1451));
 TIEHIx1_ASAP7_75t_R _35501__1452 (.H(net1452));
 TIEHIx1_ASAP7_75t_R _35502__1453 (.H(net1453));
 TIEHIx1_ASAP7_75t_R _35503__1454 (.H(net1454));
 TIEHIx1_ASAP7_75t_R _35504__1455 (.H(net1455));
 TIEHIx1_ASAP7_75t_R _35505__1456 (.H(net1456));
 TIEHIx1_ASAP7_75t_R _35506__1457 (.H(net1457));
 TIEHIx1_ASAP7_75t_R _35507__1458 (.H(net1458));
 TIEHIx1_ASAP7_75t_R _35508__1459 (.H(net1459));
 TIEHIx1_ASAP7_75t_R _35509__1460 (.H(net1460));
 TIEHIx1_ASAP7_75t_R _35510__1461 (.H(net1461));
 TIEHIx1_ASAP7_75t_R _35511__1462 (.H(net1462));
 TIEHIx1_ASAP7_75t_R _35512__1463 (.H(net1463));
 TIEHIx1_ASAP7_75t_R _35513__1464 (.H(net1464));
 TIEHIx1_ASAP7_75t_R _35514__1465 (.H(net1465));
 TIEHIx1_ASAP7_75t_R _35515__1466 (.H(net1466));
 TIEHIx1_ASAP7_75t_R _35516__1467 (.H(net1467));
 TIEHIx1_ASAP7_75t_R _35517__1468 (.H(net1468));
 TIEHIx1_ASAP7_75t_R _35518__1469 (.H(net1469));
 TIEHIx1_ASAP7_75t_R _35519__1470 (.H(net1470));
 TIEHIx1_ASAP7_75t_R _35520__1471 (.H(net1471));
 TIEHIx1_ASAP7_75t_R _35521__1472 (.H(net1472));
 TIEHIx1_ASAP7_75t_R _35522__1473 (.H(net1473));
 TIEHIx1_ASAP7_75t_R _35523__1474 (.H(net1474));
 TIEHIx1_ASAP7_75t_R _35524__1475 (.H(net1475));
 TIEHIx1_ASAP7_75t_R _35525__1476 (.H(net1476));
 TIEHIx1_ASAP7_75t_R _35526__1477 (.H(net1477));
 TIEHIx1_ASAP7_75t_R _35527__1478 (.H(net1478));
 TIEHIx1_ASAP7_75t_R _35528__1479 (.H(net1479));
 TIEHIx1_ASAP7_75t_R _35529__1480 (.H(net1480));
 TIEHIx1_ASAP7_75t_R _35530__1481 (.H(net1481));
 TIEHIx1_ASAP7_75t_R _35531__1482 (.H(net1482));
 TIEHIx1_ASAP7_75t_R _35532__1483 (.H(net1483));
 TIEHIx1_ASAP7_75t_R _35533__1484 (.H(net1484));
 TIEHIx1_ASAP7_75t_R _35534__1485 (.H(net1485));
 TIEHIx1_ASAP7_75t_R _35535__1486 (.H(net1486));
 TIEHIx1_ASAP7_75t_R _35536__1487 (.H(net1487));
 TIEHIx1_ASAP7_75t_R _35537__1488 (.H(net1488));
 TIEHIx1_ASAP7_75t_R _35538__1489 (.H(net1489));
 TIEHIx1_ASAP7_75t_R _35539__1490 (.H(net1490));
 TIEHIx1_ASAP7_75t_R _35540__1491 (.H(net1491));
 TIEHIx1_ASAP7_75t_R _35541__1492 (.H(net1492));
 TIEHIx1_ASAP7_75t_R _35542__1493 (.H(net1493));
 TIEHIx1_ASAP7_75t_R _35543__1494 (.H(net1494));
 TIEHIx1_ASAP7_75t_R _35544__1495 (.H(net1495));
 TIEHIx1_ASAP7_75t_R _35545__1496 (.H(net1496));
 TIEHIx1_ASAP7_75t_R _35546__1497 (.H(net1497));
 TIEHIx1_ASAP7_75t_R _35547__1498 (.H(net1498));
 TIEHIx1_ASAP7_75t_R _35548__1499 (.H(net1499));
 TIEHIx1_ASAP7_75t_R _35549__1500 (.H(net1500));
 TIEHIx1_ASAP7_75t_R _35550__1501 (.H(net1501));
 TIEHIx1_ASAP7_75t_R _35551__1502 (.H(net1502));
 TIEHIx1_ASAP7_75t_R _35552__1503 (.H(net1503));
 TIEHIx1_ASAP7_75t_R _35553__1504 (.H(net1504));
 TIEHIx1_ASAP7_75t_R _35554__1505 (.H(net1505));
 TIEHIx1_ASAP7_75t_R _35555__1506 (.H(net1506));
 TIEHIx1_ASAP7_75t_R _35556__1507 (.H(net1507));
 TIEHIx1_ASAP7_75t_R _35557__1508 (.H(net1508));
 TIEHIx1_ASAP7_75t_R _35558__1509 (.H(net1509));
 TIEHIx1_ASAP7_75t_R _35559__1510 (.H(net1510));
 TIEHIx1_ASAP7_75t_R _35560__1511 (.H(net1511));
 TIEHIx1_ASAP7_75t_R _35561__1512 (.H(net1512));
 TIEHIx1_ASAP7_75t_R _35562__1513 (.H(net1513));
 TIEHIx1_ASAP7_75t_R _35563__1514 (.H(net1514));
 TIEHIx1_ASAP7_75t_R _35564__1515 (.H(net1515));
 TIEHIx1_ASAP7_75t_R _35565__1516 (.H(net1516));
 TIEHIx1_ASAP7_75t_R _35566__1517 (.H(net1517));
 TIEHIx1_ASAP7_75t_R _35567__1518 (.H(net1518));
 TIEHIx1_ASAP7_75t_R _35568__1519 (.H(net1519));
 TIEHIx1_ASAP7_75t_R _35569__1520 (.H(net1520));
 TIEHIx1_ASAP7_75t_R _35570__1521 (.H(net1521));
 TIEHIx1_ASAP7_75t_R _35571__1522 (.H(net1522));
 TIEHIx1_ASAP7_75t_R _35572__1523 (.H(net1523));
 TIEHIx1_ASAP7_75t_R _35573__1524 (.H(net1524));
 TIEHIx1_ASAP7_75t_R _35574__1525 (.H(net1525));
 TIEHIx1_ASAP7_75t_R _35575__1526 (.H(net1526));
 TIEHIx1_ASAP7_75t_R _35576__1527 (.H(net1527));
 TIEHIx1_ASAP7_75t_R _35577__1528 (.H(net1528));
 TIEHIx1_ASAP7_75t_R _35578__1529 (.H(net1529));
 TIEHIx1_ASAP7_75t_R _35579__1530 (.H(net1530));
 TIEHIx1_ASAP7_75t_R _35580__1531 (.H(net1531));
 TIEHIx1_ASAP7_75t_R _35581__1532 (.H(net1532));
 TIEHIx1_ASAP7_75t_R _35582__1533 (.H(net1533));
 TIEHIx1_ASAP7_75t_R _35583__1534 (.H(net1534));
 TIEHIx1_ASAP7_75t_R _35584__1535 (.H(net1535));
 TIEHIx1_ASAP7_75t_R _35585__1536 (.H(net1536));
 TIEHIx1_ASAP7_75t_R _35586__1537 (.H(net1537));
 TIEHIx1_ASAP7_75t_R _35587__1538 (.H(net1538));
 TIEHIx1_ASAP7_75t_R _35588__1539 (.H(net1539));
 TIEHIx1_ASAP7_75t_R _35589__1540 (.H(net1540));
 TIEHIx1_ASAP7_75t_R _35590__1541 (.H(net1541));
 TIEHIx1_ASAP7_75t_R _35591__1542 (.H(net1542));
 TIEHIx1_ASAP7_75t_R _35592__1543 (.H(net1543));
 TIEHIx1_ASAP7_75t_R _35593__1544 (.H(net1544));
 TIEHIx1_ASAP7_75t_R _35594__1545 (.H(net1545));
 TIEHIx1_ASAP7_75t_R _35595__1546 (.H(net1546));
 TIEHIx1_ASAP7_75t_R _35596__1547 (.H(net1547));
 TIEHIx1_ASAP7_75t_R _35597__1548 (.H(net1548));
 TIEHIx1_ASAP7_75t_R _35598__1549 (.H(net1549));
 TIEHIx1_ASAP7_75t_R _35599__1550 (.H(net1550));
 TIEHIx1_ASAP7_75t_R _35600__1551 (.H(net1551));
 TIEHIx1_ASAP7_75t_R _35601__1552 (.H(net1552));
 TIEHIx1_ASAP7_75t_R _35602__1553 (.H(net1553));
 TIEHIx1_ASAP7_75t_R _35603__1554 (.H(net1554));
 TIEHIx1_ASAP7_75t_R _35604__1555 (.H(net1555));
 TIEHIx1_ASAP7_75t_R _35605__1556 (.H(net1556));
 TIEHIx1_ASAP7_75t_R _35606__1557 (.H(net1557));
 TIEHIx1_ASAP7_75t_R _35607__1558 (.H(net1558));
 TIEHIx1_ASAP7_75t_R _35608__1559 (.H(net1559));
 TIEHIx1_ASAP7_75t_R _35609__1560 (.H(net1560));
 TIEHIx1_ASAP7_75t_R _35610__1561 (.H(net1561));
 TIEHIx1_ASAP7_75t_R _35611__1562 (.H(net1562));
 TIEHIx1_ASAP7_75t_R _35612__1563 (.H(net1563));
 TIEHIx1_ASAP7_75t_R _35613__1564 (.H(net1564));
 TIEHIx1_ASAP7_75t_R _35614__1565 (.H(net1565));
 TIEHIx1_ASAP7_75t_R _35615__1566 (.H(net1566));
 TIEHIx1_ASAP7_75t_R _35616__1567 (.H(net1567));
 TIEHIx1_ASAP7_75t_R _35617__1568 (.H(net1568));
 TIEHIx1_ASAP7_75t_R _35618__1569 (.H(net1569));
 TIEHIx1_ASAP7_75t_R _35619__1570 (.H(net1570));
 TIEHIx1_ASAP7_75t_R _35620__1571 (.H(net1571));
 TIEHIx1_ASAP7_75t_R _35621__1572 (.H(net1572));
 TIEHIx1_ASAP7_75t_R _35622__1573 (.H(net1573));
 TIEHIx1_ASAP7_75t_R _35623__1574 (.H(net1574));
 TIEHIx1_ASAP7_75t_R _35624__1575 (.H(net1575));
 TIEHIx1_ASAP7_75t_R _35625__1576 (.H(net1576));
 TIEHIx1_ASAP7_75t_R _35626__1577 (.H(net1577));
 TIEHIx1_ASAP7_75t_R _35627__1578 (.H(net1578));
 TIEHIx1_ASAP7_75t_R _35628__1579 (.H(net1579));
 TIEHIx1_ASAP7_75t_R _35629__1580 (.H(net1580));
 TIEHIx1_ASAP7_75t_R _35630__1581 (.H(net1581));
 TIEHIx1_ASAP7_75t_R _35631__1582 (.H(net1582));
 TIEHIx1_ASAP7_75t_R _35632__1583 (.H(net1583));
 TIEHIx1_ASAP7_75t_R _35633__1584 (.H(net1584));
 TIEHIx1_ASAP7_75t_R _35634__1585 (.H(net1585));
 TIEHIx1_ASAP7_75t_R _35635__1586 (.H(net1586));
 TIEHIx1_ASAP7_75t_R _35636__1587 (.H(net1587));
 TIEHIx1_ASAP7_75t_R _35637__1588 (.H(net1588));
 TIEHIx1_ASAP7_75t_R _35638__1589 (.H(net1589));
 TIEHIx1_ASAP7_75t_R _35639__1590 (.H(net1590));
 TIEHIx1_ASAP7_75t_R _35640__1591 (.H(net1591));
 TIEHIx1_ASAP7_75t_R _35641__1592 (.H(net1592));
 TIEHIx1_ASAP7_75t_R _35642__1593 (.H(net1593));
 TIEHIx1_ASAP7_75t_R _35643__1594 (.H(net1594));
 TIEHIx1_ASAP7_75t_R _35644__1595 (.H(net1595));
 TIEHIx1_ASAP7_75t_R _35645__1596 (.H(net1596));
 TIEHIx1_ASAP7_75t_R _35646__1597 (.H(net1597));
 TIEHIx1_ASAP7_75t_R _35647__1598 (.H(net1598));
 TIEHIx1_ASAP7_75t_R _35648__1599 (.H(net1599));
 TIEHIx1_ASAP7_75t_R _35649__1600 (.H(net1600));
 TIEHIx1_ASAP7_75t_R _35650__1601 (.H(net1601));
 TIEHIx1_ASAP7_75t_R _35651__1602 (.H(net1602));
 TIEHIx1_ASAP7_75t_R _35652__1603 (.H(net1603));
 TIEHIx1_ASAP7_75t_R _35653__1604 (.H(net1604));
 TIEHIx1_ASAP7_75t_R _35654__1605 (.H(net1605));
 TIEHIx1_ASAP7_75t_R _35655__1606 (.H(net1606));
 TIEHIx1_ASAP7_75t_R _35656__1607 (.H(net1607));
 TIEHIx1_ASAP7_75t_R _35657__1608 (.H(net1608));
 TIEHIx1_ASAP7_75t_R _35658__1609 (.H(net1609));
 TIEHIx1_ASAP7_75t_R _35659__1610 (.H(net1610));
 TIEHIx1_ASAP7_75t_R _35660__1611 (.H(net1611));
 TIEHIx1_ASAP7_75t_R _35661__1612 (.H(net1612));
 TIEHIx1_ASAP7_75t_R _35662__1613 (.H(net1613));
 TIEHIx1_ASAP7_75t_R _35663__1614 (.H(net1614));
 TIEHIx1_ASAP7_75t_R _35664__1615 (.H(net1615));
 TIEHIx1_ASAP7_75t_R _35665__1616 (.H(net1616));
 TIEHIx1_ASAP7_75t_R _35666__1617 (.H(net1617));
 TIEHIx1_ASAP7_75t_R _35667__1618 (.H(net1618));
 TIEHIx1_ASAP7_75t_R _35668__1619 (.H(net1619));
 TIEHIx1_ASAP7_75t_R _35669__1620 (.H(net1620));
 TIEHIx1_ASAP7_75t_R _35670__1621 (.H(net1621));
 TIEHIx1_ASAP7_75t_R _35671__1622 (.H(net1622));
 TIEHIx1_ASAP7_75t_R _35672__1623 (.H(net1623));
 TIEHIx1_ASAP7_75t_R _35673__1624 (.H(net1624));
 TIEHIx1_ASAP7_75t_R _35674__1625 (.H(net1625));
 TIEHIx1_ASAP7_75t_R _35675__1626 (.H(net1626));
 TIEHIx1_ASAP7_75t_R _35676__1627 (.H(net1627));
 TIEHIx1_ASAP7_75t_R _35677__1628 (.H(net1628));
 TIEHIx1_ASAP7_75t_R _35678__1629 (.H(net1629));
 TIEHIx1_ASAP7_75t_R _35679__1630 (.H(net1630));
 TIEHIx1_ASAP7_75t_R _35680__1631 (.H(net1631));
 TIEHIx1_ASAP7_75t_R _35681__1632 (.H(net1632));
 TIEHIx1_ASAP7_75t_R _35682__1633 (.H(net1633));
 TIEHIx1_ASAP7_75t_R _35683__1634 (.H(net1634));
 TIEHIx1_ASAP7_75t_R _35684__1635 (.H(net1635));
 TIEHIx1_ASAP7_75t_R _35685__1636 (.H(net1636));
 TIEHIx1_ASAP7_75t_R _35686__1637 (.H(net1637));
 TIEHIx1_ASAP7_75t_R _35687__1638 (.H(net1638));
 TIEHIx1_ASAP7_75t_R _35688__1639 (.H(net1639));
 TIEHIx1_ASAP7_75t_R _35689__1640 (.H(net1640));
 TIEHIx1_ASAP7_75t_R _35690__1641 (.H(net1641));
 TIEHIx1_ASAP7_75t_R _35691__1642 (.H(net1642));
 TIEHIx1_ASAP7_75t_R _35692__1643 (.H(net1643));
 TIEHIx1_ASAP7_75t_R _35693__1644 (.H(net1644));
 TIEHIx1_ASAP7_75t_R _35694__1645 (.H(net1645));
 TIEHIx1_ASAP7_75t_R _35695__1646 (.H(net1646));
 TIEHIx1_ASAP7_75t_R _35696__1647 (.H(net1647));
 TIEHIx1_ASAP7_75t_R _35697__1648 (.H(net1648));
 TIEHIx1_ASAP7_75t_R _35698__1649 (.H(net1649));
 TIEHIx1_ASAP7_75t_R _35699__1650 (.H(net1650));
 TIEHIx1_ASAP7_75t_R _35700__1651 (.H(net1651));
 TIEHIx1_ASAP7_75t_R _35701__1652 (.H(net1652));
 TIEHIx1_ASAP7_75t_R _35702__1653 (.H(net1653));
 TIEHIx1_ASAP7_75t_R _35703__1654 (.H(net1654));
 TIEHIx1_ASAP7_75t_R _35704__1655 (.H(net1655));
 TIEHIx1_ASAP7_75t_R _35705__1656 (.H(net1656));
 TIEHIx1_ASAP7_75t_R _35706__1657 (.H(net1657));
 TIEHIx1_ASAP7_75t_R _35707__1658 (.H(net1658));
 TIEHIx1_ASAP7_75t_R _35708__1659 (.H(net1659));
 TIEHIx1_ASAP7_75t_R _35709__1660 (.H(net1660));
 TIEHIx1_ASAP7_75t_R _35710__1661 (.H(net1661));
 TIEHIx1_ASAP7_75t_R _35711__1662 (.H(net1662));
 TIEHIx1_ASAP7_75t_R _35712__1663 (.H(net1663));
 TIEHIx1_ASAP7_75t_R _35713__1664 (.H(net1664));
 TIEHIx1_ASAP7_75t_R _35714__1665 (.H(net1665));
 TIEHIx1_ASAP7_75t_R _35715__1666 (.H(net1666));
 TIEHIx1_ASAP7_75t_R _35716__1667 (.H(net1667));
 TIEHIx1_ASAP7_75t_R _35717__1668 (.H(net1668));
 TIEHIx1_ASAP7_75t_R _35718__1669 (.H(net1669));
 TIEHIx1_ASAP7_75t_R _35719__1670 (.H(net1670));
 TIEHIx1_ASAP7_75t_R _35720__1671 (.H(net1671));
 TIEHIx1_ASAP7_75t_R _35721__1672 (.H(net1672));
 TIEHIx1_ASAP7_75t_R _35722__1673 (.H(net1673));
 TIEHIx1_ASAP7_75t_R _35723__1674 (.H(net1674));
 TIEHIx1_ASAP7_75t_R _35724__1675 (.H(net1675));
 TIEHIx1_ASAP7_75t_R _35725__1676 (.H(net1676));
 TIEHIx1_ASAP7_75t_R _35726__1677 (.H(net1677));
 TIEHIx1_ASAP7_75t_R _35727__1678 (.H(net1678));
 TIEHIx1_ASAP7_75t_R _35728__1679 (.H(net1679));
 TIEHIx1_ASAP7_75t_R _35729__1680 (.H(net1680));
 TIEHIx1_ASAP7_75t_R _35730__1681 (.H(net1681));
 TIEHIx1_ASAP7_75t_R _35731__1682 (.H(net1682));
 TIEHIx1_ASAP7_75t_R _35732__1683 (.H(net1683));
 TIEHIx1_ASAP7_75t_R _35733__1684 (.H(net1684));
 TIEHIx1_ASAP7_75t_R _35734__1685 (.H(net1685));
 TIEHIx1_ASAP7_75t_R _35735__1686 (.H(net1686));
 TIEHIx1_ASAP7_75t_R _35736__1687 (.H(net1687));
 TIEHIx1_ASAP7_75t_R _35737__1688 (.H(net1688));
 TIEHIx1_ASAP7_75t_R _35738__1689 (.H(net1689));
 TIEHIx1_ASAP7_75t_R _35739__1690 (.H(net1690));
 TIEHIx1_ASAP7_75t_R _35740__1691 (.H(net1691));
 TIEHIx1_ASAP7_75t_R _35741__1692 (.H(net1692));
 TIEHIx1_ASAP7_75t_R _35742__1693 (.H(net1693));
 TIEHIx1_ASAP7_75t_R _35743__1694 (.H(net1694));
 TIEHIx1_ASAP7_75t_R _35744__1695 (.H(net1695));
 TIEHIx1_ASAP7_75t_R _35745__1696 (.H(net1696));
 TIEHIx1_ASAP7_75t_R _35746__1697 (.H(net1697));
 TIEHIx1_ASAP7_75t_R _35747__1698 (.H(net1698));
 TIEHIx1_ASAP7_75t_R _35748__1699 (.H(net1699));
 TIEHIx1_ASAP7_75t_R _35749__1700 (.H(net1700));
 TIEHIx1_ASAP7_75t_R _35750__1701 (.H(net1701));
 TIEHIx1_ASAP7_75t_R _35751__1702 (.H(net1702));
 TIEHIx1_ASAP7_75t_R _35752__1703 (.H(net1703));
 TIEHIx1_ASAP7_75t_R _35753__1704 (.H(net1704));
 TIEHIx1_ASAP7_75t_R _35754__1705 (.H(net1705));
 TIEHIx1_ASAP7_75t_R _35755__1706 (.H(net1706));
 TIEHIx1_ASAP7_75t_R _35756__1707 (.H(net1707));
 TIEHIx1_ASAP7_75t_R _35757__1708 (.H(net1708));
 TIEHIx1_ASAP7_75t_R _35758__1709 (.H(net1709));
 TIEHIx1_ASAP7_75t_R _35759__1710 (.H(net1710));
 TIEHIx1_ASAP7_75t_R _35760__1711 (.H(net1711));
 TIEHIx1_ASAP7_75t_R _35761__1712 (.H(net1712));
 TIEHIx1_ASAP7_75t_R _35762__1713 (.H(net1713));
 TIEHIx1_ASAP7_75t_R _35763__1714 (.H(net1714));
 TIEHIx1_ASAP7_75t_R _35764__1715 (.H(net1715));
 TIEHIx1_ASAP7_75t_R _35765__1716 (.H(net1716));
 TIEHIx1_ASAP7_75t_R _35766__1717 (.H(net1717));
 TIEHIx1_ASAP7_75t_R _35767__1718 (.H(net1718));
 TIEHIx1_ASAP7_75t_R _35768__1719 (.H(net1719));
 TIEHIx1_ASAP7_75t_R _35769__1720 (.H(net1720));
 TIEHIx1_ASAP7_75t_R _35770__1721 (.H(net1721));
 TIEHIx1_ASAP7_75t_R _35771__1722 (.H(net1722));
 TIEHIx1_ASAP7_75t_R _35772__1723 (.H(net1723));
 TIEHIx1_ASAP7_75t_R _35773__1724 (.H(net1724));
 TIEHIx1_ASAP7_75t_R _35774__1725 (.H(net1725));
 TIEHIx1_ASAP7_75t_R _35775__1726 (.H(net1726));
 TIEHIx1_ASAP7_75t_R _35776__1727 (.H(net1727));
 TIEHIx1_ASAP7_75t_R _35777__1728 (.H(net1728));
 TIEHIx1_ASAP7_75t_R _35778__1729 (.H(net1729));
 TIEHIx1_ASAP7_75t_R _35779__1730 (.H(net1730));
 TIEHIx1_ASAP7_75t_R _35780__1731 (.H(net1731));
 TIEHIx1_ASAP7_75t_R _35781__1732 (.H(net1732));
 TIEHIx1_ASAP7_75t_R _35782__1733 (.H(net1733));
 TIEHIx1_ASAP7_75t_R _35783__1734 (.H(net1734));
 TIEHIx1_ASAP7_75t_R _35784__1735 (.H(net1735));
 TIEHIx1_ASAP7_75t_R _35785__1736 (.H(net1736));
 TIEHIx1_ASAP7_75t_R _35786__1737 (.H(net1737));
 TIEHIx1_ASAP7_75t_R _35787__1738 (.H(net1738));
 TIEHIx1_ASAP7_75t_R _35788__1739 (.H(net1739));
 TIEHIx1_ASAP7_75t_R _35789__1740 (.H(net1740));
 TIEHIx1_ASAP7_75t_R _35790__1741 (.H(net1741));
 TIEHIx1_ASAP7_75t_R _35791__1742 (.H(net1742));
 TIEHIx1_ASAP7_75t_R _35792__1743 (.H(net1743));
 TIEHIx1_ASAP7_75t_R _35793__1744 (.H(net1744));
 TIEHIx1_ASAP7_75t_R _35824__1745 (.H(net1745));
 TIEHIx1_ASAP7_75t_R _35825__1746 (.H(net1746));
 TIEHIx1_ASAP7_75t_R _35826__1747 (.H(net1747));
 TIEHIx1_ASAP7_75t_R _35827__1748 (.H(net1748));
 TIEHIx1_ASAP7_75t_R _35828__1749 (.H(net1749));
 TIEHIx1_ASAP7_75t_R _35829__1750 (.H(net1750));
 TIEHIx1_ASAP7_75t_R _35830__1751 (.H(net1751));
 TIEHIx1_ASAP7_75t_R _35831__1752 (.H(net1752));
 TIEHIx1_ASAP7_75t_R _35832__1753 (.H(net1753));
 TIEHIx1_ASAP7_75t_R _35833__1754 (.H(net1754));
 TIEHIx1_ASAP7_75t_R _35834__1755 (.H(net1755));
 TIEHIx1_ASAP7_75t_R _35835__1756 (.H(net1756));
 TIEHIx1_ASAP7_75t_R _35836__1757 (.H(net1757));
 TIEHIx1_ASAP7_75t_R _35837__1758 (.H(net1758));
 TIEHIx1_ASAP7_75t_R _35838__1759 (.H(net1759));
 TIEHIx1_ASAP7_75t_R _35839__1760 (.H(net1760));
 TIEHIx1_ASAP7_75t_R _35840__1761 (.H(net1761));
 TIEHIx1_ASAP7_75t_R _35841__1762 (.H(net1762));
 TIEHIx1_ASAP7_75t_R _35842__1763 (.H(net1763));
 TIEHIx1_ASAP7_75t_R _35843__1764 (.H(net1764));
 TIEHIx1_ASAP7_75t_R _35844__1765 (.H(net1765));
 TIEHIx1_ASAP7_75t_R _35845__1766 (.H(net1766));
 TIEHIx1_ASAP7_75t_R _35846__1767 (.H(net1767));
 TIEHIx1_ASAP7_75t_R _35847__1768 (.H(net1768));
 TIEHIx1_ASAP7_75t_R _35848__1769 (.H(net1769));
 TIEHIx1_ASAP7_75t_R _35849__1770 (.H(net1770));
 TIEHIx1_ASAP7_75t_R _35850__1771 (.H(net1771));
 TIEHIx1_ASAP7_75t_R _35851__1772 (.H(net1772));
 TIEHIx1_ASAP7_75t_R _35852__1773 (.H(net1773));
 TIEHIx1_ASAP7_75t_R _35853__1774 (.H(net1774));
 TIEHIx1_ASAP7_75t_R _35854__1775 (.H(net1775));
 TIEHIx1_ASAP7_75t_R _35855__1776 (.H(net1776));
 TIEHIx1_ASAP7_75t_R _35856__1777 (.H(net1777));
 TIEHIx1_ASAP7_75t_R _35857__1778 (.H(net1778));
 TIEHIx1_ASAP7_75t_R _35858__1779 (.H(net1779));
 TIEHIx1_ASAP7_75t_R _35859__1780 (.H(net1780));
 TIEHIx1_ASAP7_75t_R _35860__1781 (.H(net1781));
 TIEHIx1_ASAP7_75t_R _35861__1782 (.H(net1782));
 TIEHIx1_ASAP7_75t_R _35862__1783 (.H(net1783));
 TIEHIx1_ASAP7_75t_R _35863__1784 (.H(net1784));
 TIEHIx1_ASAP7_75t_R _35864__1785 (.H(net1785));
 TIEHIx1_ASAP7_75t_R _35865__1786 (.H(net1786));
 TIEHIx1_ASAP7_75t_R _35866__1787 (.H(net1787));
 TIEHIx1_ASAP7_75t_R _35867__1788 (.H(net1788));
 TIEHIx1_ASAP7_75t_R _35868__1789 (.H(net1789));
 TIEHIx1_ASAP7_75t_R _35869__1790 (.H(net1790));
 TIEHIx1_ASAP7_75t_R _35870__1791 (.H(net1791));
 TIEHIx1_ASAP7_75t_R _35871__1792 (.H(net1792));
 TIEHIx1_ASAP7_75t_R _35872__1793 (.H(net1793));
 TIEHIx1_ASAP7_75t_R _35873__1794 (.H(net1794));
 TIEHIx1_ASAP7_75t_R _35874__1795 (.H(net1795));
 TIEHIx1_ASAP7_75t_R _35875__1796 (.H(net1796));
 TIEHIx1_ASAP7_75t_R _35876__1797 (.H(net1797));
 TIEHIx1_ASAP7_75t_R _35877__1798 (.H(net1798));
 TIEHIx1_ASAP7_75t_R _35878__1799 (.H(net1799));
 TIEHIx1_ASAP7_75t_R _35879__1800 (.H(net1800));
 TIEHIx1_ASAP7_75t_R _35880__1801 (.H(net1801));
 TIEHIx1_ASAP7_75t_R _35881__1802 (.H(net1802));
 TIEHIx1_ASAP7_75t_R _35882__1803 (.H(net1803));
 TIEHIx1_ASAP7_75t_R _35883__1804 (.H(net1804));
 TIEHIx1_ASAP7_75t_R _35884__1805 (.H(net1805));
 TIEHIx1_ASAP7_75t_R _35885__1806 (.H(net1806));
 TIEHIx1_ASAP7_75t_R _35886__1807 (.H(net1807));
 TIEHIx1_ASAP7_75t_R _35887__1808 (.H(net1808));
 TIEHIx1_ASAP7_75t_R _35888__1809 (.H(net1809));
 TIEHIx1_ASAP7_75t_R _35889__1810 (.H(net1810));
 TIEHIx1_ASAP7_75t_R _35890__1811 (.H(net1811));
 TIEHIx1_ASAP7_75t_R _35891__1812 (.H(net1812));
 TIEHIx1_ASAP7_75t_R _35892__1813 (.H(net1813));
 TIEHIx1_ASAP7_75t_R _35893__1814 (.H(net1814));
 TIEHIx1_ASAP7_75t_R _35894__1815 (.H(net1815));
 TIEHIx1_ASAP7_75t_R _35895__1816 (.H(net1816));
 TIEHIx1_ASAP7_75t_R _35896__1817 (.H(net1817));
 TIEHIx1_ASAP7_75t_R _35897__1818 (.H(net1818));
 TIEHIx1_ASAP7_75t_R _35898__1819 (.H(net1819));
 TIEHIx1_ASAP7_75t_R _35899__1820 (.H(net1820));
 TIEHIx1_ASAP7_75t_R _35900__1821 (.H(net1821));
 TIEHIx1_ASAP7_75t_R _35901__1822 (.H(net1822));
 TIEHIx1_ASAP7_75t_R _35902__1823 (.H(net1823));
 TIEHIx1_ASAP7_75t_R _35903__1824 (.H(net1824));
 TIEHIx1_ASAP7_75t_R _35904__1825 (.H(net1825));
 TIEHIx1_ASAP7_75t_R _35905__1826 (.H(net1826));
 TIEHIx1_ASAP7_75t_R _35906__1827 (.H(net1827));
 TIEHIx1_ASAP7_75t_R _35907__1828 (.H(net1828));
 TIEHIx1_ASAP7_75t_R _35908__1829 (.H(net1829));
 TIEHIx1_ASAP7_75t_R _35909__1830 (.H(net1830));
 TIEHIx1_ASAP7_75t_R _35910__1831 (.H(net1831));
 TIEHIx1_ASAP7_75t_R _35911__1832 (.H(net1832));
 TIEHIx1_ASAP7_75t_R _35912__1833 (.H(net1833));
 TIEHIx1_ASAP7_75t_R _35913__1834 (.H(net1834));
 TIEHIx1_ASAP7_75t_R _35914__1835 (.H(net1835));
 TIEHIx1_ASAP7_75t_R _35915__1836 (.H(net1836));
 TIEHIx1_ASAP7_75t_R _35916__1837 (.H(net1837));
 TIEHIx1_ASAP7_75t_R _35917__1838 (.H(net1838));
 TIEHIx1_ASAP7_75t_R _35918__1839 (.H(net1839));
 TIEHIx1_ASAP7_75t_R _35919__1840 (.H(net1840));
 TIEHIx1_ASAP7_75t_R _35920__1841 (.H(net1841));
 TIEHIx1_ASAP7_75t_R _35921__1842 (.H(net1842));
 TIEHIx1_ASAP7_75t_R _35922__1843 (.H(net1843));
 TIEHIx1_ASAP7_75t_R _35923__1844 (.H(net1844));
 TIEHIx1_ASAP7_75t_R _35924__1845 (.H(net1845));
 TIEHIx1_ASAP7_75t_R _35925__1846 (.H(net1846));
 TIEHIx1_ASAP7_75t_R _35926__1847 (.H(net1847));
 TIEHIx1_ASAP7_75t_R _35927__1848 (.H(net1848));
 TIEHIx1_ASAP7_75t_R _35928__1849 (.H(net1849));
 TIEHIx1_ASAP7_75t_R _35929__1850 (.H(net1850));
 TIEHIx1_ASAP7_75t_R _35930__1851 (.H(net1851));
 TIEHIx1_ASAP7_75t_R _35931__1852 (.H(net1852));
 TIEHIx1_ASAP7_75t_R _35932__1853 (.H(net1853));
 TIEHIx1_ASAP7_75t_R _35933__1854 (.H(net1854));
 TIEHIx1_ASAP7_75t_R _35934__1855 (.H(net1855));
 TIEHIx1_ASAP7_75t_R _35935__1856 (.H(net1856));
 TIEHIx1_ASAP7_75t_R _35936__1857 (.H(net1857));
 TIEHIx1_ASAP7_75t_R _35937__1858 (.H(net1858));
 TIEHIx1_ASAP7_75t_R _35938__1859 (.H(net1859));
 TIEHIx1_ASAP7_75t_R _35939__1860 (.H(net1860));
 TIEHIx1_ASAP7_75t_R _35940__1861 (.H(net1861));
 TIEHIx1_ASAP7_75t_R _35941__1862 (.H(net1862));
 TIEHIx1_ASAP7_75t_R _35942__1863 (.H(net1863));
 TIEHIx1_ASAP7_75t_R _35943__1864 (.H(net1864));
 TIEHIx1_ASAP7_75t_R _35944__1865 (.H(net1865));
 TIEHIx1_ASAP7_75t_R _35945__1866 (.H(net1866));
 TIEHIx1_ASAP7_75t_R _35946__1867 (.H(net1867));
 TIEHIx1_ASAP7_75t_R _35947__1868 (.H(net1868));
 TIEHIx1_ASAP7_75t_R _35948__1869 (.H(net1869));
 TIEHIx1_ASAP7_75t_R _35949__1870 (.H(net1870));
 TIEHIx1_ASAP7_75t_R _35950__1871 (.H(net1871));
 TIEHIx1_ASAP7_75t_R _35951__1872 (.H(net1872));
 TIEHIx1_ASAP7_75t_R _35952__1873 (.H(net1873));
 TIEHIx1_ASAP7_75t_R _35953__1874 (.H(net1874));
 TIEHIx1_ASAP7_75t_R _35954__1875 (.H(net1875));
 TIEHIx1_ASAP7_75t_R _35955__1876 (.H(net1876));
 TIEHIx1_ASAP7_75t_R _35956__1877 (.H(net1877));
 TIEHIx1_ASAP7_75t_R _35957__1878 (.H(net1878));
 TIEHIx1_ASAP7_75t_R _35958__1879 (.H(net1879));
 TIEHIx1_ASAP7_75t_R _35959__1880 (.H(net1880));
 TIEHIx1_ASAP7_75t_R _35960__1881 (.H(net1881));
 TIEHIx1_ASAP7_75t_R _35961__1882 (.H(net1882));
 TIEHIx1_ASAP7_75t_R _35962__1883 (.H(net1883));
 TIEHIx1_ASAP7_75t_R _35963__1884 (.H(net1884));
 TIEHIx1_ASAP7_75t_R _35964__1885 (.H(net1885));
 TIEHIx1_ASAP7_75t_R _35965__1886 (.H(net1886));
 TIEHIx1_ASAP7_75t_R _35966__1887 (.H(net1887));
 TIEHIx1_ASAP7_75t_R _35967__1888 (.H(net1888));
 TIEHIx1_ASAP7_75t_R _35968__1889 (.H(net1889));
 TIEHIx1_ASAP7_75t_R _35969__1890 (.H(net1890));
 TIEHIx1_ASAP7_75t_R _35970__1891 (.H(net1891));
 TIEHIx1_ASAP7_75t_R _35971__1892 (.H(net1892));
 TIEHIx1_ASAP7_75t_R _35972__1893 (.H(net1893));
 TIEHIx1_ASAP7_75t_R _35973__1894 (.H(net1894));
 TIEHIx1_ASAP7_75t_R _35974__1895 (.H(net1895));
 TIEHIx1_ASAP7_75t_R _35975__1896 (.H(net1896));
 TIEHIx1_ASAP7_75t_R _35976__1897 (.H(net1897));
 TIEHIx1_ASAP7_75t_R _35977__1898 (.H(net1898));
 TIEHIx1_ASAP7_75t_R _35978__1899 (.H(net1899));
 TIEHIx1_ASAP7_75t_R _35979__1900 (.H(net1900));
 TIEHIx1_ASAP7_75t_R _35980__1901 (.H(net1901));
 TIEHIx1_ASAP7_75t_R _35981__1902 (.H(net1902));
 TIEHIx1_ASAP7_75t_R _35982__1903 (.H(net1903));
 TIEHIx1_ASAP7_75t_R _35983__1904 (.H(net1904));
 TIEHIx1_ASAP7_75t_R _35984__1905 (.H(net1905));
 TIEHIx1_ASAP7_75t_R _35985__1906 (.H(net1906));
 TIEHIx1_ASAP7_75t_R _35986__1907 (.H(net1907));
 TIEHIx1_ASAP7_75t_R _35987__1908 (.H(net1908));
 TIEHIx1_ASAP7_75t_R _35988__1909 (.H(net1909));
 TIEHIx1_ASAP7_75t_R _35989__1910 (.H(net1910));
 TIEHIx1_ASAP7_75t_R _35990__1911 (.H(net1911));
 TIEHIx1_ASAP7_75t_R _35991__1912 (.H(net1912));
 TIEHIx1_ASAP7_75t_R _35992__1913 (.H(net1913));
 TIEHIx1_ASAP7_75t_R _35993__1914 (.H(net1914));
 TIEHIx1_ASAP7_75t_R _35994__1915 (.H(net1915));
 TIEHIx1_ASAP7_75t_R _35995__1916 (.H(net1916));
 TIEHIx1_ASAP7_75t_R _35996__1917 (.H(net1917));
 TIEHIx1_ASAP7_75t_R _35997__1918 (.H(net1918));
 TIEHIx1_ASAP7_75t_R _35998__1919 (.H(net1919));
 TIEHIx1_ASAP7_75t_R _35999__1920 (.H(net1920));
 TIEHIx1_ASAP7_75t_R _36000__1921 (.H(net1921));
 TIEHIx1_ASAP7_75t_R _36001__1922 (.H(net1922));
 TIEHIx1_ASAP7_75t_R _36002__1923 (.H(net1923));
 TIEHIx1_ASAP7_75t_R _36003__1924 (.H(net1924));
 TIEHIx1_ASAP7_75t_R _36004__1925 (.H(net1925));
 TIEHIx1_ASAP7_75t_R _36005__1926 (.H(net1926));
 TIEHIx1_ASAP7_75t_R _36006__1927 (.H(net1927));
 TIEHIx1_ASAP7_75t_R _36007__1928 (.H(net1928));
 TIEHIx1_ASAP7_75t_R _36008__1929 (.H(net1929));
 TIEHIx1_ASAP7_75t_R _36009__1930 (.H(net1930));
 TIEHIx1_ASAP7_75t_R _36010__1931 (.H(net1931));
 TIEHIx1_ASAP7_75t_R _36011__1932 (.H(net1932));
 TIEHIx1_ASAP7_75t_R _36012__1933 (.H(net1933));
 TIEHIx1_ASAP7_75t_R _36013__1934 (.H(net1934));
 TIEHIx1_ASAP7_75t_R _36014__1935 (.H(net1935));
 TIEHIx1_ASAP7_75t_R _36015__1936 (.H(net1936));
 TIEHIx1_ASAP7_75t_R _36016__1937 (.H(net1937));
 TIEHIx1_ASAP7_75t_R _36017__1938 (.H(net1938));
 TIEHIx1_ASAP7_75t_R _36018__1939 (.H(net1939));
 TIEHIx1_ASAP7_75t_R _36019__1940 (.H(net1940));
 TIEHIx1_ASAP7_75t_R _36020__1941 (.H(net1941));
 TIEHIx1_ASAP7_75t_R _36021__1942 (.H(net1942));
 TIEHIx1_ASAP7_75t_R _36022__1943 (.H(net1943));
 TIEHIx1_ASAP7_75t_R _36023__1944 (.H(net1944));
 TIEHIx1_ASAP7_75t_R _36024__1945 (.H(net1945));
 TIEHIx1_ASAP7_75t_R _36025__1946 (.H(net1946));
 TIEHIx1_ASAP7_75t_R _36026__1947 (.H(net1947));
 TIEHIx1_ASAP7_75t_R _36027__1948 (.H(net1948));
 TIEHIx1_ASAP7_75t_R _36028__1949 (.H(net1949));
 TIEHIx1_ASAP7_75t_R _36029__1950 (.H(net1950));
 TIEHIx1_ASAP7_75t_R _36030__1951 (.H(net1951));
 TIEHIx1_ASAP7_75t_R _36031__1952 (.H(net1952));
 TIEHIx1_ASAP7_75t_R _36032__1953 (.H(net1953));
 TIEHIx1_ASAP7_75t_R _36033__1954 (.H(net1954));
 TIEHIx1_ASAP7_75t_R _36034__1955 (.H(net1955));
 TIEHIx1_ASAP7_75t_R _36035__1956 (.H(net1956));
 TIEHIx1_ASAP7_75t_R _36036__1957 (.H(net1957));
 TIEHIx1_ASAP7_75t_R _36037__1958 (.H(net1958));
 TIEHIx1_ASAP7_75t_R _36038__1959 (.H(net1959));
 TIEHIx1_ASAP7_75t_R _36039__1960 (.H(net1960));
 TIEHIx1_ASAP7_75t_R _36040__1961 (.H(net1961));
 TIEHIx1_ASAP7_75t_R _36041__1962 (.H(net1962));
 TIEHIx1_ASAP7_75t_R _36042__1963 (.H(net1963));
 TIEHIx1_ASAP7_75t_R _36043__1964 (.H(net1964));
 TIEHIx1_ASAP7_75t_R _36044__1965 (.H(net1965));
 TIEHIx1_ASAP7_75t_R _36045__1966 (.H(net1966));
 TIEHIx1_ASAP7_75t_R _36046__1967 (.H(net1967));
 TIEHIx1_ASAP7_75t_R _36047__1968 (.H(net1968));
 TIEHIx1_ASAP7_75t_R _36048__1969 (.H(net1969));
 TIEHIx1_ASAP7_75t_R _36049__1970 (.H(net1970));
 TIEHIx1_ASAP7_75t_R _36050__1971 (.H(net1971));
 TIEHIx1_ASAP7_75t_R _36051__1972 (.H(net1972));
 TIEHIx1_ASAP7_75t_R _36052__1973 (.H(net1973));
 TIEHIx1_ASAP7_75t_R _36053__1974 (.H(net1974));
 TIEHIx1_ASAP7_75t_R _36054__1975 (.H(net1975));
 TIEHIx1_ASAP7_75t_R _36055__1976 (.H(net1976));
 TIEHIx1_ASAP7_75t_R _36056__1977 (.H(net1977));
 TIEHIx1_ASAP7_75t_R _36057__1978 (.H(net1978));
 TIEHIx1_ASAP7_75t_R _36058__1979 (.H(net1979));
 TIEHIx1_ASAP7_75t_R _36059__1980 (.H(net1980));
 TIEHIx1_ASAP7_75t_R _36060__1981 (.H(net1981));
 TIEHIx1_ASAP7_75t_R _36061__1982 (.H(net1982));
 TIEHIx1_ASAP7_75t_R _36062__1983 (.H(net1983));
 TIEHIx1_ASAP7_75t_R _36063__1984 (.H(net1984));
 TIEHIx1_ASAP7_75t_R _36064__1985 (.H(net1985));
 TIEHIx1_ASAP7_75t_R _36065__1986 (.H(net1986));
 TIEHIx1_ASAP7_75t_R _36066__1987 (.H(net1987));
 TIEHIx1_ASAP7_75t_R _36067__1988 (.H(net1988));
 TIEHIx1_ASAP7_75t_R _36068__1989 (.H(net1989));
 TIEHIx1_ASAP7_75t_R _36069__1990 (.H(net1990));
 TIEHIx1_ASAP7_75t_R _36070__1991 (.H(net1991));
 TIEHIx1_ASAP7_75t_R _36071__1992 (.H(net1992));
 TIEHIx1_ASAP7_75t_R _36072__1993 (.H(net1993));
 TIEHIx1_ASAP7_75t_R _36073__1994 (.H(net1994));
 TIEHIx1_ASAP7_75t_R _36074__1995 (.H(net1995));
 TIEHIx1_ASAP7_75t_R _36075__1996 (.H(net1996));
 TIEHIx1_ASAP7_75t_R _36076__1997 (.H(net1997));
 TIEHIx1_ASAP7_75t_R _36077__1998 (.H(net1998));
 TIEHIx1_ASAP7_75t_R _36078__1999 (.H(net1999));
 TIEHIx1_ASAP7_75t_R _36079__2000 (.H(net2000));
 TIEHIx1_ASAP7_75t_R _36080__2001 (.H(net2001));
 TIEHIx1_ASAP7_75t_R _36081__2002 (.H(net2002));
 TIEHIx1_ASAP7_75t_R _36082__2003 (.H(net2003));
 TIEHIx1_ASAP7_75t_R _36083__2004 (.H(net2004));
 TIEHIx1_ASAP7_75t_R _36084__2005 (.H(net2005));
 TIEHIx1_ASAP7_75t_R _36085__2006 (.H(net2006));
 TIEHIx1_ASAP7_75t_R _36086__2007 (.H(net2007));
 TIEHIx1_ASAP7_75t_R _36087__2008 (.H(net2008));
 TIEHIx1_ASAP7_75t_R _36088__2009 (.H(net2009));
 TIEHIx1_ASAP7_75t_R _36089__2010 (.H(net2010));
 TIEHIx1_ASAP7_75t_R _36090__2011 (.H(net2011));
 TIEHIx1_ASAP7_75t_R _36091__2012 (.H(net2012));
 TIEHIx1_ASAP7_75t_R _36092__2013 (.H(net2013));
 TIEHIx1_ASAP7_75t_R _36093__2014 (.H(net2014));
 TIEHIx1_ASAP7_75t_R _36094__2015 (.H(net2015));
 TIEHIx1_ASAP7_75t_R _36095__2016 (.H(net2016));
 TIEHIx1_ASAP7_75t_R _36096__2017 (.H(net2017));
 TIEHIx1_ASAP7_75t_R _36097__2018 (.H(net2018));
 TIEHIx1_ASAP7_75t_R _36098__2019 (.H(net2019));
 TIEHIx1_ASAP7_75t_R _36099__2020 (.H(net2020));
 TIEHIx1_ASAP7_75t_R _36100__2021 (.H(net2021));
 TIEHIx1_ASAP7_75t_R _36101__2022 (.H(net2022));
 TIEHIx1_ASAP7_75t_R _36102__2023 (.H(net2023));
 TIEHIx1_ASAP7_75t_R _36103__2024 (.H(net2024));
 TIEHIx1_ASAP7_75t_R _36104__2025 (.H(net2025));
 TIEHIx1_ASAP7_75t_R _36105__2026 (.H(net2026));
 TIEHIx1_ASAP7_75t_R _36106__2027 (.H(net2027));
 TIEHIx1_ASAP7_75t_R _36107__2028 (.H(net2028));
 TIEHIx1_ASAP7_75t_R _36108__2029 (.H(net2029));
 TIEHIx1_ASAP7_75t_R _36109__2030 (.H(net2030));
 TIEHIx1_ASAP7_75t_R _36110__2031 (.H(net2031));
 TIEHIx1_ASAP7_75t_R _36111__2032 (.H(net2032));
 TIEHIx1_ASAP7_75t_R _36112__2033 (.H(net2033));
 TIEHIx1_ASAP7_75t_R _36113__2034 (.H(net2034));
 TIEHIx1_ASAP7_75t_R _36114__2035 (.H(net2035));
 TIEHIx1_ASAP7_75t_R _36115__2036 (.H(net2036));
 TIEHIx1_ASAP7_75t_R _36116__2037 (.H(net2037));
 TIEHIx1_ASAP7_75t_R _36117__2038 (.H(net2038));
 TIEHIx1_ASAP7_75t_R _36118__2039 (.H(net2039));
 TIEHIx1_ASAP7_75t_R _36119__2040 (.H(net2040));
 TIEHIx1_ASAP7_75t_R _36120__2041 (.H(net2041));
 TIEHIx1_ASAP7_75t_R _36121__2042 (.H(net2042));
 TIEHIx1_ASAP7_75t_R _36122__2043 (.H(net2043));
 TIEHIx1_ASAP7_75t_R _36123__2044 (.H(net2044));
 TIEHIx1_ASAP7_75t_R _36124__2045 (.H(net2045));
 TIEHIx1_ASAP7_75t_R _36125__2046 (.H(net2046));
 TIEHIx1_ASAP7_75t_R _36126__2047 (.H(net2047));
 TIEHIx1_ASAP7_75t_R _36127__2048 (.H(net2048));
 TIEHIx1_ASAP7_75t_R _36128__2049 (.H(net2049));
 TIEHIx1_ASAP7_75t_R _36129__2050 (.H(net2050));
 TIEHIx1_ASAP7_75t_R _36130__2051 (.H(net2051));
 TIEHIx1_ASAP7_75t_R _36131__2052 (.H(net2052));
 TIEHIx1_ASAP7_75t_R _36132__2053 (.H(net2053));
 TIEHIx1_ASAP7_75t_R _36133__2054 (.H(net2054));
 TIEHIx1_ASAP7_75t_R _36134__2055 (.H(net2055));
 TIEHIx1_ASAP7_75t_R _36135__2056 (.H(net2056));
 TIEHIx1_ASAP7_75t_R _36136__2057 (.H(net2057));
 TIEHIx1_ASAP7_75t_R _36137__2058 (.H(net2058));
 TIEHIx1_ASAP7_75t_R _36138__2059 (.H(net2059));
 TIEHIx1_ASAP7_75t_R _36139__2060 (.H(net2060));
 TIEHIx1_ASAP7_75t_R _36140__2061 (.H(net2061));
 TIEHIx1_ASAP7_75t_R _36141__2062 (.H(net2062));
 TIEHIx1_ASAP7_75t_R _36142__2063 (.H(net2063));
 TIEHIx1_ASAP7_75t_R _36143__2064 (.H(net2064));
 TIEHIx1_ASAP7_75t_R _36144__2065 (.H(net2065));
 TIEHIx1_ASAP7_75t_R _36145__2066 (.H(net2066));
 TIEHIx1_ASAP7_75t_R _36146__2067 (.H(net2067));
 TIEHIx1_ASAP7_75t_R _36147__2068 (.H(net2068));
 TIEHIx1_ASAP7_75t_R _36148__2069 (.H(net2069));
 TIEHIx1_ASAP7_75t_R _36149__2070 (.H(net2070));
 TIEHIx1_ASAP7_75t_R _36150__2071 (.H(net2071));
 TIEHIx1_ASAP7_75t_R _36151__2072 (.H(net2072));
 TIEHIx1_ASAP7_75t_R _36152__2073 (.H(net2073));
 TIEHIx1_ASAP7_75t_R _36153__2074 (.H(net2074));
 TIEHIx1_ASAP7_75t_R _36154__2075 (.H(net2075));
 TIEHIx1_ASAP7_75t_R _36155__2076 (.H(net2076));
 TIEHIx1_ASAP7_75t_R _36156__2077 (.H(net2077));
 TIEHIx1_ASAP7_75t_R _36157__2078 (.H(net2078));
 TIEHIx1_ASAP7_75t_R _36158__2079 (.H(net2079));
 TIEHIx1_ASAP7_75t_R _36159__2080 (.H(net2080));
 TIEHIx1_ASAP7_75t_R _36160__2081 (.H(net2081));
 TIEHIx1_ASAP7_75t_R _36161__2082 (.H(net2082));
 TIEHIx1_ASAP7_75t_R _36162__2083 (.H(net2083));
 TIEHIx1_ASAP7_75t_R _36163__2084 (.H(net2084));
 TIEHIx1_ASAP7_75t_R _36164__2085 (.H(net2085));
 TIEHIx1_ASAP7_75t_R _36165__2086 (.H(net2086));
 TIEHIx1_ASAP7_75t_R _36166__2087 (.H(net2087));
 TIEHIx1_ASAP7_75t_R _36167__2088 (.H(net2088));
 TIEHIx1_ASAP7_75t_R _36168__2089 (.H(net2089));
 TIEHIx1_ASAP7_75t_R _36169__2090 (.H(net2090));
 TIEHIx1_ASAP7_75t_R _36170__2091 (.H(net2091));
 TIEHIx1_ASAP7_75t_R _36171__2092 (.H(net2092));
 TIEHIx1_ASAP7_75t_R _36172__2093 (.H(net2093));
 TIEHIx1_ASAP7_75t_R _36173__2094 (.H(net2094));
 TIEHIx1_ASAP7_75t_R _36174__2095 (.H(net2095));
 TIEHIx1_ASAP7_75t_R _36175__2096 (.H(net2096));
 TIEHIx1_ASAP7_75t_R _36176__2097 (.H(net2097));
 TIEHIx1_ASAP7_75t_R _36177__2098 (.H(net2098));
 TIEHIx1_ASAP7_75t_R _36178__2099 (.H(net2099));
 TIEHIx1_ASAP7_75t_R _36179__2100 (.H(net2100));
 TIEHIx1_ASAP7_75t_R _36180__2101 (.H(net2101));
 TIEHIx1_ASAP7_75t_R _36181__2102 (.H(net2102));
 TIEHIx1_ASAP7_75t_R _36183__2103 (.H(net2103));
 TIEHIx1_ASAP7_75t_R _36184__2104 (.H(net2104));
 TIEHIx1_ASAP7_75t_R _36185__2105 (.H(net2105));
 TIEHIx1_ASAP7_75t_R _36186__2106 (.H(net2106));
 TIEHIx1_ASAP7_75t_R _36187__2107 (.H(net2107));
 TIEHIx1_ASAP7_75t_R _36188__2108 (.H(net2108));
 TIEHIx1_ASAP7_75t_R _36222__2109 (.H(net2109));
 TIEHIx1_ASAP7_75t_R _36223__2110 (.H(net2110));
 TIEHIx1_ASAP7_75t_R _36224__2111 (.H(net2111));
 TIEHIx1_ASAP7_75t_R _36292__2112 (.H(net2112));
 TIEHIx1_ASAP7_75t_R _36325__2113 (.H(net2113));
 BUFx4_ASAP7_75t_R clkbuf_leaf_1_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_1_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_2_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_2_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_3_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_3_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_4_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_4_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_5_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_5_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_6_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_6_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_7_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_7_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_8_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_8_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_9_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_9_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_10_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_10_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_11_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_11_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_12_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_12_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_13_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_13_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_14_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_14_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_15_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_15_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_16_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_16_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_17_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_17_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_18_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_18_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_19_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_19_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_20_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_20_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_21_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_21_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_22_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_22_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_23_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_23_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_24_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_24_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_25_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_25_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_26_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_26_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_27_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_27_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_28_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_28_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_29_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_29_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_30_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_30_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_31_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_31_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_32_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_32_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_33_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_33_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_0_clk_i (.A(clk_i),
    .Y(clknet_0_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_2_0__f_clk_i (.A(clknet_0_clk_i),
    .Y(clknet_2_0__leaf_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_2_1__f_clk_i (.A(clknet_0_clk_i),
    .Y(clknet_2_1__leaf_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_2_2__f_clk_i (.A(clknet_0_clk_i),
    .Y(clknet_2_2__leaf_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_2_3__f_clk_i (.A(clknet_0_clk_i),
    .Y(clknet_2_3__leaf_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_10_clk_i (.A(clknet_leaf_0_clk_i),
    .Y(clknet_level_0_1_10_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_11_clk_i (.A(clknet_level_0_1_10_clk_i),
    .Y(clknet_level_1_1_11_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_12_clk_i (.A(clknet_level_1_1_11_clk_i),
    .Y(clknet_level_2_1_12_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_13_clk_i (.A(clknet_level_2_1_12_clk_i),
    .Y(clknet_level_3_1_13_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_24_clk_i (.A(clknet_leaf_1_clk_i),
    .Y(clknet_level_0_1_24_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_25_clk_i (.A(clknet_level_0_1_24_clk_i),
    .Y(clknet_level_1_1_25_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_26_clk_i (.A(clknet_level_1_1_25_clk_i),
    .Y(clknet_level_2_1_26_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_27_clk_i (.A(clknet_level_2_1_26_clk_i),
    .Y(clknet_level_3_1_27_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_38_clk_i (.A(clknet_leaf_2_clk_i),
    .Y(clknet_level_0_1_38_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_39_clk_i (.A(clknet_level_0_1_38_clk_i),
    .Y(clknet_level_1_1_39_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_310_clk_i (.A(clknet_level_1_1_39_clk_i),
    .Y(clknet_level_2_1_310_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_311_clk_i (.A(clknet_level_2_1_310_clk_i),
    .Y(clknet_level_3_1_311_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_412_clk_i (.A(clknet_leaf_3_clk_i),
    .Y(clknet_level_0_1_412_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_413_clk_i (.A(clknet_level_0_1_412_clk_i),
    .Y(clknet_level_1_1_413_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_414_clk_i (.A(clknet_level_1_1_413_clk_i),
    .Y(clknet_level_2_1_414_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_415_clk_i (.A(clknet_level_2_1_414_clk_i),
    .Y(clknet_level_3_1_415_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_516_clk_i (.A(clknet_leaf_4_clk_i),
    .Y(clknet_level_0_1_516_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_517_clk_i (.A(clknet_level_0_1_516_clk_i),
    .Y(clknet_level_1_1_517_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_518_clk_i (.A(clknet_level_1_1_517_clk_i),
    .Y(clknet_level_2_1_518_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_519_clk_i (.A(clknet_level_2_1_518_clk_i),
    .Y(clknet_level_3_1_519_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_620_clk_i (.A(clknet_leaf_5_clk_i),
    .Y(clknet_level_0_1_620_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_621_clk_i (.A(clknet_level_0_1_620_clk_i),
    .Y(clknet_level_1_1_621_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_622_clk_i (.A(clknet_level_1_1_621_clk_i),
    .Y(clknet_level_2_1_622_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_623_clk_i (.A(clknet_level_2_1_622_clk_i),
    .Y(clknet_level_3_1_623_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_724_clk_i (.A(clknet_leaf_6_clk_i),
    .Y(clknet_level_0_1_724_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_725_clk_i (.A(clknet_level_0_1_724_clk_i),
    .Y(clknet_level_1_1_725_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_726_clk_i (.A(clknet_level_1_1_725_clk_i),
    .Y(clknet_level_2_1_726_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_727_clk_i (.A(clknet_level_2_1_726_clk_i),
    .Y(clknet_level_3_1_727_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_828_clk_i (.A(clknet_leaf_7_clk_i),
    .Y(clknet_level_0_1_828_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_829_clk_i (.A(clknet_level_0_1_828_clk_i),
    .Y(clknet_level_1_1_829_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_830_clk_i (.A(clknet_level_1_1_829_clk_i),
    .Y(clknet_level_2_1_830_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_831_clk_i (.A(clknet_level_2_1_830_clk_i),
    .Y(clknet_level_3_1_831_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_932_clk_i (.A(clknet_leaf_8_clk_i),
    .Y(clknet_level_0_1_932_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_933_clk_i (.A(clknet_level_0_1_932_clk_i),
    .Y(clknet_level_1_1_933_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_934_clk_i (.A(clknet_level_1_1_933_clk_i),
    .Y(clknet_level_2_1_934_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_935_clk_i (.A(clknet_level_2_1_934_clk_i),
    .Y(clknet_level_3_1_935_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1036_clk_i (.A(clknet_leaf_9_clk_i),
    .Y(clknet_level_0_1_1036_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1037_clk_i (.A(clknet_level_0_1_1036_clk_i),
    .Y(clknet_level_1_1_1037_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1038_clk_i (.A(clknet_level_1_1_1037_clk_i),
    .Y(clknet_level_2_1_1038_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1039_clk_i (.A(clknet_level_2_1_1038_clk_i),
    .Y(clknet_level_3_1_1039_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1140_clk_i (.A(clknet_leaf_10_clk_i),
    .Y(clknet_level_0_1_1140_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1141_clk_i (.A(clknet_level_0_1_1140_clk_i),
    .Y(clknet_level_1_1_1141_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1142_clk_i (.A(clknet_level_1_1_1141_clk_i),
    .Y(clknet_level_2_1_1142_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1143_clk_i (.A(clknet_level_2_1_1142_clk_i),
    .Y(clknet_level_3_1_1143_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1244_clk_i (.A(clknet_leaf_11_clk_i),
    .Y(clknet_level_0_1_1244_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1245_clk_i (.A(clknet_level_0_1_1244_clk_i),
    .Y(clknet_level_1_1_1245_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1246_clk_i (.A(clknet_level_1_1_1245_clk_i),
    .Y(clknet_level_2_1_1246_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1247_clk_i (.A(clknet_level_2_1_1246_clk_i),
    .Y(clknet_level_3_1_1247_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1348_clk_i (.A(clknet_leaf_12_clk_i),
    .Y(clknet_level_0_1_1348_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1349_clk_i (.A(clknet_level_0_1_1348_clk_i),
    .Y(clknet_level_1_1_1349_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1350_clk_i (.A(clknet_level_1_1_1349_clk_i),
    .Y(clknet_level_2_1_1350_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1351_clk_i (.A(clknet_level_2_1_1350_clk_i),
    .Y(clknet_level_3_1_1351_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1452_clk_i (.A(clknet_leaf_13_clk_i),
    .Y(clknet_level_0_1_1452_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1453_clk_i (.A(clknet_level_0_1_1452_clk_i),
    .Y(clknet_level_1_1_1453_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1454_clk_i (.A(clknet_level_1_1_1453_clk_i),
    .Y(clknet_level_2_1_1454_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1455_clk_i (.A(clknet_level_2_1_1454_clk_i),
    .Y(clknet_level_3_1_1455_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1556_clk_i (.A(clknet_leaf_14_clk_i),
    .Y(clknet_level_0_1_1556_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1557_clk_i (.A(clknet_level_0_1_1556_clk_i),
    .Y(clknet_level_1_1_1557_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1558_clk_i (.A(clknet_level_1_1_1557_clk_i),
    .Y(clknet_level_2_1_1558_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1559_clk_i (.A(clknet_level_2_1_1558_clk_i),
    .Y(clknet_level_3_1_1559_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1660_clk_i (.A(clknet_leaf_15_clk_i),
    .Y(clknet_level_0_1_1660_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1661_clk_i (.A(clknet_level_0_1_1660_clk_i),
    .Y(clknet_level_1_1_1661_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1662_clk_i (.A(clknet_level_1_1_1661_clk_i),
    .Y(clknet_level_2_1_1662_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1663_clk_i (.A(clknet_level_2_1_1662_clk_i),
    .Y(clknet_level_3_1_1663_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1764_clk_i (.A(clknet_leaf_16_clk_i),
    .Y(clknet_level_0_1_1764_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1765_clk_i (.A(clknet_level_0_1_1764_clk_i),
    .Y(clknet_level_1_1_1765_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1766_clk_i (.A(clknet_level_1_1_1765_clk_i),
    .Y(clknet_level_2_1_1766_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1767_clk_i (.A(clknet_level_2_1_1766_clk_i),
    .Y(clknet_level_3_1_1767_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1868_clk_i (.A(clknet_leaf_17_clk_i),
    .Y(clknet_level_0_1_1868_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1869_clk_i (.A(clknet_level_0_1_1868_clk_i),
    .Y(clknet_level_1_1_1869_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1870_clk_i (.A(clknet_level_1_1_1869_clk_i),
    .Y(clknet_level_2_1_1870_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1871_clk_i (.A(clknet_level_2_1_1870_clk_i),
    .Y(clknet_level_3_1_1871_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1972_clk_i (.A(clknet_leaf_18_clk_i),
    .Y(clknet_level_0_1_1972_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1973_clk_i (.A(clknet_level_0_1_1972_clk_i),
    .Y(clknet_level_1_1_1973_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1974_clk_i (.A(clknet_level_1_1_1973_clk_i),
    .Y(clknet_level_2_1_1974_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1975_clk_i (.A(clknet_level_2_1_1974_clk_i),
    .Y(clknet_level_3_1_1975_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_2076_clk_i (.A(clknet_leaf_19_clk_i),
    .Y(clknet_level_0_1_2076_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_2077_clk_i (.A(clknet_level_0_1_2076_clk_i),
    .Y(clknet_level_1_1_2077_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_2078_clk_i (.A(clknet_level_1_1_2077_clk_i),
    .Y(clknet_level_2_1_2078_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_2079_clk_i (.A(clknet_level_2_1_2078_clk_i),
    .Y(clknet_level_3_1_2079_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_2180_clk_i (.A(clknet_leaf_20_clk_i),
    .Y(clknet_level_0_1_2180_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_2181_clk_i (.A(clknet_level_0_1_2180_clk_i),
    .Y(clknet_level_1_1_2181_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_2182_clk_i (.A(clknet_level_1_1_2181_clk_i),
    .Y(clknet_level_2_1_2182_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_2183_clk_i (.A(clknet_level_2_1_2182_clk_i),
    .Y(clknet_level_3_1_2183_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_2284_clk_i (.A(clknet_leaf_21_clk_i),
    .Y(clknet_level_0_1_2284_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_2285_clk_i (.A(clknet_level_0_1_2284_clk_i),
    .Y(clknet_level_1_1_2285_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_2286_clk_i (.A(clknet_level_1_1_2285_clk_i),
    .Y(clknet_level_2_1_2286_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_2287_clk_i (.A(clknet_level_2_1_2286_clk_i),
    .Y(clknet_level_3_1_2287_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_2388_clk_i (.A(clknet_leaf_22_clk_i),
    .Y(clknet_level_0_1_2388_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_2389_clk_i (.A(clknet_level_0_1_2388_clk_i),
    .Y(clknet_level_1_1_2389_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_2390_clk_i (.A(clknet_level_1_1_2389_clk_i),
    .Y(clknet_level_2_1_2390_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_2391_clk_i (.A(clknet_level_2_1_2390_clk_i),
    .Y(clknet_level_3_1_2391_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_2492_clk_i (.A(clknet_leaf_23_clk_i),
    .Y(clknet_level_0_1_2492_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_2493_clk_i (.A(clknet_level_0_1_2492_clk_i),
    .Y(clknet_level_1_1_2493_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_2494_clk_i (.A(clknet_level_1_1_2493_clk_i),
    .Y(clknet_level_2_1_2494_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_2495_clk_i (.A(clknet_level_2_1_2494_clk_i),
    .Y(clknet_level_3_1_2495_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_2596_clk_i (.A(clknet_leaf_24_clk_i),
    .Y(clknet_level_0_1_2596_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_2597_clk_i (.A(clknet_level_0_1_2596_clk_i),
    .Y(clknet_level_1_1_2597_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_2598_clk_i (.A(clknet_level_1_1_2597_clk_i),
    .Y(clknet_level_2_1_2598_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_2599_clk_i (.A(clknet_level_2_1_2598_clk_i),
    .Y(clknet_level_3_1_2599_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_26100_clk_i (.A(clknet_leaf_25_clk_i),
    .Y(clknet_level_0_1_26100_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_26101_clk_i (.A(clknet_level_0_1_26100_clk_i),
    .Y(clknet_level_1_1_26101_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_26102_clk_i (.A(clknet_level_1_1_26101_clk_i),
    .Y(clknet_level_2_1_26102_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_26103_clk_i (.A(clknet_level_2_1_26102_clk_i),
    .Y(clknet_level_3_1_26103_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_27104_clk_i (.A(clknet_leaf_26_clk_i),
    .Y(clknet_level_0_1_27104_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_27105_clk_i (.A(clknet_level_0_1_27104_clk_i),
    .Y(clknet_level_1_1_27105_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_27106_clk_i (.A(clknet_level_1_1_27105_clk_i),
    .Y(clknet_level_2_1_27106_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_27107_clk_i (.A(clknet_level_2_1_27106_clk_i),
    .Y(clknet_level_3_1_27107_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_28108_clk_i (.A(clknet_leaf_27_clk_i),
    .Y(clknet_level_0_1_28108_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_28109_clk_i (.A(clknet_level_0_1_28108_clk_i),
    .Y(clknet_level_1_1_28109_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_28110_clk_i (.A(clknet_level_1_1_28109_clk_i),
    .Y(clknet_level_2_1_28110_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_28111_clk_i (.A(clknet_level_2_1_28110_clk_i),
    .Y(clknet_level_3_1_28111_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_29112_clk_i (.A(clknet_leaf_28_clk_i),
    .Y(clknet_level_0_1_29112_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_29113_clk_i (.A(clknet_level_0_1_29112_clk_i),
    .Y(clknet_level_1_1_29113_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_29114_clk_i (.A(clknet_level_1_1_29113_clk_i),
    .Y(clknet_level_2_1_29114_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_29115_clk_i (.A(clknet_level_2_1_29114_clk_i),
    .Y(clknet_level_3_1_29115_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_30116_clk_i (.A(clknet_leaf_29_clk_i),
    .Y(clknet_level_0_1_30116_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_30117_clk_i (.A(clknet_level_0_1_30116_clk_i),
    .Y(clknet_level_1_1_30117_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_30118_clk_i (.A(clknet_level_1_1_30117_clk_i),
    .Y(clknet_level_2_1_30118_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_30119_clk_i (.A(clknet_level_2_1_30118_clk_i),
    .Y(clknet_level_3_1_30119_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_31120_clk_i (.A(clknet_leaf_30_clk_i),
    .Y(clknet_level_0_1_31120_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_31121_clk_i (.A(clknet_level_0_1_31120_clk_i),
    .Y(clknet_level_1_1_31121_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_31122_clk_i (.A(clknet_level_1_1_31121_clk_i),
    .Y(clknet_level_2_1_31122_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_31123_clk_i (.A(clknet_level_2_1_31122_clk_i),
    .Y(clknet_level_3_1_31123_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_32124_clk_i (.A(clknet_leaf_31_clk_i),
    .Y(clknet_level_0_1_32124_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_32125_clk_i (.A(clknet_level_0_1_32124_clk_i),
    .Y(clknet_level_1_1_32125_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_32126_clk_i (.A(clknet_level_1_1_32125_clk_i),
    .Y(clknet_level_2_1_32126_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_32127_clk_i (.A(clknet_level_2_1_32126_clk_i),
    .Y(clknet_level_3_1_32127_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_33128_clk_i (.A(clknet_leaf_32_clk_i),
    .Y(clknet_level_0_1_33128_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_33129_clk_i (.A(clknet_level_0_1_33128_clk_i),
    .Y(clknet_level_1_1_33129_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_33130_clk_i (.A(clknet_level_1_1_33129_clk_i),
    .Y(clknet_level_2_1_33130_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_33131_clk_i (.A(clknet_level_2_1_33130_clk_i),
    .Y(clknet_level_3_1_33131_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_34132_clk_i (.A(clknet_leaf_33_clk_i),
    .Y(clknet_level_0_1_34132_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_34133_clk_i (.A(clknet_level_0_1_34132_clk_i),
    .Y(clknet_level_1_1_34133_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_34134_clk_i (.A(clknet_level_1_1_34133_clk_i),
    .Y(clknet_level_2_1_34134_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_34135_clk_i (.A(clknet_level_2_1_34134_clk_i),
    .Y(clknet_level_3_1_34135_clk_i));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_0_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_0_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_1_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_1_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_2_core_clock_gate_i.clk_o  (.A(\clknet_2_2__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_2_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_3_core_clock_gate_i.clk_o  (.A(\clknet_2_2__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_3_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_4_core_clock_gate_i.clk_o  (.A(\clknet_2_2__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_4_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_5_core_clock_gate_i.clk_o  (.A(\clknet_2_2__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_5_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_6_core_clock_gate_i.clk_o  (.A(\clknet_2_2__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_6_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_7_core_clock_gate_i.clk_o  (.A(\clknet_2_2__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_7_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_8_core_clock_gate_i.clk_o  (.A(\clknet_2_3__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_8_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_9_core_clock_gate_i.clk_o  (.A(\clknet_2_3__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_9_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_10_core_clock_gate_i.clk_o  (.A(\clknet_2_3__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_10_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_11_core_clock_gate_i.clk_o  (.A(\clknet_2_3__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_11_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_12_core_clock_gate_i.clk_o  (.A(\clknet_2_3__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_12_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_13_core_clock_gate_i.clk_o  (.A(\clknet_2_3__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_13_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_14_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_14_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_15_core_clock_gate_i.clk_o  (.A(\clknet_2_3__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_15_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_16_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_16_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_17_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_17_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_18_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_18_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_19_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_19_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_20_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_20_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_21_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_21_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_22_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_22_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_23_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_23_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_24_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_24_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_25_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_25_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_26_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_26_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_27_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_27_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_28_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_28_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_29_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_29_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_30_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_30_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_31_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_31_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_0_core_clock_gate_i.clk_o  (.A(\core_clock_gate_i.clk_o ),
    .Y(\clknet_0_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_2_0__f_core_clock_gate_i.clk_o  (.A(\clknet_0_core_clock_gate_i.clk_o ),
    .Y(\clknet_2_0__leaf_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_2_1__f_core_clock_gate_i.clk_o  (.A(\clknet_0_core_clock_gate_i.clk_o ),
    .Y(\clknet_2_1__leaf_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_2_2__f_core_clock_gate_i.clk_o  (.A(\clknet_0_core_clock_gate_i.clk_o ),
    .Y(\clknet_2_2__leaf_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_2_3__f_core_clock_gate_i.clk_o  (.A(\clknet_0_core_clock_gate_i.clk_o ),
    .Y(\clknet_2_3__leaf_core_clock_gate_i.clk_o ));
 BUFx2_ASAP7_75t_R rebuffer1 (.A(net170),
    .Y(net2114));
 BUFx3_ASAP7_75t_R rebuffer2 (.A(net170),
    .Y(net2115));
 BUFx2_ASAP7_75t_R rebuffer3 (.A(net2115),
    .Y(net2116));
 BUFx3_ASAP7_75t_R rebuffer4 (.A(net2116),
    .Y(net2117));
 BUFx3_ASAP7_75t_R rebuffer5 (.A(net2115),
    .Y(net2118));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_420 ();
 DECAPx1_ASAP7_75t_R FILLER_0_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_446 ();
 FILLER_ASAP7_75t_R FILLER_0_452 ();
 FILLER_ASAP7_75t_R FILLER_0_460 ();
 FILLER_ASAP7_75t_R FILLER_0_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_473 ();
 FILLER_ASAP7_75t_R FILLER_0_479 ();
 FILLER_ASAP7_75t_R FILLER_0_488 ();
 DECAPx1_ASAP7_75t_R FILLER_0_496 ();
 FILLER_ASAP7_75t_R FILLER_0_507 ();
 FILLER_ASAP7_75t_R FILLER_0_515 ();
 FILLER_ASAP7_75t_R FILLER_0_523 ();
 FILLER_ASAP7_75t_R FILLER_0_531 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_0_541 ();
 FILLER_ASAP7_75t_R FILLER_0_550 ();
 FILLER_ASAP7_75t_R FILLER_0_560 ();
 FILLER_ASAP7_75t_R FILLER_0_568 ();
 FILLER_ASAP7_75t_R FILLER_0_576 ();
 FILLER_ASAP7_75t_R FILLER_0_583 ();
 FILLER_ASAP7_75t_R FILLER_0_590 ();
 DECAPx2_ASAP7_75t_R FILLER_0_600 ();
 FILLER_ASAP7_75t_R FILLER_0_606 ();
 DECAPx2_ASAP7_75t_R FILLER_0_614 ();
 DECAPx1_ASAP7_75t_R FILLER_0_627 ();
 FILLER_ASAP7_75t_R FILLER_0_636 ();
 FILLER_ASAP7_75t_R FILLER_0_643 ();
 FILLER_ASAP7_75t_R FILLER_0_650 ();
 FILLER_ASAP7_75t_R FILLER_0_657 ();
 DECAPx1_ASAP7_75t_R FILLER_0_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_670 ();
 FILLER_ASAP7_75t_R FILLER_0_677 ();
 FILLER_ASAP7_75t_R FILLER_0_685 ();
 FILLER_ASAP7_75t_R FILLER_0_693 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_0_702 ();
 DECAPx1_ASAP7_75t_R FILLER_0_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_715 ();
 FILLER_ASAP7_75t_R FILLER_0_721 ();
 DECAPx1_ASAP7_75t_R FILLER_0_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_732 ();
 FILLER_ASAP7_75t_R FILLER_0_738 ();
 FILLER_ASAP7_75t_R FILLER_0_747 ();
 FILLER_ASAP7_75t_R FILLER_0_755 ();
 FILLER_ASAP7_75t_R FILLER_0_763 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_0_770 ();
 FILLER_ASAP7_75t_R FILLER_0_778 ();
 DECAPx2_ASAP7_75t_R FILLER_0_785 ();
 FILLER_ASAP7_75t_R FILLER_0_791 ();
 FILLER_ASAP7_75t_R FILLER_0_798 ();
 DECAPx2_ASAP7_75t_R FILLER_0_807 ();
 FILLER_ASAP7_75t_R FILLER_0_819 ();
 DECAPx2_ASAP7_75t_R FILLER_0_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_832 ();
 FILLER_ASAP7_75t_R FILLER_0_840 ();
 FILLER_ASAP7_75t_R FILLER_0_848 ();
 DECAPx2_ASAP7_75t_R FILLER_0_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_862 ();
 FILLER_ASAP7_75t_R FILLER_0_870 ();
 FILLER_ASAP7_75t_R FILLER_0_878 ();
 FILLER_ASAP7_75t_R FILLER_0_885 ();
 FILLER_ASAP7_75t_R FILLER_0_894 ();
 FILLER_ASAP7_75t_R FILLER_0_902 ();
 FILLER_ASAP7_75t_R FILLER_0_909 ();
 DECAPx2_ASAP7_75t_R FILLER_0_916 ();
 FILLER_ASAP7_75t_R FILLER_0_922 ();
 DECAPx2_ASAP7_75t_R FILLER_0_926 ();
 FILLER_ASAP7_75t_R FILLER_0_932 ();
 FILLER_ASAP7_75t_R FILLER_0_940 ();
 DECAPx1_ASAP7_75t_R FILLER_0_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_951 ();
 FILLER_ASAP7_75t_R FILLER_0_959 ();
 DECAPx2_ASAP7_75t_R FILLER_0_967 ();
 FILLER_ASAP7_75t_R FILLER_0_973 ();
 FILLER_ASAP7_75t_R FILLER_0_982 ();
 FILLER_ASAP7_75t_R FILLER_0_990 ();
 DECAPx1_ASAP7_75t_R FILLER_0_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1001 ();
 FILLER_ASAP7_75t_R FILLER_0_1009 ();
 FILLER_ASAP7_75t_R FILLER_0_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_1077 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1099 ();
 FILLER_ASAP7_75t_R FILLER_0_1109 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1122 ();
 FILLER_ASAP7_75t_R FILLER_0_1130 ();
 FILLER_ASAP7_75t_R FILLER_0_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_1145 ();
 FILLER_ASAP7_75t_R FILLER_0_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1159 ();
 FILLER_ASAP7_75t_R FILLER_0_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1208 ();
 FILLER_ASAP7_75t_R FILLER_0_1221 ();
 FILLER_ASAP7_75t_R FILLER_0_1229 ();
 FILLER_ASAP7_75t_R FILLER_0_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1353 ();
 FILLER_ASAP7_75t_R FILLER_0_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_1_46 ();
 DECAPx10_ASAP7_75t_R FILLER_1_68 ();
 DECAPx10_ASAP7_75t_R FILLER_1_90 ();
 DECAPx10_ASAP7_75t_R FILLER_1_112 ();
 DECAPx10_ASAP7_75t_R FILLER_1_134 ();
 DECAPx10_ASAP7_75t_R FILLER_1_156 ();
 DECAPx10_ASAP7_75t_R FILLER_1_178 ();
 DECAPx10_ASAP7_75t_R FILLER_1_200 ();
 DECAPx10_ASAP7_75t_R FILLER_1_222 ();
 DECAPx10_ASAP7_75t_R FILLER_1_244 ();
 DECAPx10_ASAP7_75t_R FILLER_1_266 ();
 DECAPx10_ASAP7_75t_R FILLER_1_288 ();
 DECAPx10_ASAP7_75t_R FILLER_1_310 ();
 DECAPx10_ASAP7_75t_R FILLER_1_332 ();
 DECAPx10_ASAP7_75t_R FILLER_1_354 ();
 DECAPx10_ASAP7_75t_R FILLER_1_376 ();
 DECAPx10_ASAP7_75t_R FILLER_1_398 ();
 DECAPx10_ASAP7_75t_R FILLER_1_420 ();
 DECAPx1_ASAP7_75t_R FILLER_1_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_446 ();
 DECAPx1_ASAP7_75t_R FILLER_1_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_471 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_1_492 ();
 FILLER_ASAP7_75t_R FILLER_1_515 ();
 FILLER_ASAP7_75t_R FILLER_1_537 ();
 FILLER_ASAP7_75t_R FILLER_1_546 ();
 FILLER_ASAP7_75t_R FILLER_1_553 ();
 FILLER_ASAP7_75t_R FILLER_1_562 ();
 DECAPx2_ASAP7_75t_R FILLER_1_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_576 ();
 FILLER_ASAP7_75t_R FILLER_1_584 ();
 DECAPx2_ASAP7_75t_R FILLER_1_592 ();
 FILLER_ASAP7_75t_R FILLER_1_598 ();
 FILLER_ASAP7_75t_R FILLER_1_607 ();
 FILLER_ASAP7_75t_R FILLER_1_614 ();
 DECAPx1_ASAP7_75t_R FILLER_1_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_640 ();
 FILLER_ASAP7_75t_R FILLER_1_648 ();
 DECAPx2_ASAP7_75t_R FILLER_1_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_676 ();
 DECAPx1_ASAP7_75t_R FILLER_1_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_688 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_1_709 ();
 FILLER_ASAP7_75t_R FILLER_1_715 ();
 FILLER_ASAP7_75t_R FILLER_1_724 ();
 DECAPx2_ASAP7_75t_R FILLER_1_732 ();
 DECAPx2_ASAP7_75t_R FILLER_1_758 ();
 FILLER_ASAP7_75t_R FILLER_1_771 ();
 DECAPx2_ASAP7_75t_R FILLER_1_780 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_1_786 ();
 FILLER_ASAP7_75t_R FILLER_1_809 ();
 FILLER_ASAP7_75t_R FILLER_1_817 ();
 DECAPx1_ASAP7_75t_R FILLER_1_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_829 ();
 DECAPx2_ASAP7_75t_R FILLER_1_850 ();
 FILLER_ASAP7_75t_R FILLER_1_856 ();
 DECAPx1_ASAP7_75t_R FILLER_1_878 ();
 DECAPx2_ASAP7_75t_R FILLER_1_902 ();
 FILLER_ASAP7_75t_R FILLER_1_908 ();
 FILLER_ASAP7_75t_R FILLER_1_916 ();
 FILLER_ASAP7_75t_R FILLER_1_923 ();
 DECAPx1_ASAP7_75t_R FILLER_1_927 ();
 FILLER_ASAP7_75t_R FILLER_1_938 ();
 FILLER_ASAP7_75t_R FILLER_1_946 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_1_968 ();
 FILLER_ASAP7_75t_R FILLER_1_991 ();
 FILLER_ASAP7_75t_R FILLER_1_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_1_1021 ();
 FILLER_ASAP7_75t_R FILLER_1_1045 ();
 DECAPx1_ASAP7_75t_R FILLER_1_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1056 ();
 FILLER_ASAP7_75t_R FILLER_1_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_1_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_1_1110 ();
 FILLER_ASAP7_75t_R FILLER_1_1116 ();
 DECAPx2_ASAP7_75t_R FILLER_1_1138 ();
 FILLER_ASAP7_75t_R FILLER_1_1151 ();
 FILLER_ASAP7_75t_R FILLER_1_1158 ();
 FILLER_ASAP7_75t_R FILLER_1_1180 ();
 FILLER_ASAP7_75t_R FILLER_1_1187 ();
 FILLER_ASAP7_75t_R FILLER_1_1196 ();
 FILLER_ASAP7_75t_R FILLER_1_1204 ();
 FILLER_ASAP7_75t_R FILLER_1_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_1_1343 ();
 DECAPx4_ASAP7_75t_R FILLER_1_1365 ();
 FILLER_ASAP7_75t_R FILLER_1_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_2_24 ();
 DECAPx10_ASAP7_75t_R FILLER_2_46 ();
 DECAPx10_ASAP7_75t_R FILLER_2_68 ();
 DECAPx10_ASAP7_75t_R FILLER_2_90 ();
 DECAPx10_ASAP7_75t_R FILLER_2_112 ();
 DECAPx10_ASAP7_75t_R FILLER_2_134 ();
 DECAPx10_ASAP7_75t_R FILLER_2_156 ();
 DECAPx10_ASAP7_75t_R FILLER_2_178 ();
 DECAPx10_ASAP7_75t_R FILLER_2_200 ();
 DECAPx10_ASAP7_75t_R FILLER_2_222 ();
 DECAPx10_ASAP7_75t_R FILLER_2_244 ();
 DECAPx10_ASAP7_75t_R FILLER_2_266 ();
 DECAPx10_ASAP7_75t_R FILLER_2_288 ();
 DECAPx10_ASAP7_75t_R FILLER_2_310 ();
 DECAPx10_ASAP7_75t_R FILLER_2_332 ();
 DECAPx10_ASAP7_75t_R FILLER_2_354 ();
 DECAPx10_ASAP7_75t_R FILLER_2_376 ();
 DECAPx10_ASAP7_75t_R FILLER_2_398 ();
 DECAPx10_ASAP7_75t_R FILLER_2_420 ();
 DECAPx6_ASAP7_75t_R FILLER_2_442 ();
 DECAPx2_ASAP7_75t_R FILLER_2_456 ();
 FILLER_ASAP7_75t_R FILLER_2_464 ();
 DECAPx2_ASAP7_75t_R FILLER_2_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_478 ();
 FILLER_ASAP7_75t_R FILLER_2_484 ();
 FILLER_ASAP7_75t_R FILLER_2_493 ();
 FILLER_ASAP7_75t_R FILLER_2_501 ();
 FILLER_ASAP7_75t_R FILLER_2_509 ();
 DECAPx2_ASAP7_75t_R FILLER_2_518 ();
 FILLER_ASAP7_75t_R FILLER_2_530 ();
 DECAPx1_ASAP7_75t_R FILLER_2_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_543 ();
 DECAPx1_ASAP7_75t_R FILLER_2_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_568 ();
 FILLER_ASAP7_75t_R FILLER_2_589 ();
 FILLER_ASAP7_75t_R FILLER_2_611 ();
 DECAPx1_ASAP7_75t_R FILLER_2_619 ();
 DECAPx1_ASAP7_75t_R FILLER_2_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_633 ();
 DECAPx2_ASAP7_75t_R FILLER_2_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_660 ();
 FILLER_ASAP7_75t_R FILLER_2_667 ();
 FILLER_ASAP7_75t_R FILLER_2_689 ();
 FILLER_ASAP7_75t_R FILLER_2_697 ();
 DECAPx2_ASAP7_75t_R FILLER_2_705 ();
 FILLER_ASAP7_75t_R FILLER_2_711 ();
 FILLER_ASAP7_75t_R FILLER_2_733 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_2_738 ();
 FILLER_ASAP7_75t_R FILLER_2_747 ();
 DECAPx4_ASAP7_75t_R FILLER_2_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_764 ();
 DECAPx2_ASAP7_75t_R FILLER_2_785 ();
 FILLER_ASAP7_75t_R FILLER_2_796 ();
 FILLER_ASAP7_75t_R FILLER_2_803 ();
 FILLER_ASAP7_75t_R FILLER_2_810 ();
 DECAPx2_ASAP7_75t_R FILLER_2_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_823 ();
 FILLER_ASAP7_75t_R FILLER_2_831 ();
 FILLER_ASAP7_75t_R FILLER_2_838 ();
 FILLER_ASAP7_75t_R FILLER_2_845 ();
 FILLER_ASAP7_75t_R FILLER_2_853 ();
 FILLER_ASAP7_75t_R FILLER_2_861 ();
 DECAPx1_ASAP7_75t_R FILLER_2_868 ();
 DECAPx1_ASAP7_75t_R FILLER_2_879 ();
 FILLER_ASAP7_75t_R FILLER_2_888 ();
 FILLER_ASAP7_75t_R FILLER_2_896 ();
 FILLER_ASAP7_75t_R FILLER_2_904 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_2_913 ();
 FILLER_ASAP7_75t_R FILLER_2_936 ();
 FILLER_ASAP7_75t_R FILLER_2_944 ();
 DECAPx2_ASAP7_75t_R FILLER_2_951 ();
 FILLER_ASAP7_75t_R FILLER_2_964 ();
 DECAPx2_ASAP7_75t_R FILLER_2_971 ();
 FILLER_ASAP7_75t_R FILLER_2_983 ();
 FILLER_ASAP7_75t_R FILLER_2_990 ();
 DECAPx2_ASAP7_75t_R FILLER_2_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1003 ();
 FILLER_ASAP7_75t_R FILLER_2_1010 ();
 FILLER_ASAP7_75t_R FILLER_2_1017 ();
 FILLER_ASAP7_75t_R FILLER_2_1024 ();
 DECAPx1_ASAP7_75t_R FILLER_2_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_1035 ();
 DECAPx2_ASAP7_75t_R FILLER_2_1042 ();
 FILLER_ASAP7_75t_R FILLER_2_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_2_1063 ();
 FILLER_ASAP7_75t_R FILLER_2_1075 ();
 FILLER_ASAP7_75t_R FILLER_2_1083 ();
 FILLER_ASAP7_75t_R FILLER_2_1090 ();
 FILLER_ASAP7_75t_R FILLER_2_1097 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_2_1104 ();
 FILLER_ASAP7_75t_R FILLER_2_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_2_1121 ();
 FILLER_ASAP7_75t_R FILLER_2_1127 ();
 DECAPx1_ASAP7_75t_R FILLER_2_1135 ();
 FILLER_ASAP7_75t_R FILLER_2_1159 ();
 DECAPx1_ASAP7_75t_R FILLER_2_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_2_1177 ();
 FILLER_ASAP7_75t_R FILLER_2_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_2_1205 ();
 FILLER_ASAP7_75t_R FILLER_2_1211 ();
 FILLER_ASAP7_75t_R FILLER_2_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_2_1337 ();
 DECAPx6_ASAP7_75t_R FILLER_2_1359 ();
 DECAPx1_ASAP7_75t_R FILLER_2_1373 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_3_68 ();
 DECAPx10_ASAP7_75t_R FILLER_3_90 ();
 DECAPx10_ASAP7_75t_R FILLER_3_112 ();
 DECAPx10_ASAP7_75t_R FILLER_3_134 ();
 DECAPx10_ASAP7_75t_R FILLER_3_156 ();
 DECAPx10_ASAP7_75t_R FILLER_3_178 ();
 DECAPx10_ASAP7_75t_R FILLER_3_200 ();
 DECAPx10_ASAP7_75t_R FILLER_3_222 ();
 DECAPx10_ASAP7_75t_R FILLER_3_244 ();
 DECAPx10_ASAP7_75t_R FILLER_3_266 ();
 DECAPx10_ASAP7_75t_R FILLER_3_288 ();
 DECAPx10_ASAP7_75t_R FILLER_3_310 ();
 DECAPx10_ASAP7_75t_R FILLER_3_332 ();
 DECAPx10_ASAP7_75t_R FILLER_3_354 ();
 DECAPx10_ASAP7_75t_R FILLER_3_376 ();
 DECAPx10_ASAP7_75t_R FILLER_3_398 ();
 DECAPx6_ASAP7_75t_R FILLER_3_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_434 ();
 FILLER_ASAP7_75t_R FILLER_3_442 ();
 DECAPx4_ASAP7_75t_R FILLER_3_450 ();
 DECAPx2_ASAP7_75t_R FILLER_3_466 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_3_472 ();
 FILLER_ASAP7_75t_R FILLER_3_480 ();
 FILLER_ASAP7_75t_R FILLER_3_487 ();
 FILLER_ASAP7_75t_R FILLER_3_494 ();
 DECAPx1_ASAP7_75t_R FILLER_3_501 ();
 FILLER_ASAP7_75t_R FILLER_3_510 ();
 DECAPx6_ASAP7_75t_R FILLER_3_518 ();
 FILLER_ASAP7_75t_R FILLER_3_532 ();
 FILLER_ASAP7_75t_R FILLER_3_540 ();
 DECAPx1_ASAP7_75t_R FILLER_3_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_552 ();
 FILLER_ASAP7_75t_R FILLER_3_560 ();
 DECAPx2_ASAP7_75t_R FILLER_3_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_574 ();
 FILLER_ASAP7_75t_R FILLER_3_582 ();
 FILLER_ASAP7_75t_R FILLER_3_590 ();
 FILLER_ASAP7_75t_R FILLER_3_597 ();
 FILLER_ASAP7_75t_R FILLER_3_606 ();
 DECAPx2_ASAP7_75t_R FILLER_3_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_620 ();
 FILLER_ASAP7_75t_R FILLER_3_628 ();
 DECAPx2_ASAP7_75t_R FILLER_3_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_642 ();
 DECAPx10_ASAP7_75t_R FILLER_3_649 ();
 FILLER_ASAP7_75t_R FILLER_3_671 ();
 FILLER_ASAP7_75t_R FILLER_3_678 ();
 DECAPx2_ASAP7_75t_R FILLER_3_686 ();
 FILLER_ASAP7_75t_R FILLER_3_697 ();
 FILLER_ASAP7_75t_R FILLER_3_706 ();
 DECAPx2_ASAP7_75t_R FILLER_3_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_720 ();
 FILLER_ASAP7_75t_R FILLER_3_727 ();
 DECAPx2_ASAP7_75t_R FILLER_3_734 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_3_740 ();
 DECAPx4_ASAP7_75t_R FILLER_3_750 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_3_760 ();
 FILLER_ASAP7_75t_R FILLER_3_769 ();
 DECAPx10_ASAP7_75t_R FILLER_3_777 ();
 DECAPx1_ASAP7_75t_R FILLER_3_799 ();
 DECAPx2_ASAP7_75t_R FILLER_3_809 ();
 FILLER_ASAP7_75t_R FILLER_3_835 ();
 FILLER_ASAP7_75t_R FILLER_3_843 ();
 FILLER_ASAP7_75t_R FILLER_3_850 ();
 DECAPx6_ASAP7_75t_R FILLER_3_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_871 ();
 DECAPx10_ASAP7_75t_R FILLER_3_875 ();
 FILLER_ASAP7_75t_R FILLER_3_897 ();
 DECAPx2_ASAP7_75t_R FILLER_3_919 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_3_927 ();
 FILLER_ASAP7_75t_R FILLER_3_952 ();
 FILLER_ASAP7_75t_R FILLER_3_959 ();
 FILLER_ASAP7_75t_R FILLER_3_966 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_3_971 ();
 DECAPx2_ASAP7_75t_R FILLER_3_980 ();
 FILLER_ASAP7_75t_R FILLER_3_986 ();
 FILLER_ASAP7_75t_R FILLER_3_993 ();
 FILLER_ASAP7_75t_R FILLER_3_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_3_1007 ();
 DECAPx6_ASAP7_75t_R FILLER_3_1020 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_3_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_3_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_3_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1079 ();
 FILLER_ASAP7_75t_R FILLER_3_1087 ();
 DECAPx6_ASAP7_75t_R FILLER_3_1095 ();
 DECAPx6_ASAP7_75t_R FILLER_3_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1128 ();
 DECAPx6_ASAP7_75t_R FILLER_3_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_1149 ();
 FILLER_ASAP7_75t_R FILLER_3_1156 ();
 DECAPx2_ASAP7_75t_R FILLER_3_1164 ();
 FILLER_ASAP7_75t_R FILLER_3_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_3_1178 ();
 FILLER_ASAP7_75t_R FILLER_3_1187 ();
 FILLER_ASAP7_75t_R FILLER_3_1195 ();
 FILLER_ASAP7_75t_R FILLER_3_1203 ();
 FILLER_ASAP7_75t_R FILLER_3_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_3_1349 ();
 DECAPx2_ASAP7_75t_R FILLER_3_1371 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_4_68 ();
 DECAPx10_ASAP7_75t_R FILLER_4_90 ();
 DECAPx10_ASAP7_75t_R FILLER_4_112 ();
 DECAPx10_ASAP7_75t_R FILLER_4_134 ();
 DECAPx10_ASAP7_75t_R FILLER_4_156 ();
 DECAPx10_ASAP7_75t_R FILLER_4_178 ();
 DECAPx10_ASAP7_75t_R FILLER_4_200 ();
 DECAPx10_ASAP7_75t_R FILLER_4_222 ();
 DECAPx10_ASAP7_75t_R FILLER_4_244 ();
 DECAPx10_ASAP7_75t_R FILLER_4_266 ();
 DECAPx10_ASAP7_75t_R FILLER_4_288 ();
 DECAPx10_ASAP7_75t_R FILLER_4_310 ();
 DECAPx10_ASAP7_75t_R FILLER_4_332 ();
 DECAPx10_ASAP7_75t_R FILLER_4_354 ();
 DECAPx10_ASAP7_75t_R FILLER_4_376 ();
 DECAPx10_ASAP7_75t_R FILLER_4_398 ();
 DECAPx2_ASAP7_75t_R FILLER_4_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_426 ();
 DECAPx6_ASAP7_75t_R FILLER_4_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_461 ();
 FILLER_ASAP7_75t_R FILLER_4_464 ();
 DECAPx4_ASAP7_75t_R FILLER_4_472 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_4_482 ();
 FILLER_ASAP7_75t_R FILLER_4_490 ();
 DECAPx2_ASAP7_75t_R FILLER_4_500 ();
 FILLER_ASAP7_75t_R FILLER_4_511 ();
 DECAPx6_ASAP7_75t_R FILLER_4_519 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_4_539 ();
 FILLER_ASAP7_75t_R FILLER_4_547 ();
 FILLER_ASAP7_75t_R FILLER_4_554 ();
 FILLER_ASAP7_75t_R FILLER_4_561 ();
 FILLER_ASAP7_75t_R FILLER_4_568 ();
 DECAPx4_ASAP7_75t_R FILLER_4_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_585 ();
 DECAPx2_ASAP7_75t_R FILLER_4_591 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_4_597 ();
 DECAPx2_ASAP7_75t_R FILLER_4_605 ();
 FILLER_ASAP7_75t_R FILLER_4_611 ();
 DECAPx10_ASAP7_75t_R FILLER_4_618 ();
 FILLER_ASAP7_75t_R FILLER_4_640 ();
 FILLER_ASAP7_75t_R FILLER_4_649 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_4_657 ();
 FILLER_ASAP7_75t_R FILLER_4_667 ();
 DECAPx1_ASAP7_75t_R FILLER_4_675 ();
 FILLER_ASAP7_75t_R FILLER_4_686 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_4_694 ();
 FILLER_ASAP7_75t_R FILLER_4_702 ();
 DECAPx4_ASAP7_75t_R FILLER_4_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_719 ();
 DECAPx10_ASAP7_75t_R FILLER_4_726 ();
 DECAPx6_ASAP7_75t_R FILLER_4_748 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_4_762 ();
 DECAPx4_ASAP7_75t_R FILLER_4_773 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_4_783 ();
 FILLER_ASAP7_75t_R FILLER_4_806 ();
 FILLER_ASAP7_75t_R FILLER_4_815 ();
 DECAPx1_ASAP7_75t_R FILLER_4_822 ();
 FILLER_ASAP7_75t_R FILLER_4_832 ();
 DECAPx2_ASAP7_75t_R FILLER_4_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_846 ();
 FILLER_ASAP7_75t_R FILLER_4_854 ();
 DECAPx10_ASAP7_75t_R FILLER_4_862 ();
 DECAPx10_ASAP7_75t_R FILLER_4_884 ();
 DECAPx1_ASAP7_75t_R FILLER_4_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_910 ();
 FILLER_ASAP7_75t_R FILLER_4_919 ();
 DECAPx2_ASAP7_75t_R FILLER_4_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_933 ();
 FILLER_ASAP7_75t_R FILLER_4_954 ();
 FILLER_ASAP7_75t_R FILLER_4_962 ();
 FILLER_ASAP7_75t_R FILLER_4_969 ();
 DECAPx4_ASAP7_75t_R FILLER_4_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_986 ();
 DECAPx4_ASAP7_75t_R FILLER_4_994 ();
 FILLER_ASAP7_75t_R FILLER_4_1004 ();
 FILLER_ASAP7_75t_R FILLER_4_1012 ();
 DECAPx6_ASAP7_75t_R FILLER_4_1034 ();
 DECAPx1_ASAP7_75t_R FILLER_4_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_1052 ();
 FILLER_ASAP7_75t_R FILLER_4_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_4_1067 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_4_1073 ();
 FILLER_ASAP7_75t_R FILLER_4_1096 ();
 DECAPx1_ASAP7_75t_R FILLER_4_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_4_1181 ();
 FILLER_ASAP7_75t_R FILLER_4_1187 ();
 DECAPx1_ASAP7_75t_R FILLER_4_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_4_1205 ();
 FILLER_ASAP7_75t_R FILLER_4_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_4_1351 ();
 DECAPx1_ASAP7_75t_R FILLER_4_1373 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 DECAPx10_ASAP7_75t_R FILLER_5_24 ();
 DECAPx10_ASAP7_75t_R FILLER_5_46 ();
 DECAPx10_ASAP7_75t_R FILLER_5_68 ();
 DECAPx10_ASAP7_75t_R FILLER_5_90 ();
 DECAPx10_ASAP7_75t_R FILLER_5_112 ();
 DECAPx10_ASAP7_75t_R FILLER_5_134 ();
 DECAPx10_ASAP7_75t_R FILLER_5_156 ();
 DECAPx10_ASAP7_75t_R FILLER_5_178 ();
 DECAPx10_ASAP7_75t_R FILLER_5_200 ();
 DECAPx10_ASAP7_75t_R FILLER_5_222 ();
 DECAPx10_ASAP7_75t_R FILLER_5_244 ();
 DECAPx10_ASAP7_75t_R FILLER_5_266 ();
 DECAPx10_ASAP7_75t_R FILLER_5_288 ();
 DECAPx10_ASAP7_75t_R FILLER_5_310 ();
 DECAPx10_ASAP7_75t_R FILLER_5_332 ();
 DECAPx10_ASAP7_75t_R FILLER_5_354 ();
 DECAPx10_ASAP7_75t_R FILLER_5_376 ();
 DECAPx10_ASAP7_75t_R FILLER_5_398 ();
 DECAPx6_ASAP7_75t_R FILLER_5_420 ();
 DECAPx2_ASAP7_75t_R FILLER_5_434 ();
 DECAPx6_ASAP7_75t_R FILLER_5_446 ();
 DECAPx2_ASAP7_75t_R FILLER_5_480 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_5_486 ();
 DECAPx1_ASAP7_75t_R FILLER_5_509 ();
 DECAPx4_ASAP7_75t_R FILLER_5_521 ();
 FILLER_ASAP7_75t_R FILLER_5_531 ();
 DECAPx6_ASAP7_75t_R FILLER_5_541 ();
 FILLER_ASAP7_75t_R FILLER_5_563 ();
 DECAPx1_ASAP7_75t_R FILLER_5_571 ();
 FILLER_ASAP7_75t_R FILLER_5_583 ();
 DECAPx2_ASAP7_75t_R FILLER_5_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_597 ();
 FILLER_ASAP7_75t_R FILLER_5_606 ();
 DECAPx1_ASAP7_75t_R FILLER_5_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_618 ();
 FILLER_ASAP7_75t_R FILLER_5_627 ();
 DECAPx10_ASAP7_75t_R FILLER_5_635 ();
 DECAPx10_ASAP7_75t_R FILLER_5_657 ();
 DECAPx4_ASAP7_75t_R FILLER_5_685 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_5_695 ();
 FILLER_ASAP7_75t_R FILLER_5_706 ();
 DECAPx2_ASAP7_75t_R FILLER_5_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_720 ();
 FILLER_ASAP7_75t_R FILLER_5_728 ();
 DECAPx2_ASAP7_75t_R FILLER_5_736 ();
 FILLER_ASAP7_75t_R FILLER_5_750 ();
 DECAPx1_ASAP7_75t_R FILLER_5_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_762 ();
 DECAPx10_ASAP7_75t_R FILLER_5_783 ();
 FILLER_ASAP7_75t_R FILLER_5_811 ();
 DECAPx6_ASAP7_75t_R FILLER_5_819 ();
 DECAPx1_ASAP7_75t_R FILLER_5_833 ();
 FILLER_ASAP7_75t_R FILLER_5_857 ();
 DECAPx1_ASAP7_75t_R FILLER_5_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_871 ();
 FILLER_ASAP7_75t_R FILLER_5_880 ();
 DECAPx10_ASAP7_75t_R FILLER_5_888 ();
 DECAPx6_ASAP7_75t_R FILLER_5_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_924 ();
 FILLER_ASAP7_75t_R FILLER_5_927 ();
 DECAPx2_ASAP7_75t_R FILLER_5_951 ();
 FILLER_ASAP7_75t_R FILLER_5_965 ();
 FILLER_ASAP7_75t_R FILLER_5_973 ();
 FILLER_ASAP7_75t_R FILLER_5_995 ();
 DECAPx1_ASAP7_75t_R FILLER_5_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1007 ();
 FILLER_ASAP7_75t_R FILLER_5_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1022 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1044 ();
 DECAPx6_ASAP7_75t_R FILLER_5_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_5_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1086 ();
 DECAPx4_ASAP7_75t_R FILLER_5_1093 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_5_1103 ();
 FILLER_ASAP7_75t_R FILLER_5_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_5_1156 ();
 DECAPx1_ASAP7_75t_R FILLER_5_1170 ();
 DECAPx4_ASAP7_75t_R FILLER_5_1186 ();
 FILLER_ASAP7_75t_R FILLER_5_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_5_1334 ();
 DECAPx6_ASAP7_75t_R FILLER_5_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_5_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_6_24 ();
 DECAPx10_ASAP7_75t_R FILLER_6_46 ();
 DECAPx10_ASAP7_75t_R FILLER_6_68 ();
 DECAPx10_ASAP7_75t_R FILLER_6_90 ();
 DECAPx10_ASAP7_75t_R FILLER_6_112 ();
 DECAPx10_ASAP7_75t_R FILLER_6_134 ();
 DECAPx10_ASAP7_75t_R FILLER_6_156 ();
 DECAPx10_ASAP7_75t_R FILLER_6_178 ();
 DECAPx10_ASAP7_75t_R FILLER_6_200 ();
 DECAPx10_ASAP7_75t_R FILLER_6_222 ();
 DECAPx10_ASAP7_75t_R FILLER_6_244 ();
 DECAPx10_ASAP7_75t_R FILLER_6_266 ();
 DECAPx10_ASAP7_75t_R FILLER_6_288 ();
 DECAPx10_ASAP7_75t_R FILLER_6_310 ();
 DECAPx10_ASAP7_75t_R FILLER_6_332 ();
 DECAPx10_ASAP7_75t_R FILLER_6_354 ();
 DECAPx10_ASAP7_75t_R FILLER_6_376 ();
 DECAPx10_ASAP7_75t_R FILLER_6_398 ();
 DECAPx6_ASAP7_75t_R FILLER_6_420 ();
 DECAPx2_ASAP7_75t_R FILLER_6_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_440 ();
 DECAPx6_ASAP7_75t_R FILLER_6_448 ();
 FILLER_ASAP7_75t_R FILLER_6_464 ();
 FILLER_ASAP7_75t_R FILLER_6_472 ();
 DECAPx4_ASAP7_75t_R FILLER_6_477 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_6_487 ();
 DECAPx2_ASAP7_75t_R FILLER_6_496 ();
 FILLER_ASAP7_75t_R FILLER_6_502 ();
 FILLER_ASAP7_75t_R FILLER_6_524 ();
 FILLER_ASAP7_75t_R FILLER_6_546 ();
 FILLER_ASAP7_75t_R FILLER_6_568 ();
 FILLER_ASAP7_75t_R FILLER_6_590 ();
 FILLER_ASAP7_75t_R FILLER_6_612 ();
 DECAPx1_ASAP7_75t_R FILLER_6_634 ();
 FILLER_ASAP7_75t_R FILLER_6_646 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_6_654 ();
 FILLER_ASAP7_75t_R FILLER_6_665 ();
 DECAPx1_ASAP7_75t_R FILLER_6_673 ();
 DECAPx2_ASAP7_75t_R FILLER_6_685 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_6_691 ();
 DECAPx2_ASAP7_75t_R FILLER_6_714 ();
 FILLER_ASAP7_75t_R FILLER_6_720 ();
 DECAPx2_ASAP7_75t_R FILLER_6_730 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_6_736 ();
 DECAPx1_ASAP7_75t_R FILLER_6_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_763 ();
 DECAPx10_ASAP7_75t_R FILLER_6_770 ();
 DECAPx10_ASAP7_75t_R FILLER_6_792 ();
 DECAPx10_ASAP7_75t_R FILLER_6_814 ();
 DECAPx6_ASAP7_75t_R FILLER_6_836 ();
 DECAPx4_ASAP7_75t_R FILLER_6_856 ();
 DECAPx6_ASAP7_75t_R FILLER_6_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_900 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_6_910 ();
 DECAPx4_ASAP7_75t_R FILLER_6_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_935 ();
 DECAPx4_ASAP7_75t_R FILLER_6_943 ();
 FILLER_ASAP7_75t_R FILLER_6_953 ();
 DECAPx10_ASAP7_75t_R FILLER_6_961 ();
 DECAPx2_ASAP7_75t_R FILLER_6_983 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_6_989 ();
 FILLER_ASAP7_75t_R FILLER_6_998 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1028 ();
 DECAPx2_ASAP7_75t_R FILLER_6_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_6_1063 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_6_1069 ();
 FILLER_ASAP7_75t_R FILLER_6_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1087 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_6_1109 ();
 DECAPx1_ASAP7_75t_R FILLER_6_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1122 ();
 DECAPx2_ASAP7_75t_R FILLER_6_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_6_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_1161 ();
 FILLER_ASAP7_75t_R FILLER_6_1182 ();
 FILLER_ASAP7_75t_R FILLER_6_1191 ();
 DECAPx4_ASAP7_75t_R FILLER_6_1199 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_6_1209 ();
 DECAPx4_ASAP7_75t_R FILLER_6_1218 ();
 FILLER_ASAP7_75t_R FILLER_6_1228 ();
 FILLER_ASAP7_75t_R FILLER_6_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_6_1355 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 DECAPx10_ASAP7_75t_R FILLER_7_24 ();
 DECAPx10_ASAP7_75t_R FILLER_7_46 ();
 DECAPx10_ASAP7_75t_R FILLER_7_68 ();
 DECAPx10_ASAP7_75t_R FILLER_7_90 ();
 DECAPx10_ASAP7_75t_R FILLER_7_112 ();
 DECAPx10_ASAP7_75t_R FILLER_7_134 ();
 DECAPx10_ASAP7_75t_R FILLER_7_156 ();
 DECAPx10_ASAP7_75t_R FILLER_7_178 ();
 DECAPx10_ASAP7_75t_R FILLER_7_200 ();
 DECAPx10_ASAP7_75t_R FILLER_7_222 ();
 DECAPx10_ASAP7_75t_R FILLER_7_244 ();
 DECAPx10_ASAP7_75t_R FILLER_7_266 ();
 DECAPx10_ASAP7_75t_R FILLER_7_288 ();
 DECAPx10_ASAP7_75t_R FILLER_7_310 ();
 DECAPx10_ASAP7_75t_R FILLER_7_332 ();
 DECAPx10_ASAP7_75t_R FILLER_7_354 ();
 DECAPx10_ASAP7_75t_R FILLER_7_376 ();
 DECAPx10_ASAP7_75t_R FILLER_7_398 ();
 DECAPx6_ASAP7_75t_R FILLER_7_420 ();
 DECAPx1_ASAP7_75t_R FILLER_7_434 ();
 FILLER_ASAP7_75t_R FILLER_7_444 ();
 DECAPx6_ASAP7_75t_R FILLER_7_454 ();
 FILLER_ASAP7_75t_R FILLER_7_468 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_7_473 ();
 DECAPx2_ASAP7_75t_R FILLER_7_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_502 ();
 DECAPx10_ASAP7_75t_R FILLER_7_506 ();
 DECAPx4_ASAP7_75t_R FILLER_7_528 ();
 FILLER_ASAP7_75t_R FILLER_7_538 ();
 DECAPx10_ASAP7_75t_R FILLER_7_543 ();
 DECAPx4_ASAP7_75t_R FILLER_7_565 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_7_575 ();
 DECAPx6_ASAP7_75t_R FILLER_7_581 ();
 DECAPx2_ASAP7_75t_R FILLER_7_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_601 ();
 DECAPx10_ASAP7_75t_R FILLER_7_605 ();
 FILLER_ASAP7_75t_R FILLER_7_627 ();
 FILLER_ASAP7_75t_R FILLER_7_649 ();
 FILLER_ASAP7_75t_R FILLER_7_671 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_7_693 ();
 DECAPx6_ASAP7_75t_R FILLER_7_699 ();
 DECAPx2_ASAP7_75t_R FILLER_7_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_719 ();
 DECAPx10_ASAP7_75t_R FILLER_7_740 ();
 FILLER_ASAP7_75t_R FILLER_7_765 ();
 DECAPx6_ASAP7_75t_R FILLER_7_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_784 ();
 DECAPx10_ASAP7_75t_R FILLER_7_792 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_7_814 ();
 FILLER_ASAP7_75t_R FILLER_7_825 ();
 DECAPx10_ASAP7_75t_R FILLER_7_833 ();
 DECAPx6_ASAP7_75t_R FILLER_7_855 ();
 FILLER_ASAP7_75t_R FILLER_7_869 ();
 FILLER_ASAP7_75t_R FILLER_7_878 ();
 DECAPx1_ASAP7_75t_R FILLER_7_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_890 ();
 FILLER_ASAP7_75t_R FILLER_7_911 ();
 DECAPx2_ASAP7_75t_R FILLER_7_919 ();
 FILLER_ASAP7_75t_R FILLER_7_927 ();
 DECAPx6_ASAP7_75t_R FILLER_7_936 ();
 DECAPx1_ASAP7_75t_R FILLER_7_957 ();
 DECAPx4_ASAP7_75t_R FILLER_7_969 ();
 DECAPx10_ASAP7_75t_R FILLER_7_985 ();
 DECAPx4_ASAP7_75t_R FILLER_7_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_7_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_1034 ();
 FILLER_ASAP7_75t_R FILLER_7_1044 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_7_1054 ();
 FILLER_ASAP7_75t_R FILLER_7_1069 ();
 DECAPx2_ASAP7_75t_R FILLER_7_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_1097 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_7_1104 ();
 DECAPx6_ASAP7_75t_R FILLER_7_1113 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_7_1134 ();
 FILLER_ASAP7_75t_R FILLER_7_1149 ();
 FILLER_ASAP7_75t_R FILLER_7_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_7_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_7_1182 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_7_1188 ();
 DECAPx4_ASAP7_75t_R FILLER_7_1200 ();
 FILLER_ASAP7_75t_R FILLER_7_1216 ();
 FILLER_ASAP7_75t_R FILLER_7_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_7_1340 ();
 DECAPx6_ASAP7_75t_R FILLER_7_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_8_2 ();
 DECAPx10_ASAP7_75t_R FILLER_8_24 ();
 DECAPx10_ASAP7_75t_R FILLER_8_46 ();
 DECAPx10_ASAP7_75t_R FILLER_8_68 ();
 DECAPx10_ASAP7_75t_R FILLER_8_90 ();
 DECAPx10_ASAP7_75t_R FILLER_8_112 ();
 DECAPx10_ASAP7_75t_R FILLER_8_134 ();
 DECAPx10_ASAP7_75t_R FILLER_8_156 ();
 DECAPx10_ASAP7_75t_R FILLER_8_178 ();
 DECAPx10_ASAP7_75t_R FILLER_8_200 ();
 DECAPx10_ASAP7_75t_R FILLER_8_222 ();
 DECAPx10_ASAP7_75t_R FILLER_8_244 ();
 DECAPx10_ASAP7_75t_R FILLER_8_266 ();
 DECAPx10_ASAP7_75t_R FILLER_8_288 ();
 DECAPx10_ASAP7_75t_R FILLER_8_310 ();
 DECAPx10_ASAP7_75t_R FILLER_8_332 ();
 DECAPx10_ASAP7_75t_R FILLER_8_354 ();
 DECAPx10_ASAP7_75t_R FILLER_8_376 ();
 DECAPx10_ASAP7_75t_R FILLER_8_398 ();
 DECAPx6_ASAP7_75t_R FILLER_8_420 ();
 DECAPx1_ASAP7_75t_R FILLER_8_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_438 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_459 ();
 DECAPx1_ASAP7_75t_R FILLER_8_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_468 ();
 DECAPx10_ASAP7_75t_R FILLER_8_481 ();
 DECAPx6_ASAP7_75t_R FILLER_8_503 ();
 DECAPx1_ASAP7_75t_R FILLER_8_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_521 ();
 DECAPx6_ASAP7_75t_R FILLER_8_525 ();
 DECAPx10_ASAP7_75t_R FILLER_8_551 ();
 FILLER_ASAP7_75t_R FILLER_8_573 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_587 ();
 DECAPx10_ASAP7_75t_R FILLER_8_593 ();
 DECAPx10_ASAP7_75t_R FILLER_8_615 ();
 DECAPx10_ASAP7_75t_R FILLER_8_637 ();
 DECAPx2_ASAP7_75t_R FILLER_8_659 ();
 DECAPx10_ASAP7_75t_R FILLER_8_668 ();
 DECAPx10_ASAP7_75t_R FILLER_8_690 ();
 DECAPx10_ASAP7_75t_R FILLER_8_712 ();
 DECAPx4_ASAP7_75t_R FILLER_8_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_744 ();
 FILLER_ASAP7_75t_R FILLER_8_765 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_773 ();
 FILLER_ASAP7_75t_R FILLER_8_782 ();
 FILLER_ASAP7_75t_R FILLER_8_804 ();
 FILLER_ASAP7_75t_R FILLER_8_826 ();
 FILLER_ASAP7_75t_R FILLER_8_837 ();
 DECAPx2_ASAP7_75t_R FILLER_8_842 ();
 FILLER_ASAP7_75t_R FILLER_8_848 ();
 DECAPx10_ASAP7_75t_R FILLER_8_858 ();
 DECAPx4_ASAP7_75t_R FILLER_8_880 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_890 ();
 FILLER_ASAP7_75t_R FILLER_8_901 ();
 FILLER_ASAP7_75t_R FILLER_8_911 ();
 DECAPx1_ASAP7_75t_R FILLER_8_920 ();
 FILLER_ASAP7_75t_R FILLER_8_944 ();
 FILLER_ASAP7_75t_R FILLER_8_966 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_974 ();
 DECAPx1_ASAP7_75t_R FILLER_8_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1001 ();
 FILLER_ASAP7_75t_R FILLER_8_1022 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_8_1054 ();
 FILLER_ASAP7_75t_R FILLER_8_1060 ();
 FILLER_ASAP7_75t_R FILLER_8_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_8_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_8_1116 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_8_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1141 ();
 FILLER_ASAP7_75t_R FILLER_8_1149 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_1157 ();
 DECAPx6_ASAP7_75t_R FILLER_8_1169 ();
 FILLER_ASAP7_75t_R FILLER_8_1183 ();
 FILLER_ASAP7_75t_R FILLER_8_1192 ();
 DECAPx4_ASAP7_75t_R FILLER_8_1200 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_8_1222 ();
 FILLER_ASAP7_75t_R FILLER_8_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_8_1348 ();
 DECAPx2_ASAP7_75t_R FILLER_8_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_9_2 ();
 DECAPx10_ASAP7_75t_R FILLER_9_24 ();
 DECAPx10_ASAP7_75t_R FILLER_9_46 ();
 DECAPx10_ASAP7_75t_R FILLER_9_68 ();
 DECAPx10_ASAP7_75t_R FILLER_9_90 ();
 DECAPx10_ASAP7_75t_R FILLER_9_112 ();
 DECAPx10_ASAP7_75t_R FILLER_9_134 ();
 DECAPx10_ASAP7_75t_R FILLER_9_156 ();
 DECAPx10_ASAP7_75t_R FILLER_9_178 ();
 DECAPx10_ASAP7_75t_R FILLER_9_200 ();
 DECAPx10_ASAP7_75t_R FILLER_9_222 ();
 DECAPx10_ASAP7_75t_R FILLER_9_244 ();
 DECAPx10_ASAP7_75t_R FILLER_9_266 ();
 DECAPx10_ASAP7_75t_R FILLER_9_288 ();
 DECAPx10_ASAP7_75t_R FILLER_9_310 ();
 DECAPx10_ASAP7_75t_R FILLER_9_332 ();
 DECAPx10_ASAP7_75t_R FILLER_9_354 ();
 DECAPx10_ASAP7_75t_R FILLER_9_376 ();
 DECAPx10_ASAP7_75t_R FILLER_9_398 ();
 DECAPx10_ASAP7_75t_R FILLER_9_420 ();
 DECAPx2_ASAP7_75t_R FILLER_9_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_448 ();
 DECAPx1_ASAP7_75t_R FILLER_9_459 ();
 FILLER_ASAP7_75t_R FILLER_9_475 ();
 DECAPx2_ASAP7_75t_R FILLER_9_480 ();
 DECAPx2_ASAP7_75t_R FILLER_9_489 ();
 FILLER_ASAP7_75t_R FILLER_9_495 ();
 DECAPx4_ASAP7_75t_R FILLER_9_503 ();
 FILLER_ASAP7_75t_R FILLER_9_516 ();
 FILLER_ASAP7_75t_R FILLER_9_530 ();
 DECAPx1_ASAP7_75t_R FILLER_9_539 ();
 FILLER_ASAP7_75t_R FILLER_9_563 ();
 DECAPx2_ASAP7_75t_R FILLER_9_568 ();
 FILLER_ASAP7_75t_R FILLER_9_574 ();
 FILLER_ASAP7_75t_R FILLER_9_596 ();
 FILLER_ASAP7_75t_R FILLER_9_610 ();
 DECAPx1_ASAP7_75t_R FILLER_9_615 ();
 DECAPx10_ASAP7_75t_R FILLER_9_631 ();
 DECAPx4_ASAP7_75t_R FILLER_9_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_663 ();
 DECAPx2_ASAP7_75t_R FILLER_9_676 ();
 DECAPx1_ASAP7_75t_R FILLER_9_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_689 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_9_702 ();
 FILLER_ASAP7_75t_R FILLER_9_708 ();
 DECAPx4_ASAP7_75t_R FILLER_9_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_727 ();
 DECAPx2_ASAP7_75t_R FILLER_9_734 ();
 DECAPx2_ASAP7_75t_R FILLER_9_752 ();
 FILLER_ASAP7_75t_R FILLER_9_765 ();
 DECAPx2_ASAP7_75t_R FILLER_9_775 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_9_781 ();
 FILLER_ASAP7_75t_R FILLER_9_791 ();
 DECAPx6_ASAP7_75t_R FILLER_9_799 ();
 DECAPx2_ASAP7_75t_R FILLER_9_813 ();
 FILLER_ASAP7_75t_R FILLER_9_827 ();
 DECAPx2_ASAP7_75t_R FILLER_9_832 ();
 FILLER_ASAP7_75t_R FILLER_9_838 ();
 DECAPx4_ASAP7_75t_R FILLER_9_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_870 ();
 DECAPx10_ASAP7_75t_R FILLER_9_878 ();
 DECAPx2_ASAP7_75t_R FILLER_9_900 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_9_906 ();
 DECAPx4_ASAP7_75t_R FILLER_9_915 ();
 FILLER_ASAP7_75t_R FILLER_9_927 ();
 DECAPx10_ASAP7_75t_R FILLER_9_935 ();
 DECAPx4_ASAP7_75t_R FILLER_9_957 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_9_967 ();
 DECAPx1_ASAP7_75t_R FILLER_9_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_986 ();
 FILLER_ASAP7_75t_R FILLER_9_993 ();
 DECAPx6_ASAP7_75t_R FILLER_9_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_9_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1019 ();
 FILLER_ASAP7_75t_R FILLER_9_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_9_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1038 ();
 FILLER_ASAP7_75t_R FILLER_9_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1055 ();
 DECAPx4_ASAP7_75t_R FILLER_9_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1087 ();
 DECAPx4_ASAP7_75t_R FILLER_9_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1162 ();
 DECAPx2_ASAP7_75t_R FILLER_9_1184 ();
 FILLER_ASAP7_75t_R FILLER_9_1190 ();
 FILLER_ASAP7_75t_R FILLER_9_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_9_1340 ();
 DECAPx6_ASAP7_75t_R FILLER_9_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_10_2 ();
 DECAPx10_ASAP7_75t_R FILLER_10_24 ();
 DECAPx10_ASAP7_75t_R FILLER_10_46 ();
 DECAPx10_ASAP7_75t_R FILLER_10_68 ();
 DECAPx10_ASAP7_75t_R FILLER_10_90 ();
 DECAPx10_ASAP7_75t_R FILLER_10_112 ();
 DECAPx10_ASAP7_75t_R FILLER_10_134 ();
 DECAPx10_ASAP7_75t_R FILLER_10_156 ();
 DECAPx10_ASAP7_75t_R FILLER_10_178 ();
 DECAPx10_ASAP7_75t_R FILLER_10_200 ();
 DECAPx10_ASAP7_75t_R FILLER_10_222 ();
 DECAPx10_ASAP7_75t_R FILLER_10_244 ();
 DECAPx10_ASAP7_75t_R FILLER_10_266 ();
 DECAPx10_ASAP7_75t_R FILLER_10_288 ();
 DECAPx10_ASAP7_75t_R FILLER_10_310 ();
 DECAPx10_ASAP7_75t_R FILLER_10_332 ();
 DECAPx10_ASAP7_75t_R FILLER_10_354 ();
 DECAPx10_ASAP7_75t_R FILLER_10_376 ();
 DECAPx10_ASAP7_75t_R FILLER_10_398 ();
 DECAPx10_ASAP7_75t_R FILLER_10_420 ();
 DECAPx6_ASAP7_75t_R FILLER_10_442 ();
 DECAPx2_ASAP7_75t_R FILLER_10_456 ();
 FILLER_ASAP7_75t_R FILLER_10_464 ();
 FILLER_ASAP7_75t_R FILLER_10_486 ();
 DECAPx1_ASAP7_75t_R FILLER_10_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_498 ();
 FILLER_ASAP7_75t_R FILLER_10_507 ();
 DECAPx2_ASAP7_75t_R FILLER_10_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_521 ();
 FILLER_ASAP7_75t_R FILLER_10_542 ();
 DECAPx6_ASAP7_75t_R FILLER_10_550 ();
 DECAPx1_ASAP7_75t_R FILLER_10_564 ();
 DECAPx4_ASAP7_75t_R FILLER_10_574 ();
 DECAPx2_ASAP7_75t_R FILLER_10_590 ();
 FILLER_ASAP7_75t_R FILLER_10_596 ();
 DECAPx1_ASAP7_75t_R FILLER_10_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_622 ();
 FILLER_ASAP7_75t_R FILLER_10_643 ();
 DECAPx4_ASAP7_75t_R FILLER_10_651 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_10_661 ();
 FILLER_ASAP7_75t_R FILLER_10_684 ();
 FILLER_ASAP7_75t_R FILLER_10_706 ();
 FILLER_ASAP7_75t_R FILLER_10_728 ();
 DECAPx2_ASAP7_75t_R FILLER_10_737 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_10_743 ();
 DECAPx6_ASAP7_75t_R FILLER_10_752 ();
 FILLER_ASAP7_75t_R FILLER_10_766 ();
 DECAPx6_ASAP7_75t_R FILLER_10_788 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_10_802 ();
 DECAPx10_ASAP7_75t_R FILLER_10_811 ();
 DECAPx6_ASAP7_75t_R FILLER_10_833 ();
 DECAPx1_ASAP7_75t_R FILLER_10_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_851 ();
 DECAPx4_ASAP7_75t_R FILLER_10_858 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_10_868 ();
 FILLER_ASAP7_75t_R FILLER_10_891 ();
 DECAPx4_ASAP7_75t_R FILLER_10_899 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_10_909 ();
 DECAPx4_ASAP7_75t_R FILLER_10_918 ();
 DECAPx4_ASAP7_75t_R FILLER_10_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_944 ();
 DECAPx10_ASAP7_75t_R FILLER_10_951 ();
 DECAPx10_ASAP7_75t_R FILLER_10_973 ();
 DECAPx6_ASAP7_75t_R FILLER_10_995 ();
 FILLER_ASAP7_75t_R FILLER_10_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_10_1080 ();
 DECAPx6_ASAP7_75t_R FILLER_10_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_10_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1121 ();
 FILLER_ASAP7_75t_R FILLER_10_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_10_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_10_1158 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_10_1164 ();
 FILLER_ASAP7_75t_R FILLER_10_1175 ();
 DECAPx2_ASAP7_75t_R FILLER_10_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_10_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1213 ();
 FILLER_ASAP7_75t_R FILLER_10_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_10_1340 ();
 DECAPx6_ASAP7_75t_R FILLER_10_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_11_2 ();
 DECAPx10_ASAP7_75t_R FILLER_11_24 ();
 DECAPx10_ASAP7_75t_R FILLER_11_46 ();
 DECAPx10_ASAP7_75t_R FILLER_11_68 ();
 DECAPx10_ASAP7_75t_R FILLER_11_90 ();
 DECAPx10_ASAP7_75t_R FILLER_11_112 ();
 DECAPx10_ASAP7_75t_R FILLER_11_134 ();
 DECAPx10_ASAP7_75t_R FILLER_11_156 ();
 DECAPx10_ASAP7_75t_R FILLER_11_178 ();
 DECAPx10_ASAP7_75t_R FILLER_11_200 ();
 DECAPx10_ASAP7_75t_R FILLER_11_222 ();
 DECAPx10_ASAP7_75t_R FILLER_11_244 ();
 DECAPx10_ASAP7_75t_R FILLER_11_266 ();
 DECAPx10_ASAP7_75t_R FILLER_11_288 ();
 DECAPx10_ASAP7_75t_R FILLER_11_310 ();
 DECAPx10_ASAP7_75t_R FILLER_11_332 ();
 DECAPx10_ASAP7_75t_R FILLER_11_354 ();
 DECAPx10_ASAP7_75t_R FILLER_11_376 ();
 DECAPx10_ASAP7_75t_R FILLER_11_398 ();
 DECAPx4_ASAP7_75t_R FILLER_11_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_430 ();
 FILLER_ASAP7_75t_R FILLER_11_438 ();
 FILLER_ASAP7_75t_R FILLER_11_447 ();
 DECAPx10_ASAP7_75t_R FILLER_11_455 ();
 DECAPx1_ASAP7_75t_R FILLER_11_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_481 ();
 FILLER_ASAP7_75t_R FILLER_11_488 ();
 DECAPx2_ASAP7_75t_R FILLER_11_498 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_504 ();
 DECAPx2_ASAP7_75t_R FILLER_11_514 ();
 FILLER_ASAP7_75t_R FILLER_11_520 ();
 DECAPx6_ASAP7_75t_R FILLER_11_528 ();
 DECAPx2_ASAP7_75t_R FILLER_11_550 ();
 FILLER_ASAP7_75t_R FILLER_11_556 ();
 FILLER_ASAP7_75t_R FILLER_11_561 ();
 DECAPx1_ASAP7_75t_R FILLER_11_571 ();
 DECAPx1_ASAP7_75t_R FILLER_11_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_585 ();
 DECAPx6_ASAP7_75t_R FILLER_11_592 ();
 DECAPx1_ASAP7_75t_R FILLER_11_606 ();
 DECAPx2_ASAP7_75t_R FILLER_11_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_622 ();
 FILLER_ASAP7_75t_R FILLER_11_626 ();
 DECAPx4_ASAP7_75t_R FILLER_11_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_641 ();
 FILLER_ASAP7_75t_R FILLER_11_645 ();
 DECAPx2_ASAP7_75t_R FILLER_11_655 ();
 FILLER_ASAP7_75t_R FILLER_11_661 ();
 DECAPx10_ASAP7_75t_R FILLER_11_669 ();
 DECAPx10_ASAP7_75t_R FILLER_11_691 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_713 ();
 DECAPx6_ASAP7_75t_R FILLER_11_722 ();
 DECAPx1_ASAP7_75t_R FILLER_11_736 ();
 FILLER_ASAP7_75t_R FILLER_11_746 ();
 DECAPx10_ASAP7_75t_R FILLER_11_755 ();
 DECAPx10_ASAP7_75t_R FILLER_11_777 ();
 FILLER_ASAP7_75t_R FILLER_11_805 ();
 DECAPx2_ASAP7_75t_R FILLER_11_816 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_822 ();
 FILLER_ASAP7_75t_R FILLER_11_834 ();
 DECAPx1_ASAP7_75t_R FILLER_11_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_848 ();
 DECAPx6_ASAP7_75t_R FILLER_11_858 ();
 FILLER_ASAP7_75t_R FILLER_11_878 ();
 FILLER_ASAP7_75t_R FILLER_11_886 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_891 ();
 DECAPx4_ASAP7_75t_R FILLER_11_900 ();
 DECAPx2_ASAP7_75t_R FILLER_11_916 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_922 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_927 ();
 FILLER_ASAP7_75t_R FILLER_11_942 ();
 DECAPx2_ASAP7_75t_R FILLER_11_964 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_970 ();
 FILLER_ASAP7_75t_R FILLER_11_982 ();
 FILLER_ASAP7_75t_R FILLER_11_992 ();
 DECAPx2_ASAP7_75t_R FILLER_11_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_1006 ();
 FILLER_ASAP7_75t_R FILLER_11_1014 ();
 DECAPx4_ASAP7_75t_R FILLER_11_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_1032 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_1045 ();
 DECAPx4_ASAP7_75t_R FILLER_11_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_1064 ();
 FILLER_ASAP7_75t_R FILLER_11_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_11_1081 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_1087 ();
 DECAPx2_ASAP7_75t_R FILLER_11_1098 ();
 FILLER_ASAP7_75t_R FILLER_11_1104 ();
 DECAPx4_ASAP7_75t_R FILLER_11_1112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_1122 ();
 FILLER_ASAP7_75t_R FILLER_11_1133 ();
 FILLER_ASAP7_75t_R FILLER_11_1141 ();
 FILLER_ASAP7_75t_R FILLER_11_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_11_1185 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_1191 ();
 DECAPx4_ASAP7_75t_R FILLER_11_1202 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_1212 ();
 FILLER_ASAP7_75t_R FILLER_11_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_11_1355 ();
 DECAPx10_ASAP7_75t_R FILLER_12_2 ();
 DECAPx10_ASAP7_75t_R FILLER_12_24 ();
 DECAPx10_ASAP7_75t_R FILLER_12_46 ();
 DECAPx10_ASAP7_75t_R FILLER_12_68 ();
 DECAPx10_ASAP7_75t_R FILLER_12_90 ();
 DECAPx10_ASAP7_75t_R FILLER_12_112 ();
 DECAPx10_ASAP7_75t_R FILLER_12_134 ();
 DECAPx10_ASAP7_75t_R FILLER_12_156 ();
 DECAPx10_ASAP7_75t_R FILLER_12_178 ();
 DECAPx10_ASAP7_75t_R FILLER_12_200 ();
 DECAPx10_ASAP7_75t_R FILLER_12_222 ();
 DECAPx10_ASAP7_75t_R FILLER_12_244 ();
 DECAPx10_ASAP7_75t_R FILLER_12_266 ();
 DECAPx10_ASAP7_75t_R FILLER_12_288 ();
 DECAPx10_ASAP7_75t_R FILLER_12_310 ();
 DECAPx10_ASAP7_75t_R FILLER_12_332 ();
 DECAPx10_ASAP7_75t_R FILLER_12_354 ();
 DECAPx10_ASAP7_75t_R FILLER_12_376 ();
 DECAPx10_ASAP7_75t_R FILLER_12_398 ();
 FILLER_ASAP7_75t_R FILLER_12_420 ();
 DECAPx2_ASAP7_75t_R FILLER_12_442 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_448 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_459 ();
 DECAPx10_ASAP7_75t_R FILLER_12_464 ();
 DECAPx2_ASAP7_75t_R FILLER_12_494 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_500 ();
 FILLER_ASAP7_75t_R FILLER_12_509 ();
 DECAPx6_ASAP7_75t_R FILLER_12_517 ();
 DECAPx1_ASAP7_75t_R FILLER_12_531 ();
 FILLER_ASAP7_75t_R FILLER_12_541 ();
 DECAPx4_ASAP7_75t_R FILLER_12_549 ();
 FILLER_ASAP7_75t_R FILLER_12_559 ();
 DECAPx6_ASAP7_75t_R FILLER_12_567 ();
 DECAPx2_ASAP7_75t_R FILLER_12_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_587 ();
 DECAPx10_ASAP7_75t_R FILLER_12_596 ();
 DECAPx1_ASAP7_75t_R FILLER_12_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_622 ();
 DECAPx6_ASAP7_75t_R FILLER_12_629 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_651 ();
 FILLER_ASAP7_75t_R FILLER_12_660 ();
 FILLER_ASAP7_75t_R FILLER_12_668 ();
 DECAPx10_ASAP7_75t_R FILLER_12_676 ();
 DECAPx1_ASAP7_75t_R FILLER_12_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_702 ();
 DECAPx6_ASAP7_75t_R FILLER_12_709 ();
 FILLER_ASAP7_75t_R FILLER_12_723 ();
 FILLER_ASAP7_75t_R FILLER_12_733 ();
 DECAPx4_ASAP7_75t_R FILLER_12_741 ();
 DECAPx1_ASAP7_75t_R FILLER_12_759 ();
 FILLER_ASAP7_75t_R FILLER_12_769 ();
 DECAPx4_ASAP7_75t_R FILLER_12_777 ();
 FILLER_ASAP7_75t_R FILLER_12_807 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_816 ();
 FILLER_ASAP7_75t_R FILLER_12_839 ();
 FILLER_ASAP7_75t_R FILLER_12_847 ();
 FILLER_ASAP7_75t_R FILLER_12_861 ();
 FILLER_ASAP7_75t_R FILLER_12_869 ();
 DECAPx4_ASAP7_75t_R FILLER_12_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_890 ();
 FILLER_ASAP7_75t_R FILLER_12_897 ();
 FILLER_ASAP7_75t_R FILLER_12_907 ();
 DECAPx2_ASAP7_75t_R FILLER_12_915 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_933 ();
 FILLER_ASAP7_75t_R FILLER_12_948 ();
 FILLER_ASAP7_75t_R FILLER_12_956 ();
 FILLER_ASAP7_75t_R FILLER_12_964 ();
 DECAPx1_ASAP7_75t_R FILLER_12_972 ();
 DECAPx1_ASAP7_75t_R FILLER_12_996 ();
 DECAPx2_ASAP7_75t_R FILLER_12_1006 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_1012 ();
 FILLER_ASAP7_75t_R FILLER_12_1024 ();
 DECAPx1_ASAP7_75t_R FILLER_12_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1038 ();
 FILLER_ASAP7_75t_R FILLER_12_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_12_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1085 ();
 FILLER_ASAP7_75t_R FILLER_12_1106 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_12_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_1144 ();
 FILLER_ASAP7_75t_R FILLER_12_1151 ();
 DECAPx6_ASAP7_75t_R FILLER_12_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_12_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_12_1351 ();
 DECAPx1_ASAP7_75t_R FILLER_12_1373 ();
 DECAPx10_ASAP7_75t_R FILLER_13_2 ();
 DECAPx10_ASAP7_75t_R FILLER_13_24 ();
 DECAPx10_ASAP7_75t_R FILLER_13_46 ();
 DECAPx10_ASAP7_75t_R FILLER_13_68 ();
 DECAPx10_ASAP7_75t_R FILLER_13_90 ();
 DECAPx10_ASAP7_75t_R FILLER_13_112 ();
 DECAPx10_ASAP7_75t_R FILLER_13_134 ();
 DECAPx10_ASAP7_75t_R FILLER_13_156 ();
 DECAPx10_ASAP7_75t_R FILLER_13_178 ();
 DECAPx10_ASAP7_75t_R FILLER_13_200 ();
 DECAPx10_ASAP7_75t_R FILLER_13_222 ();
 DECAPx10_ASAP7_75t_R FILLER_13_244 ();
 DECAPx10_ASAP7_75t_R FILLER_13_266 ();
 DECAPx10_ASAP7_75t_R FILLER_13_288 ();
 DECAPx10_ASAP7_75t_R FILLER_13_310 ();
 DECAPx10_ASAP7_75t_R FILLER_13_332 ();
 DECAPx10_ASAP7_75t_R FILLER_13_354 ();
 DECAPx10_ASAP7_75t_R FILLER_13_376 ();
 DECAPx10_ASAP7_75t_R FILLER_13_398 ();
 DECAPx4_ASAP7_75t_R FILLER_13_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_430 ();
 FILLER_ASAP7_75t_R FILLER_13_437 ();
 DECAPx1_ASAP7_75t_R FILLER_13_445 ();
 FILLER_ASAP7_75t_R FILLER_13_469 ();
 DECAPx10_ASAP7_75t_R FILLER_13_474 ();
 DECAPx2_ASAP7_75t_R FILLER_13_496 ();
 DECAPx4_ASAP7_75t_R FILLER_13_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_524 ();
 DECAPx1_ASAP7_75t_R FILLER_13_533 ();
 FILLER_ASAP7_75t_R FILLER_13_543 ();
 DECAPx1_ASAP7_75t_R FILLER_13_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_555 ();
 DECAPx1_ASAP7_75t_R FILLER_13_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_572 ();
 DECAPx6_ASAP7_75t_R FILLER_13_579 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_593 ();
 DECAPx2_ASAP7_75t_R FILLER_13_599 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_605 ();
 DECAPx2_ASAP7_75t_R FILLER_13_614 ();
 FILLER_ASAP7_75t_R FILLER_13_620 ();
 DECAPx4_ASAP7_75t_R FILLER_13_630 ();
 DECAPx10_ASAP7_75t_R FILLER_13_652 ();
 DECAPx2_ASAP7_75t_R FILLER_13_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_680 ();
 DECAPx2_ASAP7_75t_R FILLER_13_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_690 ();
 FILLER_ASAP7_75t_R FILLER_13_697 ();
 FILLER_ASAP7_75t_R FILLER_13_705 ();
 DECAPx2_ASAP7_75t_R FILLER_13_714 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_720 ();
 DECAPx4_ASAP7_75t_R FILLER_13_743 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_753 ();
 DECAPx2_ASAP7_75t_R FILLER_13_762 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_775 ();
 FILLER_ASAP7_75t_R FILLER_13_786 ();
 DECAPx4_ASAP7_75t_R FILLER_13_794 ();
 FILLER_ASAP7_75t_R FILLER_13_804 ();
 DECAPx4_ASAP7_75t_R FILLER_13_814 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_824 ();
 DECAPx6_ASAP7_75t_R FILLER_13_835 ();
 DECAPx6_ASAP7_75t_R FILLER_13_857 ();
 DECAPx10_ASAP7_75t_R FILLER_13_877 ();
 DECAPx1_ASAP7_75t_R FILLER_13_899 ();
 FILLER_ASAP7_75t_R FILLER_13_923 ();
 FILLER_ASAP7_75t_R FILLER_13_927 ();
 DECAPx6_ASAP7_75t_R FILLER_13_938 ();
 DECAPx1_ASAP7_75t_R FILLER_13_952 ();
 FILLER_ASAP7_75t_R FILLER_13_962 ();
 DECAPx1_ASAP7_75t_R FILLER_13_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_975 ();
 FILLER_ASAP7_75t_R FILLER_13_984 ();
 DECAPx6_ASAP7_75t_R FILLER_13_992 ();
 DECAPx2_ASAP7_75t_R FILLER_13_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1012 ();
 FILLER_ASAP7_75t_R FILLER_13_1033 ();
 FILLER_ASAP7_75t_R FILLER_13_1041 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_1049 ();
 DECAPx4_ASAP7_75t_R FILLER_13_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1068 ();
 DECAPx6_ASAP7_75t_R FILLER_13_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_13_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_13_1124 ();
 FILLER_ASAP7_75t_R FILLER_13_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1162 ();
 DECAPx1_ASAP7_75t_R FILLER_13_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1197 ();
 FILLER_ASAP7_75t_R FILLER_13_1219 ();
 DECAPx4_ASAP7_75t_R FILLER_13_1229 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_13_1355 ();
 DECAPx10_ASAP7_75t_R FILLER_14_2 ();
 DECAPx10_ASAP7_75t_R FILLER_14_24 ();
 DECAPx10_ASAP7_75t_R FILLER_14_46 ();
 DECAPx10_ASAP7_75t_R FILLER_14_68 ();
 DECAPx10_ASAP7_75t_R FILLER_14_90 ();
 DECAPx10_ASAP7_75t_R FILLER_14_112 ();
 DECAPx10_ASAP7_75t_R FILLER_14_134 ();
 DECAPx10_ASAP7_75t_R FILLER_14_156 ();
 DECAPx10_ASAP7_75t_R FILLER_14_178 ();
 DECAPx10_ASAP7_75t_R FILLER_14_200 ();
 DECAPx10_ASAP7_75t_R FILLER_14_222 ();
 DECAPx10_ASAP7_75t_R FILLER_14_244 ();
 DECAPx10_ASAP7_75t_R FILLER_14_266 ();
 DECAPx10_ASAP7_75t_R FILLER_14_288 ();
 DECAPx10_ASAP7_75t_R FILLER_14_310 ();
 DECAPx10_ASAP7_75t_R FILLER_14_332 ();
 DECAPx10_ASAP7_75t_R FILLER_14_354 ();
 DECAPx10_ASAP7_75t_R FILLER_14_376 ();
 DECAPx10_ASAP7_75t_R FILLER_14_398 ();
 DECAPx6_ASAP7_75t_R FILLER_14_420 ();
 DECAPx1_ASAP7_75t_R FILLER_14_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_438 ();
 DECAPx6_ASAP7_75t_R FILLER_14_446 ();
 FILLER_ASAP7_75t_R FILLER_14_460 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_14_464 ();
 DECAPx6_ASAP7_75t_R FILLER_14_479 ();
 DECAPx2_ASAP7_75t_R FILLER_14_499 ();
 FILLER_ASAP7_75t_R FILLER_14_505 ();
 FILLER_ASAP7_75t_R FILLER_14_527 ();
 DECAPx4_ASAP7_75t_R FILLER_14_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_545 ();
 DECAPx1_ASAP7_75t_R FILLER_14_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_557 ();
 FILLER_ASAP7_75t_R FILLER_14_578 ();
 FILLER_ASAP7_75t_R FILLER_14_588 ();
 FILLER_ASAP7_75t_R FILLER_14_597 ();
 FILLER_ASAP7_75t_R FILLER_14_605 ();
 DECAPx2_ASAP7_75t_R FILLER_14_615 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_14_621 ();
 DECAPx4_ASAP7_75t_R FILLER_14_631 ();
 FILLER_ASAP7_75t_R FILLER_14_641 ();
 DECAPx6_ASAP7_75t_R FILLER_14_663 ();
 DECAPx1_ASAP7_75t_R FILLER_14_689 ();
 DECAPx2_ASAP7_75t_R FILLER_14_699 ();
 FILLER_ASAP7_75t_R FILLER_14_705 ();
 DECAPx10_ASAP7_75t_R FILLER_14_715 ();
 DECAPx10_ASAP7_75t_R FILLER_14_737 ();
 DECAPx10_ASAP7_75t_R FILLER_14_759 ();
 DECAPx10_ASAP7_75t_R FILLER_14_781 ();
 DECAPx10_ASAP7_75t_R FILLER_14_803 ();
 DECAPx10_ASAP7_75t_R FILLER_14_825 ();
 DECAPx4_ASAP7_75t_R FILLER_14_847 ();
 DECAPx4_ASAP7_75t_R FILLER_14_863 ();
 FILLER_ASAP7_75t_R FILLER_14_873 ();
 FILLER_ASAP7_75t_R FILLER_14_881 ();
 FILLER_ASAP7_75t_R FILLER_14_895 ();
 DECAPx10_ASAP7_75t_R FILLER_14_903 ();
 FILLER_ASAP7_75t_R FILLER_14_925 ();
 DECAPx10_ASAP7_75t_R FILLER_14_933 ();
 DECAPx10_ASAP7_75t_R FILLER_14_955 ();
 DECAPx6_ASAP7_75t_R FILLER_14_977 ();
 DECAPx2_ASAP7_75t_R FILLER_14_991 ();
 FILLER_ASAP7_75t_R FILLER_14_1003 ();
 DECAPx4_ASAP7_75t_R FILLER_14_1011 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_14_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1054 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_14_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1087 ();
 DECAPx2_ASAP7_75t_R FILLER_14_1109 ();
 FILLER_ASAP7_75t_R FILLER_14_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_14_1145 ();
 DECAPx4_ASAP7_75t_R FILLER_14_1154 ();
 FILLER_ASAP7_75t_R FILLER_14_1164 ();
 DECAPx4_ASAP7_75t_R FILLER_14_1174 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_14_1184 ();
 DECAPx4_ASAP7_75t_R FILLER_14_1207 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_14_1217 ();
 FILLER_ASAP7_75t_R FILLER_14_1240 ();
 FILLER_ASAP7_75t_R FILLER_14_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_14_1343 ();
 DECAPx4_ASAP7_75t_R FILLER_14_1365 ();
 FILLER_ASAP7_75t_R FILLER_14_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_15_2 ();
 DECAPx10_ASAP7_75t_R FILLER_15_24 ();
 DECAPx10_ASAP7_75t_R FILLER_15_46 ();
 DECAPx10_ASAP7_75t_R FILLER_15_68 ();
 DECAPx10_ASAP7_75t_R FILLER_15_90 ();
 DECAPx10_ASAP7_75t_R FILLER_15_112 ();
 DECAPx10_ASAP7_75t_R FILLER_15_134 ();
 DECAPx10_ASAP7_75t_R FILLER_15_156 ();
 DECAPx10_ASAP7_75t_R FILLER_15_178 ();
 DECAPx10_ASAP7_75t_R FILLER_15_200 ();
 DECAPx10_ASAP7_75t_R FILLER_15_222 ();
 DECAPx10_ASAP7_75t_R FILLER_15_244 ();
 DECAPx10_ASAP7_75t_R FILLER_15_266 ();
 DECAPx10_ASAP7_75t_R FILLER_15_288 ();
 DECAPx10_ASAP7_75t_R FILLER_15_310 ();
 DECAPx10_ASAP7_75t_R FILLER_15_332 ();
 DECAPx10_ASAP7_75t_R FILLER_15_354 ();
 DECAPx10_ASAP7_75t_R FILLER_15_376 ();
 DECAPx10_ASAP7_75t_R FILLER_15_398 ();
 DECAPx2_ASAP7_75t_R FILLER_15_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_426 ();
 DECAPx2_ASAP7_75t_R FILLER_15_434 ();
 DECAPx10_ASAP7_75t_R FILLER_15_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_469 ();
 FILLER_ASAP7_75t_R FILLER_15_490 ();
 FILLER_ASAP7_75t_R FILLER_15_500 ();
 DECAPx1_ASAP7_75t_R FILLER_15_508 ();
 DECAPx1_ASAP7_75t_R FILLER_15_518 ();
 DECAPx10_ASAP7_75t_R FILLER_15_525 ();
 DECAPx6_ASAP7_75t_R FILLER_15_547 ();
 DECAPx10_ASAP7_75t_R FILLER_15_564 ();
 DECAPx6_ASAP7_75t_R FILLER_15_586 ();
 FILLER_ASAP7_75t_R FILLER_15_600 ();
 FILLER_ASAP7_75t_R FILLER_15_608 ();
 FILLER_ASAP7_75t_R FILLER_15_617 ();
 DECAPx6_ASAP7_75t_R FILLER_15_625 ();
 DECAPx1_ASAP7_75t_R FILLER_15_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_643 ();
 DECAPx2_ASAP7_75t_R FILLER_15_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_653 ();
 FILLER_ASAP7_75t_R FILLER_15_660 ();
 DECAPx1_ASAP7_75t_R FILLER_15_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_674 ();
 FILLER_ASAP7_75t_R FILLER_15_695 ();
 DECAPx4_ASAP7_75t_R FILLER_15_700 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_15_710 ();
 FILLER_ASAP7_75t_R FILLER_15_719 ();
 DECAPx2_ASAP7_75t_R FILLER_15_727 ();
 DECAPx4_ASAP7_75t_R FILLER_15_753 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_15_763 ();
 FILLER_ASAP7_75t_R FILLER_15_786 ();
 DECAPx6_ASAP7_75t_R FILLER_15_794 ();
 DECAPx1_ASAP7_75t_R FILLER_15_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_812 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_15_819 ();
 DECAPx6_ASAP7_75t_R FILLER_15_834 ();
 FILLER_ASAP7_75t_R FILLER_15_848 ();
 FILLER_ASAP7_75t_R FILLER_15_870 ();
 DECAPx2_ASAP7_75t_R FILLER_15_878 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_15_884 ();
 FILLER_ASAP7_75t_R FILLER_15_907 ();
 DECAPx4_ASAP7_75t_R FILLER_15_915 ();
 FILLER_ASAP7_75t_R FILLER_15_927 ();
 FILLER_ASAP7_75t_R FILLER_15_937 ();
 FILLER_ASAP7_75t_R FILLER_15_945 ();
 DECAPx2_ASAP7_75t_R FILLER_15_953 ();
 DECAPx4_ASAP7_75t_R FILLER_15_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_975 ();
 FILLER_ASAP7_75t_R FILLER_15_986 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1008 ();
 DECAPx6_ASAP7_75t_R FILLER_15_1030 ();
 FILLER_ASAP7_75t_R FILLER_15_1052 ();
 DECAPx1_ASAP7_75t_R FILLER_15_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1066 ();
 DECAPx1_ASAP7_75t_R FILLER_15_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1074 ();
 FILLER_ASAP7_75t_R FILLER_15_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_15_1103 ();
 FILLER_ASAP7_75t_R FILLER_15_1109 ();
 FILLER_ASAP7_75t_R FILLER_15_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1149 ();
 DECAPx1_ASAP7_75t_R FILLER_15_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1163 ();
 FILLER_ASAP7_75t_R FILLER_15_1184 ();
 DECAPx1_ASAP7_75t_R FILLER_15_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_15_1211 ();
 FILLER_ASAP7_75t_R FILLER_15_1217 ();
 DECAPx6_ASAP7_75t_R FILLER_15_1225 ();
 FILLER_ASAP7_75t_R FILLER_15_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_15_1337 ();
 DECAPx6_ASAP7_75t_R FILLER_15_1359 ();
 DECAPx1_ASAP7_75t_R FILLER_15_1373 ();
 DECAPx10_ASAP7_75t_R FILLER_16_2 ();
 DECAPx10_ASAP7_75t_R FILLER_16_24 ();
 DECAPx10_ASAP7_75t_R FILLER_16_46 ();
 DECAPx10_ASAP7_75t_R FILLER_16_68 ();
 DECAPx10_ASAP7_75t_R FILLER_16_90 ();
 DECAPx10_ASAP7_75t_R FILLER_16_112 ();
 DECAPx10_ASAP7_75t_R FILLER_16_134 ();
 DECAPx10_ASAP7_75t_R FILLER_16_156 ();
 DECAPx10_ASAP7_75t_R FILLER_16_178 ();
 DECAPx10_ASAP7_75t_R FILLER_16_200 ();
 DECAPx10_ASAP7_75t_R FILLER_16_222 ();
 DECAPx10_ASAP7_75t_R FILLER_16_244 ();
 DECAPx10_ASAP7_75t_R FILLER_16_266 ();
 DECAPx10_ASAP7_75t_R FILLER_16_288 ();
 DECAPx10_ASAP7_75t_R FILLER_16_310 ();
 DECAPx10_ASAP7_75t_R FILLER_16_332 ();
 DECAPx10_ASAP7_75t_R FILLER_16_354 ();
 DECAPx10_ASAP7_75t_R FILLER_16_376 ();
 DECAPx10_ASAP7_75t_R FILLER_16_398 ();
 FILLER_ASAP7_75t_R FILLER_16_440 ();
 FILLER_ASAP7_75t_R FILLER_16_448 ();
 DECAPx1_ASAP7_75t_R FILLER_16_458 ();
 DECAPx2_ASAP7_75t_R FILLER_16_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_470 ();
 DECAPx1_ASAP7_75t_R FILLER_16_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_478 ();
 DECAPx2_ASAP7_75t_R FILLER_16_485 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_16_491 ();
 FILLER_ASAP7_75t_R FILLER_16_500 ();
 DECAPx1_ASAP7_75t_R FILLER_16_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_514 ();
 DECAPx4_ASAP7_75t_R FILLER_16_521 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_16_531 ();
 DECAPx10_ASAP7_75t_R FILLER_16_541 ();
 DECAPx6_ASAP7_75t_R FILLER_16_563 ();
 DECAPx2_ASAP7_75t_R FILLER_16_577 ();
 FILLER_ASAP7_75t_R FILLER_16_590 ();
 DECAPx10_ASAP7_75t_R FILLER_16_598 ();
 DECAPx2_ASAP7_75t_R FILLER_16_620 ();
 FILLER_ASAP7_75t_R FILLER_16_626 ();
 DECAPx4_ASAP7_75t_R FILLER_16_635 ();
 FILLER_ASAP7_75t_R FILLER_16_645 ();
 DECAPx10_ASAP7_75t_R FILLER_16_653 ();
 DECAPx6_ASAP7_75t_R FILLER_16_675 ();
 DECAPx2_ASAP7_75t_R FILLER_16_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_695 ();
 FILLER_ASAP7_75t_R FILLER_16_702 ();
 FILLER_ASAP7_75t_R FILLER_16_712 ();
 FILLER_ASAP7_75t_R FILLER_16_720 ();
 DECAPx1_ASAP7_75t_R FILLER_16_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_742 ();
 FILLER_ASAP7_75t_R FILLER_16_751 ();
 DECAPx2_ASAP7_75t_R FILLER_16_759 ();
 FILLER_ASAP7_75t_R FILLER_16_774 ();
 FILLER_ASAP7_75t_R FILLER_16_782 ();
 DECAPx1_ASAP7_75t_R FILLER_16_790 ();
 FILLER_ASAP7_75t_R FILLER_16_814 ();
 FILLER_ASAP7_75t_R FILLER_16_828 ();
 FILLER_ASAP7_75t_R FILLER_16_839 ();
 FILLER_ASAP7_75t_R FILLER_16_847 ();
 FILLER_ASAP7_75t_R FILLER_16_855 ();
 DECAPx1_ASAP7_75t_R FILLER_16_863 ();
 DECAPx1_ASAP7_75t_R FILLER_16_875 ();
 FILLER_ASAP7_75t_R FILLER_16_891 ();
 DECAPx6_ASAP7_75t_R FILLER_16_899 ();
 DECAPx2_ASAP7_75t_R FILLER_16_913 ();
 FILLER_ASAP7_75t_R FILLER_16_939 ();
 DECAPx4_ASAP7_75t_R FILLER_16_949 ();
 DECAPx2_ASAP7_75t_R FILLER_16_979 ();
 DECAPx2_ASAP7_75t_R FILLER_16_1007 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_16_1013 ();
 FILLER_ASAP7_75t_R FILLER_16_1028 ();
 FILLER_ASAP7_75t_R FILLER_16_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_16_1043 ();
 FILLER_ASAP7_75t_R FILLER_16_1067 ();
 FILLER_ASAP7_75t_R FILLER_16_1077 ();
 FILLER_ASAP7_75t_R FILLER_16_1086 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_16_1094 ();
 FILLER_ASAP7_75t_R FILLER_16_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_16_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_16_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1141 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_16_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_16_1154 ();
 FILLER_ASAP7_75t_R FILLER_16_1166 ();
 DECAPx6_ASAP7_75t_R FILLER_16_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_1188 ();
 DECAPx2_ASAP7_75t_R FILLER_16_1195 ();
 FILLER_ASAP7_75t_R FILLER_16_1201 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_16_1206 ();
 FILLER_ASAP7_75t_R FILLER_16_1215 ();
 FILLER_ASAP7_75t_R FILLER_16_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_16_1342 ();
 DECAPx4_ASAP7_75t_R FILLER_16_1364 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_16_1374 ();
 DECAPx10_ASAP7_75t_R FILLER_17_2 ();
 DECAPx10_ASAP7_75t_R FILLER_17_24 ();
 DECAPx10_ASAP7_75t_R FILLER_17_46 ();
 DECAPx10_ASAP7_75t_R FILLER_17_68 ();
 DECAPx10_ASAP7_75t_R FILLER_17_90 ();
 DECAPx10_ASAP7_75t_R FILLER_17_112 ();
 DECAPx10_ASAP7_75t_R FILLER_17_134 ();
 DECAPx10_ASAP7_75t_R FILLER_17_156 ();
 DECAPx10_ASAP7_75t_R FILLER_17_178 ();
 DECAPx10_ASAP7_75t_R FILLER_17_200 ();
 DECAPx10_ASAP7_75t_R FILLER_17_222 ();
 DECAPx10_ASAP7_75t_R FILLER_17_244 ();
 DECAPx10_ASAP7_75t_R FILLER_17_266 ();
 DECAPx10_ASAP7_75t_R FILLER_17_288 ();
 DECAPx10_ASAP7_75t_R FILLER_17_310 ();
 DECAPx10_ASAP7_75t_R FILLER_17_332 ();
 DECAPx10_ASAP7_75t_R FILLER_17_354 ();
 DECAPx10_ASAP7_75t_R FILLER_17_376 ();
 DECAPx10_ASAP7_75t_R FILLER_17_398 ();
 DECAPx2_ASAP7_75t_R FILLER_17_420 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_17_426 ();
 DECAPx4_ASAP7_75t_R FILLER_17_435 ();
 FILLER_ASAP7_75t_R FILLER_17_445 ();
 DECAPx10_ASAP7_75t_R FILLER_17_467 ();
 DECAPx6_ASAP7_75t_R FILLER_17_489 ();
 DECAPx1_ASAP7_75t_R FILLER_17_503 ();
 DECAPx1_ASAP7_75t_R FILLER_17_514 ();
 DECAPx4_ASAP7_75t_R FILLER_17_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_535 ();
 FILLER_ASAP7_75t_R FILLER_17_543 ();
 DECAPx2_ASAP7_75t_R FILLER_17_551 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_17_557 ();
 DECAPx2_ASAP7_75t_R FILLER_17_567 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_17_573 ();
 FILLER_ASAP7_75t_R FILLER_17_596 ();
 DECAPx1_ASAP7_75t_R FILLER_17_604 ();
 DECAPx4_ASAP7_75t_R FILLER_17_615 ();
 DECAPx1_ASAP7_75t_R FILLER_17_645 ();
 DECAPx2_ASAP7_75t_R FILLER_17_655 ();
 FILLER_ASAP7_75t_R FILLER_17_661 ();
 FILLER_ASAP7_75t_R FILLER_17_671 ();
 DECAPx10_ASAP7_75t_R FILLER_17_680 ();
 DECAPx10_ASAP7_75t_R FILLER_17_702 ();
 DECAPx4_ASAP7_75t_R FILLER_17_724 ();
 FILLER_ASAP7_75t_R FILLER_17_734 ();
 FILLER_ASAP7_75t_R FILLER_17_745 ();
 DECAPx4_ASAP7_75t_R FILLER_17_753 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_17_763 ();
 DECAPx2_ASAP7_75t_R FILLER_17_774 ();
 DECAPx6_ASAP7_75t_R FILLER_17_796 ();
 DECAPx1_ASAP7_75t_R FILLER_17_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_814 ();
 FILLER_ASAP7_75t_R FILLER_17_821 ();
 FILLER_ASAP7_75t_R FILLER_17_829 ();
 FILLER_ASAP7_75t_R FILLER_17_834 ();
 DECAPx2_ASAP7_75t_R FILLER_17_844 ();
 DECAPx10_ASAP7_75t_R FILLER_17_858 ();
 DECAPx10_ASAP7_75t_R FILLER_17_880 ();
 DECAPx2_ASAP7_75t_R FILLER_17_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_908 ();
 DECAPx2_ASAP7_75t_R FILLER_17_917 ();
 FILLER_ASAP7_75t_R FILLER_17_923 ();
 DECAPx6_ASAP7_75t_R FILLER_17_927 ();
 FILLER_ASAP7_75t_R FILLER_17_941 ();
 DECAPx2_ASAP7_75t_R FILLER_17_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_955 ();
 FILLER_ASAP7_75t_R FILLER_17_963 ();
 DECAPx6_ASAP7_75t_R FILLER_17_971 ();
 DECAPx1_ASAP7_75t_R FILLER_17_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_989 ();
 FILLER_ASAP7_75t_R FILLER_17_998 ();
 FILLER_ASAP7_75t_R FILLER_17_1006 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_17_1011 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_17_1020 ();
 DECAPx1_ASAP7_75t_R FILLER_17_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1059 ();
 DECAPx6_ASAP7_75t_R FILLER_17_1081 ();
 DECAPx1_ASAP7_75t_R FILLER_17_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_17_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_1108 ();
 FILLER_ASAP7_75t_R FILLER_17_1115 ();
 DECAPx6_ASAP7_75t_R FILLER_17_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_17_1199 ();
 FILLER_ASAP7_75t_R FILLER_17_1205 ();
 FILLER_ASAP7_75t_R FILLER_17_1210 ();
 FILLER_ASAP7_75t_R FILLER_17_1221 ();
 FILLER_ASAP7_75t_R FILLER_17_1235 ();
 FILLER_ASAP7_75t_R FILLER_17_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_17_1343 ();
 DECAPx4_ASAP7_75t_R FILLER_17_1365 ();
 FILLER_ASAP7_75t_R FILLER_17_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_18_2 ();
 DECAPx10_ASAP7_75t_R FILLER_18_24 ();
 DECAPx10_ASAP7_75t_R FILLER_18_46 ();
 DECAPx10_ASAP7_75t_R FILLER_18_68 ();
 DECAPx10_ASAP7_75t_R FILLER_18_90 ();
 DECAPx10_ASAP7_75t_R FILLER_18_112 ();
 DECAPx10_ASAP7_75t_R FILLER_18_134 ();
 DECAPx10_ASAP7_75t_R FILLER_18_156 ();
 DECAPx10_ASAP7_75t_R FILLER_18_178 ();
 DECAPx10_ASAP7_75t_R FILLER_18_200 ();
 DECAPx10_ASAP7_75t_R FILLER_18_222 ();
 DECAPx10_ASAP7_75t_R FILLER_18_244 ();
 DECAPx10_ASAP7_75t_R FILLER_18_266 ();
 DECAPx10_ASAP7_75t_R FILLER_18_288 ();
 DECAPx10_ASAP7_75t_R FILLER_18_310 ();
 DECAPx10_ASAP7_75t_R FILLER_18_332 ();
 DECAPx10_ASAP7_75t_R FILLER_18_354 ();
 DECAPx10_ASAP7_75t_R FILLER_18_376 ();
 DECAPx10_ASAP7_75t_R FILLER_18_398 ();
 DECAPx10_ASAP7_75t_R FILLER_18_420 ();
 DECAPx1_ASAP7_75t_R FILLER_18_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_446 ();
 DECAPx2_ASAP7_75t_R FILLER_18_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_18_459 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_18_464 ();
 DECAPx6_ASAP7_75t_R FILLER_18_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_493 ();
 DECAPx10_ASAP7_75t_R FILLER_18_500 ();
 DECAPx1_ASAP7_75t_R FILLER_18_522 ();
 DECAPx1_ASAP7_75t_R FILLER_18_546 ();
 FILLER_ASAP7_75t_R FILLER_18_570 ();
 DECAPx4_ASAP7_75t_R FILLER_18_578 ();
 DECAPx2_ASAP7_75t_R FILLER_18_595 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_18_601 ();
 DECAPx6_ASAP7_75t_R FILLER_18_624 ();
 FILLER_ASAP7_75t_R FILLER_18_638 ();
 DECAPx2_ASAP7_75t_R FILLER_18_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_653 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_18_661 ();
 DECAPx2_ASAP7_75t_R FILLER_18_671 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_18_677 ();
 FILLER_ASAP7_75t_R FILLER_18_686 ();
 DECAPx10_ASAP7_75t_R FILLER_18_694 ();
 DECAPx1_ASAP7_75t_R FILLER_18_716 ();
 DECAPx10_ASAP7_75t_R FILLER_18_726 ();
 DECAPx6_ASAP7_75t_R FILLER_18_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_762 ();
 DECAPx10_ASAP7_75t_R FILLER_18_775 ();
 DECAPx4_ASAP7_75t_R FILLER_18_797 ();
 DECAPx10_ASAP7_75t_R FILLER_18_810 ();
 FILLER_ASAP7_75t_R FILLER_18_832 ();
 DECAPx4_ASAP7_75t_R FILLER_18_854 ();
 DECAPx4_ASAP7_75t_R FILLER_18_876 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_18_886 ();
 FILLER_ASAP7_75t_R FILLER_18_895 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_18_903 ();
 DECAPx6_ASAP7_75t_R FILLER_18_926 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_18_946 ();
 FILLER_ASAP7_75t_R FILLER_18_952 ();
 DECAPx4_ASAP7_75t_R FILLER_18_963 ();
 FILLER_ASAP7_75t_R FILLER_18_973 ();
 DECAPx4_ASAP7_75t_R FILLER_18_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_991 ();
 DECAPx2_ASAP7_75t_R FILLER_18_998 ();
 FILLER_ASAP7_75t_R FILLER_18_1004 ();
 FILLER_ASAP7_75t_R FILLER_18_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_18_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_18_1058 ();
 FILLER_ASAP7_75t_R FILLER_18_1064 ();
 DECAPx6_ASAP7_75t_R FILLER_18_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1096 ();
 DECAPx6_ASAP7_75t_R FILLER_18_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_18_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1138 ();
 DECAPx1_ASAP7_75t_R FILLER_18_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_18_1158 ();
 FILLER_ASAP7_75t_R FILLER_18_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_18_1180 ();
 FILLER_ASAP7_75t_R FILLER_18_1187 ();
 DECAPx6_ASAP7_75t_R FILLER_18_1198 ();
 DECAPx6_ASAP7_75t_R FILLER_18_1215 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_18_1229 ();
 FILLER_ASAP7_75t_R FILLER_18_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_18_1345 ();
 DECAPx4_ASAP7_75t_R FILLER_18_1367 ();
 DECAPx10_ASAP7_75t_R FILLER_19_2 ();
 DECAPx10_ASAP7_75t_R FILLER_19_24 ();
 DECAPx10_ASAP7_75t_R FILLER_19_46 ();
 DECAPx10_ASAP7_75t_R FILLER_19_68 ();
 DECAPx10_ASAP7_75t_R FILLER_19_90 ();
 DECAPx10_ASAP7_75t_R FILLER_19_112 ();
 DECAPx10_ASAP7_75t_R FILLER_19_134 ();
 DECAPx10_ASAP7_75t_R FILLER_19_156 ();
 DECAPx10_ASAP7_75t_R FILLER_19_178 ();
 DECAPx10_ASAP7_75t_R FILLER_19_200 ();
 DECAPx10_ASAP7_75t_R FILLER_19_222 ();
 DECAPx10_ASAP7_75t_R FILLER_19_244 ();
 DECAPx10_ASAP7_75t_R FILLER_19_266 ();
 DECAPx10_ASAP7_75t_R FILLER_19_288 ();
 DECAPx10_ASAP7_75t_R FILLER_19_310 ();
 DECAPx10_ASAP7_75t_R FILLER_19_332 ();
 DECAPx10_ASAP7_75t_R FILLER_19_354 ();
 DECAPx10_ASAP7_75t_R FILLER_19_376 ();
 DECAPx10_ASAP7_75t_R FILLER_19_398 ();
 DECAPx2_ASAP7_75t_R FILLER_19_420 ();
 FILLER_ASAP7_75t_R FILLER_19_426 ();
 DECAPx1_ASAP7_75t_R FILLER_19_435 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_19_445 ();
 DECAPx4_ASAP7_75t_R FILLER_19_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_464 ();
 FILLER_ASAP7_75t_R FILLER_19_468 ();
 FILLER_ASAP7_75t_R FILLER_19_490 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_19_495 ();
 FILLER_ASAP7_75t_R FILLER_19_504 ();
 DECAPx10_ASAP7_75t_R FILLER_19_512 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_19_534 ();
 DECAPx6_ASAP7_75t_R FILLER_19_543 ();
 DECAPx1_ASAP7_75t_R FILLER_19_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_561 ();
 FILLER_ASAP7_75t_R FILLER_19_569 ();
 DECAPx2_ASAP7_75t_R FILLER_19_577 ();
 FILLER_ASAP7_75t_R FILLER_19_591 ();
 DECAPx4_ASAP7_75t_R FILLER_19_599 ();
 FILLER_ASAP7_75t_R FILLER_19_609 ();
 DECAPx6_ASAP7_75t_R FILLER_19_617 ();
 DECAPx2_ASAP7_75t_R FILLER_19_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_637 ();
 DECAPx1_ASAP7_75t_R FILLER_19_644 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_19_651 ();
 DECAPx2_ASAP7_75t_R FILLER_19_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_680 ();
 FILLER_ASAP7_75t_R FILLER_19_687 ();
 DECAPx1_ASAP7_75t_R FILLER_19_697 ();
 FILLER_ASAP7_75t_R FILLER_19_709 ();
 DECAPx1_ASAP7_75t_R FILLER_19_717 ();
 DECAPx6_ASAP7_75t_R FILLER_19_737 ();
 DECAPx1_ASAP7_75t_R FILLER_19_751 ();
 DECAPx6_ASAP7_75t_R FILLER_19_762 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_19_776 ();
 DECAPx6_ASAP7_75t_R FILLER_19_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_799 ();
 FILLER_ASAP7_75t_R FILLER_19_804 ();
 DECAPx10_ASAP7_75t_R FILLER_19_816 ();
 DECAPx10_ASAP7_75t_R FILLER_19_838 ();
 DECAPx4_ASAP7_75t_R FILLER_19_860 ();
 FILLER_ASAP7_75t_R FILLER_19_870 ();
 FILLER_ASAP7_75t_R FILLER_19_892 ();
 DECAPx2_ASAP7_75t_R FILLER_19_900 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_19_906 ();
 FILLER_ASAP7_75t_R FILLER_19_915 ();
 FILLER_ASAP7_75t_R FILLER_19_923 ();
 DECAPx10_ASAP7_75t_R FILLER_19_927 ();
 DECAPx1_ASAP7_75t_R FILLER_19_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_953 ();
 DECAPx2_ASAP7_75t_R FILLER_19_957 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_19_963 ();
 FILLER_ASAP7_75t_R FILLER_19_978 ();
 DECAPx6_ASAP7_75t_R FILLER_19_988 ();
 DECAPx1_ASAP7_75t_R FILLER_19_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_19_1010 ();
 DECAPx1_ASAP7_75t_R FILLER_19_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_19_1035 ();
 DECAPx1_ASAP7_75t_R FILLER_19_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_19_1057 ();
 FILLER_ASAP7_75t_R FILLER_19_1063 ();
 FILLER_ASAP7_75t_R FILLER_19_1073 ();
 FILLER_ASAP7_75t_R FILLER_19_1095 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_19_1103 ();
 DECAPx2_ASAP7_75t_R FILLER_19_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1115 ();
 FILLER_ASAP7_75t_R FILLER_19_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_19_1132 ();
 FILLER_ASAP7_75t_R FILLER_19_1156 ();
 DECAPx1_ASAP7_75t_R FILLER_19_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_1170 ();
 FILLER_ASAP7_75t_R FILLER_19_1191 ();
 DECAPx4_ASAP7_75t_R FILLER_19_1196 ();
 FILLER_ASAP7_75t_R FILLER_19_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_19_1346 ();
 DECAPx2_ASAP7_75t_R FILLER_19_1368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_19_1374 ();
 DECAPx10_ASAP7_75t_R FILLER_20_2 ();
 DECAPx10_ASAP7_75t_R FILLER_20_24 ();
 DECAPx10_ASAP7_75t_R FILLER_20_46 ();
 DECAPx10_ASAP7_75t_R FILLER_20_68 ();
 DECAPx10_ASAP7_75t_R FILLER_20_90 ();
 DECAPx10_ASAP7_75t_R FILLER_20_112 ();
 DECAPx10_ASAP7_75t_R FILLER_20_134 ();
 DECAPx10_ASAP7_75t_R FILLER_20_156 ();
 DECAPx10_ASAP7_75t_R FILLER_20_178 ();
 DECAPx10_ASAP7_75t_R FILLER_20_200 ();
 DECAPx10_ASAP7_75t_R FILLER_20_222 ();
 DECAPx10_ASAP7_75t_R FILLER_20_244 ();
 DECAPx10_ASAP7_75t_R FILLER_20_266 ();
 DECAPx10_ASAP7_75t_R FILLER_20_288 ();
 DECAPx10_ASAP7_75t_R FILLER_20_310 ();
 DECAPx10_ASAP7_75t_R FILLER_20_332 ();
 DECAPx10_ASAP7_75t_R FILLER_20_354 ();
 DECAPx10_ASAP7_75t_R FILLER_20_376 ();
 DECAPx10_ASAP7_75t_R FILLER_20_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_420 ();
 FILLER_ASAP7_75t_R FILLER_20_441 ();
 FILLER_ASAP7_75t_R FILLER_20_450 ();
 FILLER_ASAP7_75t_R FILLER_20_460 ();
 DECAPx10_ASAP7_75t_R FILLER_20_464 ();
 DECAPx4_ASAP7_75t_R FILLER_20_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_496 ();
 FILLER_ASAP7_75t_R FILLER_20_503 ();
 DECAPx10_ASAP7_75t_R FILLER_20_512 ();
 FILLER_ASAP7_75t_R FILLER_20_542 ();
 DECAPx10_ASAP7_75t_R FILLER_20_550 ();
 DECAPx2_ASAP7_75t_R FILLER_20_572 ();
 FILLER_ASAP7_75t_R FILLER_20_578 ();
 DECAPx2_ASAP7_75t_R FILLER_20_600 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_606 ();
 FILLER_ASAP7_75t_R FILLER_20_616 ();
 DECAPx1_ASAP7_75t_R FILLER_20_624 ();
 DECAPx10_ASAP7_75t_R FILLER_20_636 ();
 DECAPx2_ASAP7_75t_R FILLER_20_658 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_664 ();
 DECAPx4_ASAP7_75t_R FILLER_20_673 ();
 FILLER_ASAP7_75t_R FILLER_20_683 ();
 DECAPx10_ASAP7_75t_R FILLER_20_691 ();
 DECAPx6_ASAP7_75t_R FILLER_20_713 ();
 DECAPx1_ASAP7_75t_R FILLER_20_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_731 ();
 FILLER_ASAP7_75t_R FILLER_20_741 ();
 DECAPx1_ASAP7_75t_R FILLER_20_749 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_773 ();
 FILLER_ASAP7_75t_R FILLER_20_802 ();
 DECAPx1_ASAP7_75t_R FILLER_20_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_834 ();
 DECAPx10_ASAP7_75t_R FILLER_20_838 ();
 DECAPx1_ASAP7_75t_R FILLER_20_860 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_870 ();
 DECAPx10_ASAP7_75t_R FILLER_20_879 ();
 DECAPx4_ASAP7_75t_R FILLER_20_901 ();
 DECAPx6_ASAP7_75t_R FILLER_20_914 ();
 FILLER_ASAP7_75t_R FILLER_20_940 ();
 DECAPx6_ASAP7_75t_R FILLER_20_950 ();
 DECAPx1_ASAP7_75t_R FILLER_20_970 ();
 DECAPx4_ASAP7_75t_R FILLER_20_994 ();
 FILLER_ASAP7_75t_R FILLER_20_1004 ();
 FILLER_ASAP7_75t_R FILLER_20_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1027 ();
 FILLER_ASAP7_75t_R FILLER_20_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1046 ();
 FILLER_ASAP7_75t_R FILLER_20_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1069 ();
 FILLER_ASAP7_75t_R FILLER_20_1075 ();
 DECAPx4_ASAP7_75t_R FILLER_20_1085 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_1095 ();
 FILLER_ASAP7_75t_R FILLER_20_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_1121 ();
 DECAPx4_ASAP7_75t_R FILLER_20_1142 ();
 FILLER_ASAP7_75t_R FILLER_20_1152 ();
 DECAPx4_ASAP7_75t_R FILLER_20_1157 ();
 FILLER_ASAP7_75t_R FILLER_20_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1180 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_1186 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1195 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_1201 ();
 FILLER_ASAP7_75t_R FILLER_20_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1215 ();
 FILLER_ASAP7_75t_R FILLER_20_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_20_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_20_1369 ();
 FILLER_ASAP7_75t_R FILLER_20_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_21_2 ();
 DECAPx10_ASAP7_75t_R FILLER_21_24 ();
 DECAPx10_ASAP7_75t_R FILLER_21_46 ();
 DECAPx10_ASAP7_75t_R FILLER_21_68 ();
 DECAPx10_ASAP7_75t_R FILLER_21_90 ();
 DECAPx10_ASAP7_75t_R FILLER_21_112 ();
 DECAPx10_ASAP7_75t_R FILLER_21_134 ();
 DECAPx10_ASAP7_75t_R FILLER_21_156 ();
 DECAPx10_ASAP7_75t_R FILLER_21_178 ();
 DECAPx10_ASAP7_75t_R FILLER_21_200 ();
 DECAPx10_ASAP7_75t_R FILLER_21_222 ();
 DECAPx10_ASAP7_75t_R FILLER_21_244 ();
 DECAPx10_ASAP7_75t_R FILLER_21_266 ();
 DECAPx10_ASAP7_75t_R FILLER_21_288 ();
 DECAPx10_ASAP7_75t_R FILLER_21_310 ();
 DECAPx10_ASAP7_75t_R FILLER_21_332 ();
 DECAPx10_ASAP7_75t_R FILLER_21_354 ();
 DECAPx10_ASAP7_75t_R FILLER_21_376 ();
 DECAPx10_ASAP7_75t_R FILLER_21_398 ();
 DECAPx4_ASAP7_75t_R FILLER_21_420 ();
 FILLER_ASAP7_75t_R FILLER_21_430 ();
 DECAPx6_ASAP7_75t_R FILLER_21_438 ();
 FILLER_ASAP7_75t_R FILLER_21_452 ();
 DECAPx10_ASAP7_75t_R FILLER_21_474 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_21_496 ();
 DECAPx4_ASAP7_75t_R FILLER_21_507 ();
 DECAPx2_ASAP7_75t_R FILLER_21_524 ();
 DECAPx2_ASAP7_75t_R FILLER_21_550 ();
 FILLER_ASAP7_75t_R FILLER_21_556 ();
 FILLER_ASAP7_75t_R FILLER_21_566 ();
 DECAPx10_ASAP7_75t_R FILLER_21_574 ();
 DECAPx10_ASAP7_75t_R FILLER_21_596 ();
 DECAPx1_ASAP7_75t_R FILLER_21_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_622 ();
 DECAPx2_ASAP7_75t_R FILLER_21_643 ();
 FILLER_ASAP7_75t_R FILLER_21_649 ();
 FILLER_ASAP7_75t_R FILLER_21_658 ();
 DECAPx1_ASAP7_75t_R FILLER_21_666 ();
 FILLER_ASAP7_75t_R FILLER_21_677 ();
 DECAPx2_ASAP7_75t_R FILLER_21_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_691 ();
 DECAPx2_ASAP7_75t_R FILLER_21_698 ();
 DECAPx10_ASAP7_75t_R FILLER_21_711 ();
 DECAPx1_ASAP7_75t_R FILLER_21_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_737 ();
 FILLER_ASAP7_75t_R FILLER_21_746 ();
 DECAPx2_ASAP7_75t_R FILLER_21_754 ();
 DECAPx4_ASAP7_75t_R FILLER_21_766 ();
 FILLER_ASAP7_75t_R FILLER_21_776 ();
 FILLER_ASAP7_75t_R FILLER_21_784 ();
 FILLER_ASAP7_75t_R FILLER_21_808 ();
 DECAPx1_ASAP7_75t_R FILLER_21_816 ();
 FILLER_ASAP7_75t_R FILLER_21_846 ();
 FILLER_ASAP7_75t_R FILLER_21_854 ();
 DECAPx10_ASAP7_75t_R FILLER_21_859 ();
 DECAPx10_ASAP7_75t_R FILLER_21_881 ();
 FILLER_ASAP7_75t_R FILLER_21_903 ();
 FILLER_ASAP7_75t_R FILLER_21_908 ();
 DECAPx2_ASAP7_75t_R FILLER_21_919 ();
 DECAPx2_ASAP7_75t_R FILLER_21_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_933 ();
 DECAPx10_ASAP7_75t_R FILLER_21_954 ();
 DECAPx10_ASAP7_75t_R FILLER_21_976 ();
 DECAPx2_ASAP7_75t_R FILLER_21_998 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_21_1004 ();
 DECAPx6_ASAP7_75t_R FILLER_21_1010 ();
 FILLER_ASAP7_75t_R FILLER_21_1024 ();
 FILLER_ASAP7_75t_R FILLER_21_1046 ();
 FILLER_ASAP7_75t_R FILLER_21_1054 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_21_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1068 ();
 DECAPx6_ASAP7_75t_R FILLER_21_1090 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_21_1104 ();
 DECAPx4_ASAP7_75t_R FILLER_21_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1171 ();
 DECAPx6_ASAP7_75t_R FILLER_21_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1207 ();
 FILLER_ASAP7_75t_R FILLER_21_1217 ();
 DECAPx1_ASAP7_75t_R FILLER_21_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_21_1338 ();
 DECAPx6_ASAP7_75t_R FILLER_21_1360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_21_1374 ();
 DECAPx10_ASAP7_75t_R FILLER_22_2 ();
 DECAPx10_ASAP7_75t_R FILLER_22_24 ();
 DECAPx10_ASAP7_75t_R FILLER_22_46 ();
 DECAPx10_ASAP7_75t_R FILLER_22_68 ();
 DECAPx10_ASAP7_75t_R FILLER_22_90 ();
 DECAPx10_ASAP7_75t_R FILLER_22_112 ();
 DECAPx10_ASAP7_75t_R FILLER_22_134 ();
 DECAPx10_ASAP7_75t_R FILLER_22_156 ();
 DECAPx10_ASAP7_75t_R FILLER_22_178 ();
 DECAPx10_ASAP7_75t_R FILLER_22_200 ();
 DECAPx10_ASAP7_75t_R FILLER_22_222 ();
 DECAPx10_ASAP7_75t_R FILLER_22_244 ();
 DECAPx10_ASAP7_75t_R FILLER_22_266 ();
 DECAPx10_ASAP7_75t_R FILLER_22_288 ();
 DECAPx10_ASAP7_75t_R FILLER_22_310 ();
 DECAPx10_ASAP7_75t_R FILLER_22_332 ();
 DECAPx10_ASAP7_75t_R FILLER_22_354 ();
 DECAPx10_ASAP7_75t_R FILLER_22_376 ();
 DECAPx10_ASAP7_75t_R FILLER_22_398 ();
 DECAPx10_ASAP7_75t_R FILLER_22_420 ();
 DECAPx6_ASAP7_75t_R FILLER_22_442 ();
 DECAPx2_ASAP7_75t_R FILLER_22_456 ();
 DECAPx2_ASAP7_75t_R FILLER_22_464 ();
 FILLER_ASAP7_75t_R FILLER_22_473 ();
 DECAPx4_ASAP7_75t_R FILLER_22_487 ();
 DECAPx2_ASAP7_75t_R FILLER_22_503 ();
 DECAPx4_ASAP7_75t_R FILLER_22_529 ();
 DECAPx4_ASAP7_75t_R FILLER_22_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_552 ();
 DECAPx2_ASAP7_75t_R FILLER_22_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_579 ();
 DECAPx6_ASAP7_75t_R FILLER_22_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_606 ();
 FILLER_ASAP7_75t_R FILLER_22_615 ();
 DECAPx2_ASAP7_75t_R FILLER_22_623 ();
 DECAPx4_ASAP7_75t_R FILLER_22_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_642 ();
 DECAPx4_ASAP7_75t_R FILLER_22_663 ();
 DECAPx2_ASAP7_75t_R FILLER_22_679 ();
 FILLER_ASAP7_75t_R FILLER_22_685 ();
 DECAPx1_ASAP7_75t_R FILLER_22_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_699 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_22_720 ();
 DECAPx4_ASAP7_75t_R FILLER_22_743 ();
 FILLER_ASAP7_75t_R FILLER_22_757 ();
 DECAPx6_ASAP7_75t_R FILLER_22_769 ();
 FILLER_ASAP7_75t_R FILLER_22_787 ();
 FILLER_ASAP7_75t_R FILLER_22_796 ();
 DECAPx2_ASAP7_75t_R FILLER_22_801 ();
 FILLER_ASAP7_75t_R FILLER_22_807 ();
 FILLER_ASAP7_75t_R FILLER_22_817 ();
 FILLER_ASAP7_75t_R FILLER_22_822 ();
 DECAPx2_ASAP7_75t_R FILLER_22_827 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_22_833 ();
 DECAPx2_ASAP7_75t_R FILLER_22_843 ();
 FILLER_ASAP7_75t_R FILLER_22_852 ();
 FILLER_ASAP7_75t_R FILLER_22_863 ();
 DECAPx2_ASAP7_75t_R FILLER_22_871 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_22_877 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_22_883 ();
 FILLER_ASAP7_75t_R FILLER_22_893 ();
 DECAPx10_ASAP7_75t_R FILLER_22_901 ();
 DECAPx1_ASAP7_75t_R FILLER_22_923 ();
 FILLER_ASAP7_75t_R FILLER_22_933 ();
 DECAPx6_ASAP7_75t_R FILLER_22_941 ();
 FILLER_ASAP7_75t_R FILLER_22_955 ();
 FILLER_ASAP7_75t_R FILLER_22_965 ();
 FILLER_ASAP7_75t_R FILLER_22_973 ();
 DECAPx4_ASAP7_75t_R FILLER_22_981 ();
 FILLER_ASAP7_75t_R FILLER_22_991 ();
 DECAPx4_ASAP7_75t_R FILLER_22_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_22_1060 ();
 DECAPx2_ASAP7_75t_R FILLER_22_1072 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_22_1078 ();
 DECAPx6_ASAP7_75t_R FILLER_22_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_22_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1109 ();
 DECAPx6_ASAP7_75t_R FILLER_22_1118 ();
 DECAPx1_ASAP7_75t_R FILLER_22_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_22_1144 ();
 DECAPx4_ASAP7_75t_R FILLER_22_1154 ();
 FILLER_ASAP7_75t_R FILLER_22_1172 ();
 DECAPx4_ASAP7_75t_R FILLER_22_1177 ();
 FILLER_ASAP7_75t_R FILLER_22_1199 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_22_1207 ();
 DECAPx6_ASAP7_75t_R FILLER_22_1213 ();
 FILLER_ASAP7_75t_R FILLER_22_1230 ();
 DECAPx2_ASAP7_75t_R FILLER_22_1240 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_22_1246 ();
 FILLER_ASAP7_75t_R FILLER_22_1275 ();
 FILLER_ASAP7_75t_R FILLER_22_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_22_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_23_2 ();
 DECAPx10_ASAP7_75t_R FILLER_23_24 ();
 DECAPx10_ASAP7_75t_R FILLER_23_46 ();
 DECAPx10_ASAP7_75t_R FILLER_23_68 ();
 DECAPx10_ASAP7_75t_R FILLER_23_90 ();
 DECAPx10_ASAP7_75t_R FILLER_23_112 ();
 DECAPx10_ASAP7_75t_R FILLER_23_134 ();
 DECAPx10_ASAP7_75t_R FILLER_23_156 ();
 DECAPx10_ASAP7_75t_R FILLER_23_178 ();
 DECAPx10_ASAP7_75t_R FILLER_23_200 ();
 DECAPx10_ASAP7_75t_R FILLER_23_222 ();
 DECAPx10_ASAP7_75t_R FILLER_23_244 ();
 DECAPx10_ASAP7_75t_R FILLER_23_266 ();
 DECAPx10_ASAP7_75t_R FILLER_23_288 ();
 DECAPx10_ASAP7_75t_R FILLER_23_310 ();
 DECAPx10_ASAP7_75t_R FILLER_23_332 ();
 DECAPx10_ASAP7_75t_R FILLER_23_354 ();
 DECAPx10_ASAP7_75t_R FILLER_23_376 ();
 DECAPx10_ASAP7_75t_R FILLER_23_398 ();
 DECAPx2_ASAP7_75t_R FILLER_23_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_426 ();
 DECAPx6_ASAP7_75t_R FILLER_23_433 ();
 DECAPx2_ASAP7_75t_R FILLER_23_447 ();
 FILLER_ASAP7_75t_R FILLER_23_460 ();
 DECAPx2_ASAP7_75t_R FILLER_23_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_474 ();
 FILLER_ASAP7_75t_R FILLER_23_478 ();
 FILLER_ASAP7_75t_R FILLER_23_500 ();
 DECAPx4_ASAP7_75t_R FILLER_23_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_518 ();
 DECAPx4_ASAP7_75t_R FILLER_23_525 ();
 DECAPx10_ASAP7_75t_R FILLER_23_547 ();
 DECAPx2_ASAP7_75t_R FILLER_23_569 ();
 FILLER_ASAP7_75t_R FILLER_23_575 ();
 FILLER_ASAP7_75t_R FILLER_23_580 ();
 FILLER_ASAP7_75t_R FILLER_23_602 ();
 FILLER_ASAP7_75t_R FILLER_23_624 ();
 DECAPx6_ASAP7_75t_R FILLER_23_638 ();
 DECAPx1_ASAP7_75t_R FILLER_23_652 ();
 DECAPx4_ASAP7_75t_R FILLER_23_662 ();
 FILLER_ASAP7_75t_R FILLER_23_672 ();
 DECAPx2_ASAP7_75t_R FILLER_23_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_688 ();
 DECAPx6_ASAP7_75t_R FILLER_23_696 ();
 DECAPx10_ASAP7_75t_R FILLER_23_716 ();
 DECAPx6_ASAP7_75t_R FILLER_23_738 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_23_752 ();
 FILLER_ASAP7_75t_R FILLER_23_761 ();
 DECAPx2_ASAP7_75t_R FILLER_23_783 ();
 FILLER_ASAP7_75t_R FILLER_23_789 ();
 FILLER_ASAP7_75t_R FILLER_23_805 ();
 DECAPx1_ASAP7_75t_R FILLER_23_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_819 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_23_846 ();
 FILLER_ASAP7_75t_R FILLER_23_855 ();
 DECAPx1_ASAP7_75t_R FILLER_23_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_869 ();
 FILLER_ASAP7_75t_R FILLER_23_876 ();
 FILLER_ASAP7_75t_R FILLER_23_887 ();
 DECAPx6_ASAP7_75t_R FILLER_23_909 ();
 FILLER_ASAP7_75t_R FILLER_23_923 ();
 FILLER_ASAP7_75t_R FILLER_23_927 ();
 DECAPx6_ASAP7_75t_R FILLER_23_937 ();
 FILLER_ASAP7_75t_R FILLER_23_951 ();
 DECAPx2_ASAP7_75t_R FILLER_23_973 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_23_979 ();
 DECAPx6_ASAP7_75t_R FILLER_23_989 ();
 FILLER_ASAP7_75t_R FILLER_23_1003 ();
 DECAPx6_ASAP7_75t_R FILLER_23_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_23_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1038 ();
 FILLER_ASAP7_75t_R FILLER_23_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_23_1102 ();
 FILLER_ASAP7_75t_R FILLER_23_1128 ();
 FILLER_ASAP7_75t_R FILLER_23_1150 ();
 DECAPx4_ASAP7_75t_R FILLER_23_1178 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_23_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1217 ();
 DECAPx4_ASAP7_75t_R FILLER_23_1239 ();
 FILLER_ASAP7_75t_R FILLER_23_1256 ();
 FILLER_ASAP7_75t_R FILLER_23_1264 ();
 FILLER_ASAP7_75t_R FILLER_23_1292 ();
 FILLER_ASAP7_75t_R FILLER_23_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_23_1351 ();
 DECAPx1_ASAP7_75t_R FILLER_23_1373 ();
 DECAPx10_ASAP7_75t_R FILLER_24_2 ();
 DECAPx10_ASAP7_75t_R FILLER_24_24 ();
 DECAPx10_ASAP7_75t_R FILLER_24_46 ();
 DECAPx10_ASAP7_75t_R FILLER_24_68 ();
 DECAPx10_ASAP7_75t_R FILLER_24_90 ();
 DECAPx10_ASAP7_75t_R FILLER_24_112 ();
 DECAPx10_ASAP7_75t_R FILLER_24_134 ();
 DECAPx10_ASAP7_75t_R FILLER_24_156 ();
 DECAPx10_ASAP7_75t_R FILLER_24_178 ();
 DECAPx10_ASAP7_75t_R FILLER_24_200 ();
 DECAPx10_ASAP7_75t_R FILLER_24_222 ();
 DECAPx10_ASAP7_75t_R FILLER_24_244 ();
 DECAPx10_ASAP7_75t_R FILLER_24_266 ();
 DECAPx10_ASAP7_75t_R FILLER_24_288 ();
 DECAPx10_ASAP7_75t_R FILLER_24_310 ();
 DECAPx10_ASAP7_75t_R FILLER_24_332 ();
 DECAPx10_ASAP7_75t_R FILLER_24_354 ();
 DECAPx10_ASAP7_75t_R FILLER_24_376 ();
 DECAPx10_ASAP7_75t_R FILLER_24_398 ();
 DECAPx1_ASAP7_75t_R FILLER_24_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_424 ();
 DECAPx2_ASAP7_75t_R FILLER_24_432 ();
 DECAPx1_ASAP7_75t_R FILLER_24_458 ();
 FILLER_ASAP7_75t_R FILLER_24_464 ();
 DECAPx2_ASAP7_75t_R FILLER_24_473 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_485 ();
 DECAPx6_ASAP7_75t_R FILLER_24_496 ();
 DECAPx2_ASAP7_75t_R FILLER_24_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_516 ();
 FILLER_ASAP7_75t_R FILLER_24_524 ();
 DECAPx1_ASAP7_75t_R FILLER_24_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_536 ();
 DECAPx1_ASAP7_75t_R FILLER_24_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_561 ();
 DECAPx4_ASAP7_75t_R FILLER_24_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_575 ();
 FILLER_ASAP7_75t_R FILLER_24_582 ();
 DECAPx2_ASAP7_75t_R FILLER_24_587 ();
 DECAPx10_ASAP7_75t_R FILLER_24_599 ();
 DECAPx2_ASAP7_75t_R FILLER_24_621 ();
 FILLER_ASAP7_75t_R FILLER_24_647 ();
 DECAPx1_ASAP7_75t_R FILLER_24_652 ();
 DECAPx2_ASAP7_75t_R FILLER_24_663 ();
 FILLER_ASAP7_75t_R FILLER_24_669 ();
 FILLER_ASAP7_75t_R FILLER_24_691 ();
 DECAPx2_ASAP7_75t_R FILLER_24_701 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_707 ();
 FILLER_ASAP7_75t_R FILLER_24_720 ();
 DECAPx2_ASAP7_75t_R FILLER_24_730 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_736 ();
 DECAPx6_ASAP7_75t_R FILLER_24_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_763 ();
 DECAPx2_ASAP7_75t_R FILLER_24_772 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_778 ();
 DECAPx1_ASAP7_75t_R FILLER_24_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_794 ();
 DECAPx4_ASAP7_75t_R FILLER_24_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_815 ();
 FILLER_ASAP7_75t_R FILLER_24_822 ();
 DECAPx2_ASAP7_75t_R FILLER_24_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_833 ();
 DECAPx6_ASAP7_75t_R FILLER_24_837 ();
 DECAPx1_ASAP7_75t_R FILLER_24_851 ();
 DECAPx4_ASAP7_75t_R FILLER_24_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_885 ();
 FILLER_ASAP7_75t_R FILLER_24_892 ();
 DECAPx1_ASAP7_75t_R FILLER_24_897 ();
 FILLER_ASAP7_75t_R FILLER_24_907 ();
 FILLER_ASAP7_75t_R FILLER_24_916 ();
 FILLER_ASAP7_75t_R FILLER_24_924 ();
 FILLER_ASAP7_75t_R FILLER_24_946 ();
 DECAPx2_ASAP7_75t_R FILLER_24_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_960 ();
 FILLER_ASAP7_75t_R FILLER_24_987 ();
 FILLER_ASAP7_75t_R FILLER_24_997 ();
 FILLER_ASAP7_75t_R FILLER_24_1005 ();
 DECAPx1_ASAP7_75t_R FILLER_24_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_24_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1060 ();
 FILLER_ASAP7_75t_R FILLER_24_1082 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_1090 ();
 FILLER_ASAP7_75t_R FILLER_24_1099 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_24_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1122 ();
 FILLER_ASAP7_75t_R FILLER_24_1129 ();
 FILLER_ASAP7_75t_R FILLER_24_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_24_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_24_1158 ();
 FILLER_ASAP7_75t_R FILLER_24_1168 ();
 DECAPx4_ASAP7_75t_R FILLER_24_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1190 ();
 DECAPx4_ASAP7_75t_R FILLER_24_1199 ();
 FILLER_ASAP7_75t_R FILLER_24_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_24_1219 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_1225 ();
 FILLER_ASAP7_75t_R FILLER_24_1234 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_1242 ();
 DECAPx2_ASAP7_75t_R FILLER_24_1255 ();
 FILLER_ASAP7_75t_R FILLER_24_1261 ();
 FILLER_ASAP7_75t_R FILLER_24_1266 ();
 DECAPx2_ASAP7_75t_R FILLER_24_1276 ();
 FILLER_ASAP7_75t_R FILLER_24_1282 ();
 FILLER_ASAP7_75t_R FILLER_24_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_24_1340 ();
 DECAPx6_ASAP7_75t_R FILLER_24_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_25_2 ();
 DECAPx10_ASAP7_75t_R FILLER_25_24 ();
 DECAPx10_ASAP7_75t_R FILLER_25_46 ();
 DECAPx10_ASAP7_75t_R FILLER_25_68 ();
 DECAPx10_ASAP7_75t_R FILLER_25_90 ();
 DECAPx10_ASAP7_75t_R FILLER_25_112 ();
 DECAPx10_ASAP7_75t_R FILLER_25_134 ();
 DECAPx10_ASAP7_75t_R FILLER_25_156 ();
 DECAPx10_ASAP7_75t_R FILLER_25_178 ();
 DECAPx10_ASAP7_75t_R FILLER_25_200 ();
 DECAPx10_ASAP7_75t_R FILLER_25_222 ();
 DECAPx10_ASAP7_75t_R FILLER_25_244 ();
 DECAPx10_ASAP7_75t_R FILLER_25_266 ();
 DECAPx10_ASAP7_75t_R FILLER_25_288 ();
 DECAPx10_ASAP7_75t_R FILLER_25_310 ();
 DECAPx10_ASAP7_75t_R FILLER_25_332 ();
 DECAPx10_ASAP7_75t_R FILLER_25_354 ();
 DECAPx10_ASAP7_75t_R FILLER_25_376 ();
 DECAPx6_ASAP7_75t_R FILLER_25_398 ();
 DECAPx2_ASAP7_75t_R FILLER_25_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_418 ();
 FILLER_ASAP7_75t_R FILLER_25_439 ();
 DECAPx2_ASAP7_75t_R FILLER_25_448 ();
 DECAPx1_ASAP7_75t_R FILLER_25_460 ();
 DECAPx10_ASAP7_75t_R FILLER_25_470 ();
 DECAPx10_ASAP7_75t_R FILLER_25_492 ();
 FILLER_ASAP7_75t_R FILLER_25_514 ();
 FILLER_ASAP7_75t_R FILLER_25_524 ();
 DECAPx6_ASAP7_75t_R FILLER_25_532 ();
 FILLER_ASAP7_75t_R FILLER_25_546 ();
 DECAPx2_ASAP7_75t_R FILLER_25_551 ();
 DECAPx10_ASAP7_75t_R FILLER_25_569 ();
 DECAPx10_ASAP7_75t_R FILLER_25_591 ();
 DECAPx10_ASAP7_75t_R FILLER_25_613 ();
 DECAPx6_ASAP7_75t_R FILLER_25_635 ();
 DECAPx2_ASAP7_75t_R FILLER_25_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_655 ();
 DECAPx10_ASAP7_75t_R FILLER_25_662 ();
 FILLER_ASAP7_75t_R FILLER_25_684 ();
 DECAPx6_ASAP7_75t_R FILLER_25_689 ();
 FILLER_ASAP7_75t_R FILLER_25_703 ();
 FILLER_ASAP7_75t_R FILLER_25_711 ();
 FILLER_ASAP7_75t_R FILLER_25_733 ();
 FILLER_ASAP7_75t_R FILLER_25_747 ();
 DECAPx2_ASAP7_75t_R FILLER_25_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_762 ();
 DECAPx6_ASAP7_75t_R FILLER_25_770 ();
 DECAPx2_ASAP7_75t_R FILLER_25_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_790 ();
 FILLER_ASAP7_75t_R FILLER_25_795 ();
 DECAPx1_ASAP7_75t_R FILLER_25_807 ();
 FILLER_ASAP7_75t_R FILLER_25_817 ();
 DECAPx1_ASAP7_75t_R FILLER_25_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_831 ();
 DECAPx10_ASAP7_75t_R FILLER_25_835 ();
 DECAPx10_ASAP7_75t_R FILLER_25_857 ();
 DECAPx10_ASAP7_75t_R FILLER_25_879 ();
 DECAPx10_ASAP7_75t_R FILLER_25_901 ();
 FILLER_ASAP7_75t_R FILLER_25_923 ();
 FILLER_ASAP7_75t_R FILLER_25_927 ();
 DECAPx4_ASAP7_75t_R FILLER_25_935 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_25_945 ();
 DECAPx10_ASAP7_75t_R FILLER_25_954 ();
 DECAPx2_ASAP7_75t_R FILLER_25_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_985 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_25_992 ();
 FILLER_ASAP7_75t_R FILLER_25_1021 ();
 FILLER_ASAP7_75t_R FILLER_25_1029 ();
 DECAPx4_ASAP7_75t_R FILLER_25_1038 ();
 FILLER_ASAP7_75t_R FILLER_25_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_25_1169 ();
 FILLER_ASAP7_75t_R FILLER_25_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1184 ();
 DECAPx1_ASAP7_75t_R FILLER_25_1206 ();
 DECAPx6_ASAP7_75t_R FILLER_25_1230 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_25_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1253 ();
 DECAPx4_ASAP7_75t_R FILLER_25_1275 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_25_1285 ();
 FILLER_ASAP7_75t_R FILLER_25_1294 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_25_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_25_1335 ();
 DECAPx6_ASAP7_75t_R FILLER_25_1357 ();
 DECAPx2_ASAP7_75t_R FILLER_25_1371 ();
 DECAPx10_ASAP7_75t_R FILLER_26_2 ();
 DECAPx10_ASAP7_75t_R FILLER_26_24 ();
 DECAPx10_ASAP7_75t_R FILLER_26_46 ();
 DECAPx10_ASAP7_75t_R FILLER_26_68 ();
 DECAPx10_ASAP7_75t_R FILLER_26_90 ();
 DECAPx10_ASAP7_75t_R FILLER_26_112 ();
 DECAPx10_ASAP7_75t_R FILLER_26_134 ();
 DECAPx10_ASAP7_75t_R FILLER_26_156 ();
 DECAPx10_ASAP7_75t_R FILLER_26_178 ();
 DECAPx4_ASAP7_75t_R FILLER_26_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_210 ();
 DECAPx10_ASAP7_75t_R FILLER_26_237 ();
 DECAPx10_ASAP7_75t_R FILLER_26_259 ();
 DECAPx10_ASAP7_75t_R FILLER_26_281 ();
 DECAPx10_ASAP7_75t_R FILLER_26_303 ();
 DECAPx10_ASAP7_75t_R FILLER_26_325 ();
 DECAPx10_ASAP7_75t_R FILLER_26_347 ();
 DECAPx10_ASAP7_75t_R FILLER_26_369 ();
 DECAPx10_ASAP7_75t_R FILLER_26_391 ();
 DECAPx10_ASAP7_75t_R FILLER_26_413 ();
 DECAPx1_ASAP7_75t_R FILLER_26_441 ();
 DECAPx4_ASAP7_75t_R FILLER_26_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_461 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_26_464 ();
 DECAPx4_ASAP7_75t_R FILLER_26_475 ();
 DECAPx1_ASAP7_75t_R FILLER_26_497 ();
 DECAPx4_ASAP7_75t_R FILLER_26_504 ();
 DECAPx10_ASAP7_75t_R FILLER_26_534 ();
 DECAPx1_ASAP7_75t_R FILLER_26_576 ();
 DECAPx2_ASAP7_75t_R FILLER_26_586 ();
 FILLER_ASAP7_75t_R FILLER_26_592 ();
 DECAPx4_ASAP7_75t_R FILLER_26_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_612 ();
 FILLER_ASAP7_75t_R FILLER_26_619 ();
 DECAPx4_ASAP7_75t_R FILLER_26_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_639 ();
 DECAPx4_ASAP7_75t_R FILLER_26_646 ();
 DECAPx10_ASAP7_75t_R FILLER_26_664 ();
 DECAPx2_ASAP7_75t_R FILLER_26_698 ();
 DECAPx2_ASAP7_75t_R FILLER_26_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_713 ();
 DECAPx6_ASAP7_75t_R FILLER_26_717 ();
 DECAPx2_ASAP7_75t_R FILLER_26_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_737 ();
 FILLER_ASAP7_75t_R FILLER_26_745 ();
 DECAPx4_ASAP7_75t_R FILLER_26_754 ();
 FILLER_ASAP7_75t_R FILLER_26_764 ();
 FILLER_ASAP7_75t_R FILLER_26_774 ();
 DECAPx10_ASAP7_75t_R FILLER_26_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_804 ();
 DECAPx2_ASAP7_75t_R FILLER_26_811 ();
 FILLER_ASAP7_75t_R FILLER_26_843 ();
 DECAPx4_ASAP7_75t_R FILLER_26_853 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_26_863 ();
 DECAPx2_ASAP7_75t_R FILLER_26_872 ();
 FILLER_ASAP7_75t_R FILLER_26_878 ();
 FILLER_ASAP7_75t_R FILLER_26_886 ();
 DECAPx6_ASAP7_75t_R FILLER_26_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_910 ();
 FILLER_ASAP7_75t_R FILLER_26_917 ();
 DECAPx6_ASAP7_75t_R FILLER_26_925 ();
 DECAPx2_ASAP7_75t_R FILLER_26_939 ();
 FILLER_ASAP7_75t_R FILLER_26_953 ();
 DECAPx10_ASAP7_75t_R FILLER_26_958 ();
 DECAPx4_ASAP7_75t_R FILLER_26_980 ();
 FILLER_ASAP7_75t_R FILLER_26_990 ();
 DECAPx4_ASAP7_75t_R FILLER_26_999 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1012 ();
 DECAPx4_ASAP7_75t_R FILLER_26_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1044 ();
 FILLER_ASAP7_75t_R FILLER_26_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1093 ();
 FILLER_ASAP7_75t_R FILLER_26_1115 ();
 FILLER_ASAP7_75t_R FILLER_26_1126 ();
 DECAPx6_ASAP7_75t_R FILLER_26_1131 ();
 DECAPx1_ASAP7_75t_R FILLER_26_1152 ();
 DECAPx1_ASAP7_75t_R FILLER_26_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1169 ();
 FILLER_ASAP7_75t_R FILLER_26_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1204 ();
 DECAPx6_ASAP7_75t_R FILLER_26_1226 ();
 DECAPx2_ASAP7_75t_R FILLER_26_1240 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_26_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_26_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1279 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1301 ();
 FILLER_ASAP7_75t_R FILLER_26_1308 ();
 DECAPx2_ASAP7_75t_R FILLER_26_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_26_1349 ();
 DECAPx2_ASAP7_75t_R FILLER_26_1371 ();
 DECAPx10_ASAP7_75t_R FILLER_27_2 ();
 DECAPx10_ASAP7_75t_R FILLER_27_24 ();
 DECAPx10_ASAP7_75t_R FILLER_27_46 ();
 DECAPx6_ASAP7_75t_R FILLER_27_68 ();
 FILLER_ASAP7_75t_R FILLER_27_82 ();
 FILLER_ASAP7_75t_R FILLER_27_90 ();
 DECAPx4_ASAP7_75t_R FILLER_27_95 ();
 FILLER_ASAP7_75t_R FILLER_27_105 ();
 DECAPx10_ASAP7_75t_R FILLER_27_113 ();
 DECAPx10_ASAP7_75t_R FILLER_27_135 ();
 DECAPx10_ASAP7_75t_R FILLER_27_157 ();
 DECAPx10_ASAP7_75t_R FILLER_27_179 ();
 DECAPx10_ASAP7_75t_R FILLER_27_201 ();
 FILLER_ASAP7_75t_R FILLER_27_223 ();
 DECAPx1_ASAP7_75t_R FILLER_27_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_232 ();
 DECAPx2_ASAP7_75t_R FILLER_27_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_265 ();
 DECAPx10_ASAP7_75t_R FILLER_27_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_294 ();
 DECAPx10_ASAP7_75t_R FILLER_27_301 ();
 FILLER_ASAP7_75t_R FILLER_27_323 ();
 FILLER_ASAP7_75t_R FILLER_27_331 ();
 DECAPx10_ASAP7_75t_R FILLER_27_339 ();
 DECAPx2_ASAP7_75t_R FILLER_27_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_367 ();
 DECAPx10_ASAP7_75t_R FILLER_27_374 ();
 DECAPx10_ASAP7_75t_R FILLER_27_396 ();
 DECAPx10_ASAP7_75t_R FILLER_27_418 ();
 DECAPx2_ASAP7_75t_R FILLER_27_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_446 ();
 DECAPx4_ASAP7_75t_R FILLER_27_455 ();
 DECAPx1_ASAP7_75t_R FILLER_27_485 ();
 DECAPx10_ASAP7_75t_R FILLER_27_509 ();
 DECAPx1_ASAP7_75t_R FILLER_27_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_535 ();
 FILLER_ASAP7_75t_R FILLER_27_542 ();
 DECAPx6_ASAP7_75t_R FILLER_27_550 ();
 DECAPx1_ASAP7_75t_R FILLER_27_564 ();
 FILLER_ASAP7_75t_R FILLER_27_574 ();
 FILLER_ASAP7_75t_R FILLER_27_584 ();
 FILLER_ASAP7_75t_R FILLER_27_592 ();
 FILLER_ASAP7_75t_R FILLER_27_600 ();
 FILLER_ASAP7_75t_R FILLER_27_614 ();
 FILLER_ASAP7_75t_R FILLER_27_619 ();
 FILLER_ASAP7_75t_R FILLER_27_627 ();
 DECAPx2_ASAP7_75t_R FILLER_27_635 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_27_649 ();
 DECAPx6_ASAP7_75t_R FILLER_27_672 ();
 DECAPx1_ASAP7_75t_R FILLER_27_686 ();
 DECAPx1_ASAP7_75t_R FILLER_27_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_714 ();
 DECAPx6_ASAP7_75t_R FILLER_27_730 ();
 DECAPx2_ASAP7_75t_R FILLER_27_744 ();
 DECAPx4_ASAP7_75t_R FILLER_27_760 ();
 FILLER_ASAP7_75t_R FILLER_27_796 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_27_804 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_27_815 ();
 DECAPx6_ASAP7_75t_R FILLER_27_824 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_27_838 ();
 FILLER_ASAP7_75t_R FILLER_27_861 ();
 DECAPx4_ASAP7_75t_R FILLER_27_869 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_27_879 ();
 DECAPx2_ASAP7_75t_R FILLER_27_894 ();
 FILLER_ASAP7_75t_R FILLER_27_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_27_922 ();
 DECAPx2_ASAP7_75t_R FILLER_27_927 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_27_933 ();
 DECAPx1_ASAP7_75t_R FILLER_27_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_966 ();
 DECAPx2_ASAP7_75t_R FILLER_27_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_980 ();
 FILLER_ASAP7_75t_R FILLER_27_991 ();
 DECAPx2_ASAP7_75t_R FILLER_27_999 ();
 FILLER_ASAP7_75t_R FILLER_27_1005 ();
 DECAPx4_ASAP7_75t_R FILLER_27_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_1026 ();
 FILLER_ASAP7_75t_R FILLER_27_1030 ();
 FILLER_ASAP7_75t_R FILLER_27_1038 ();
 FILLER_ASAP7_75t_R FILLER_27_1046 ();
 DECAPx6_ASAP7_75t_R FILLER_27_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_27_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_27_1083 ();
 FILLER_ASAP7_75t_R FILLER_27_1097 ();
 FILLER_ASAP7_75t_R FILLER_27_1125 ();
 FILLER_ASAP7_75t_R FILLER_27_1153 ();
 DECAPx6_ASAP7_75t_R FILLER_27_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_27_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_1190 ();
 FILLER_ASAP7_75t_R FILLER_27_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_27_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_27_1209 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_27_1215 ();
 FILLER_ASAP7_75t_R FILLER_27_1227 ();
 DECAPx1_ASAP7_75t_R FILLER_27_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_1239 ();
 DECAPx1_ASAP7_75t_R FILLER_27_1250 ();
 FILLER_ASAP7_75t_R FILLER_27_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_27_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_28_2 ();
 DECAPx10_ASAP7_75t_R FILLER_28_24 ();
 DECAPx6_ASAP7_75t_R FILLER_28_46 ();
 FILLER_ASAP7_75t_R FILLER_28_60 ();
 FILLER_ASAP7_75t_R FILLER_28_68 ();
 FILLER_ASAP7_75t_R FILLER_28_96 ();
 DECAPx10_ASAP7_75t_R FILLER_28_124 ();
 DECAPx10_ASAP7_75t_R FILLER_28_146 ();
 DECAPx10_ASAP7_75t_R FILLER_28_174 ();
 DECAPx2_ASAP7_75t_R FILLER_28_196 ();
 FILLER_ASAP7_75t_R FILLER_28_202 ();
 DECAPx2_ASAP7_75t_R FILLER_28_210 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_222 ();
 DECAPx2_ASAP7_75t_R FILLER_28_231 ();
 FILLER_ASAP7_75t_R FILLER_28_243 ();
 DECAPx1_ASAP7_75t_R FILLER_28_251 ();
 DECAPx2_ASAP7_75t_R FILLER_28_281 ();
 FILLER_ASAP7_75t_R FILLER_28_287 ();
 DECAPx1_ASAP7_75t_R FILLER_28_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_319 ();
 DECAPx1_ASAP7_75t_R FILLER_28_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_350 ();
 FILLER_ASAP7_75t_R FILLER_28_357 ();
 FILLER_ASAP7_75t_R FILLER_28_362 ();
 DECAPx1_ASAP7_75t_R FILLER_28_390 ();
 FILLER_ASAP7_75t_R FILLER_28_397 ();
 DECAPx2_ASAP7_75t_R FILLER_28_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_431 ();
 FILLER_ASAP7_75t_R FILLER_28_438 ();
 FILLER_ASAP7_75t_R FILLER_28_460 ();
 DECAPx6_ASAP7_75t_R FILLER_28_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_478 ();
 FILLER_ASAP7_75t_R FILLER_28_487 ();
 DECAPx4_ASAP7_75t_R FILLER_28_492 ();
 DECAPx6_ASAP7_75t_R FILLER_28_508 ();
 DECAPx2_ASAP7_75t_R FILLER_28_522 ();
 FILLER_ASAP7_75t_R FILLER_28_534 ();
 DECAPx2_ASAP7_75t_R FILLER_28_544 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_550 ();
 DECAPx6_ASAP7_75t_R FILLER_28_559 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_576 ();
 DECAPx6_ASAP7_75t_R FILLER_28_585 ();
 DECAPx1_ASAP7_75t_R FILLER_28_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_603 ();
 DECAPx6_ASAP7_75t_R FILLER_28_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_638 ();
 DECAPx6_ASAP7_75t_R FILLER_28_645 ();
 DECAPx2_ASAP7_75t_R FILLER_28_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_665 ();
 FILLER_ASAP7_75t_R FILLER_28_669 ();
 DECAPx1_ASAP7_75t_R FILLER_28_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_687 ();
 DECAPx6_ASAP7_75t_R FILLER_28_691 ();
 DECAPx1_ASAP7_75t_R FILLER_28_705 ();
 FILLER_ASAP7_75t_R FILLER_28_721 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_729 ();
 DECAPx10_ASAP7_75t_R FILLER_28_744 ();
 FILLER_ASAP7_75t_R FILLER_28_773 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_782 ();
 DECAPx6_ASAP7_75t_R FILLER_28_823 ();
 FILLER_ASAP7_75t_R FILLER_28_849 ();
 DECAPx1_ASAP7_75t_R FILLER_28_858 ();
 FILLER_ASAP7_75t_R FILLER_28_868 ();
 DECAPx2_ASAP7_75t_R FILLER_28_877 ();
 FILLER_ASAP7_75t_R FILLER_28_883 ();
 DECAPx6_ASAP7_75t_R FILLER_28_905 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_919 ();
 DECAPx6_ASAP7_75t_R FILLER_28_931 ();
 DECAPx1_ASAP7_75t_R FILLER_28_951 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_965 ();
 DECAPx4_ASAP7_75t_R FILLER_28_994 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_1004 ();
 FILLER_ASAP7_75t_R FILLER_28_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1060 ();
 DECAPx1_ASAP7_75t_R FILLER_28_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1074 ();
 FILLER_ASAP7_75t_R FILLER_28_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_28_1086 ();
 FILLER_ASAP7_75t_R FILLER_28_1098 ();
 FILLER_ASAP7_75t_R FILLER_28_1107 ();
 FILLER_ASAP7_75t_R FILLER_28_1115 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_28_1132 ();
 FILLER_ASAP7_75t_R FILLER_28_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_28_1143 ();
 FILLER_ASAP7_75t_R FILLER_28_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_28_1157 ();
 FILLER_ASAP7_75t_R FILLER_28_1163 ();
 DECAPx4_ASAP7_75t_R FILLER_28_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_1181 ();
 DECAPx2_ASAP7_75t_R FILLER_28_1185 ();
 FILLER_ASAP7_75t_R FILLER_28_1191 ();
 FILLER_ASAP7_75t_R FILLER_28_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_28_1247 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_1253 ();
 FILLER_ASAP7_75t_R FILLER_28_1262 ();
 FILLER_ASAP7_75t_R FILLER_28_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_28_1318 ();
 DECAPx4_ASAP7_75t_R FILLER_28_1340 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_1350 ();
 FILLER_ASAP7_75t_R FILLER_28_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_29_2 ();
 DECAPx4_ASAP7_75t_R FILLER_29_24 ();
 FILLER_ASAP7_75t_R FILLER_29_34 ();
 FILLER_ASAP7_75t_R FILLER_29_42 ();
 FILLER_ASAP7_75t_R FILLER_29_70 ();
 DECAPx1_ASAP7_75t_R FILLER_29_75 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_85 ();
 DECAPx4_ASAP7_75t_R FILLER_29_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_101 ();
 DECAPx1_ASAP7_75t_R FILLER_29_108 ();
 DECAPx4_ASAP7_75t_R FILLER_29_115 ();
 FILLER_ASAP7_75t_R FILLER_29_125 ();
 DECAPx1_ASAP7_75t_R FILLER_29_153 ();
 DECAPx4_ASAP7_75t_R FILLER_29_183 ();
 FILLER_ASAP7_75t_R FILLER_29_193 ();
 DECAPx4_ASAP7_75t_R FILLER_29_221 ();
 DECAPx4_ASAP7_75t_R FILLER_29_234 ();
 FILLER_ASAP7_75t_R FILLER_29_244 ();
 FILLER_ASAP7_75t_R FILLER_29_249 ();
 DECAPx2_ASAP7_75t_R FILLER_29_254 ();
 FILLER_ASAP7_75t_R FILLER_29_266 ();
 FILLER_ASAP7_75t_R FILLER_29_271 ();
 DECAPx4_ASAP7_75t_R FILLER_29_276 ();
 DECAPx2_ASAP7_75t_R FILLER_29_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_298 ();
 FILLER_ASAP7_75t_R FILLER_29_302 ();
 DECAPx1_ASAP7_75t_R FILLER_29_310 ();
 DECAPx2_ASAP7_75t_R FILLER_29_320 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_332 ();
 FILLER_ASAP7_75t_R FILLER_29_338 ();
 DECAPx1_ASAP7_75t_R FILLER_29_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_370 ();
 FILLER_ASAP7_75t_R FILLER_29_377 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_382 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_411 ();
 FILLER_ASAP7_75t_R FILLER_29_417 ();
 DECAPx6_ASAP7_75t_R FILLER_29_445 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_459 ();
 DECAPx10_ASAP7_75t_R FILLER_29_465 ();
 FILLER_ASAP7_75t_R FILLER_29_487 ();
 DECAPx10_ASAP7_75t_R FILLER_29_492 ();
 DECAPx2_ASAP7_75t_R FILLER_29_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_520 ();
 FILLER_ASAP7_75t_R FILLER_29_524 ();
 DECAPx4_ASAP7_75t_R FILLER_29_529 ();
 FILLER_ASAP7_75t_R FILLER_29_539 ();
 DECAPx1_ASAP7_75t_R FILLER_29_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_551 ();
 DECAPx10_ASAP7_75t_R FILLER_29_558 ();
 DECAPx10_ASAP7_75t_R FILLER_29_580 ();
 DECAPx1_ASAP7_75t_R FILLER_29_602 ();
 DECAPx4_ASAP7_75t_R FILLER_29_609 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_619 ();
 FILLER_ASAP7_75t_R FILLER_29_628 ();
 DECAPx6_ASAP7_75t_R FILLER_29_638 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_652 ();
 DECAPx4_ASAP7_75t_R FILLER_29_661 ();
 FILLER_ASAP7_75t_R FILLER_29_674 ();
 DECAPx6_ASAP7_75t_R FILLER_29_696 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_710 ();
 DECAPx2_ASAP7_75t_R FILLER_29_733 ();
 FILLER_ASAP7_75t_R FILLER_29_753 ();
 FILLER_ASAP7_75t_R FILLER_29_761 ();
 DECAPx6_ASAP7_75t_R FILLER_29_769 ();
 FILLER_ASAP7_75t_R FILLER_29_783 ();
 DECAPx2_ASAP7_75t_R FILLER_29_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_794 ();
 DECAPx1_ASAP7_75t_R FILLER_29_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_807 ();
 FILLER_ASAP7_75t_R FILLER_29_834 ();
 DECAPx4_ASAP7_75t_R FILLER_29_842 ();
 FILLER_ASAP7_75t_R FILLER_29_864 ();
 DECAPx10_ASAP7_75t_R FILLER_29_874 ();
 DECAPx10_ASAP7_75t_R FILLER_29_896 ();
 FILLER_ASAP7_75t_R FILLER_29_918 ();
 FILLER_ASAP7_75t_R FILLER_29_923 ();
 FILLER_ASAP7_75t_R FILLER_29_927 ();
 DECAPx2_ASAP7_75t_R FILLER_29_955 ();
 FILLER_ASAP7_75t_R FILLER_29_961 ();
 FILLER_ASAP7_75t_R FILLER_29_969 ();
 DECAPx2_ASAP7_75t_R FILLER_29_977 ();
 DECAPx10_ASAP7_75t_R FILLER_29_986 ();
 DECAPx1_ASAP7_75t_R FILLER_29_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1018 ();
 DECAPx4_ASAP7_75t_R FILLER_29_1040 ();
 FILLER_ASAP7_75t_R FILLER_29_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_29_1058 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_29_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1082 ();
 DECAPx4_ASAP7_75t_R FILLER_29_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_29_1117 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1132 ();
 DECAPx2_ASAP7_75t_R FILLER_29_1154 ();
 FILLER_ASAP7_75t_R FILLER_29_1160 ();
 FILLER_ASAP7_75t_R FILLER_29_1165 ();
 DECAPx6_ASAP7_75t_R FILLER_29_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1211 ();
 FILLER_ASAP7_75t_R FILLER_29_1236 ();
 DECAPx1_ASAP7_75t_R FILLER_29_1241 ();
 FILLER_ASAP7_75t_R FILLER_29_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_29_1259 ();
 DECAPx2_ASAP7_75t_R FILLER_29_1273 ();
 DECAPx1_ASAP7_75t_R FILLER_29_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1286 ();
 FILLER_ASAP7_75t_R FILLER_29_1293 ();
 DECAPx1_ASAP7_75t_R FILLER_29_1303 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1307 ();
 FILLER_ASAP7_75t_R FILLER_29_1314 ();
 DECAPx2_ASAP7_75t_R FILLER_29_1323 ();
 FILLER_ASAP7_75t_R FILLER_29_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_29_1334 ();
 DECAPx6_ASAP7_75t_R FILLER_29_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_29_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_30_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_24 ();
 FILLER_ASAP7_75t_R FILLER_30_53 ();
 FILLER_ASAP7_75t_R FILLER_30_62 ();
 FILLER_ASAP7_75t_R FILLER_30_70 ();
 FILLER_ASAP7_75t_R FILLER_30_75 ();
 DECAPx10_ASAP7_75t_R FILLER_30_80 ();
 DECAPx1_ASAP7_75t_R FILLER_30_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_106 ();
 FILLER_ASAP7_75t_R FILLER_30_110 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_118 ();
 DECAPx2_ASAP7_75t_R FILLER_30_124 ();
 FILLER_ASAP7_75t_R FILLER_30_130 ();
 FILLER_ASAP7_75t_R FILLER_30_138 ();
 FILLER_ASAP7_75t_R FILLER_30_146 ();
 FILLER_ASAP7_75t_R FILLER_30_151 ();
 DECAPx1_ASAP7_75t_R FILLER_30_159 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_169 ();
 DECAPx1_ASAP7_75t_R FILLER_30_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_179 ();
 FILLER_ASAP7_75t_R FILLER_30_186 ();
 DECAPx2_ASAP7_75t_R FILLER_30_194 ();
 DECAPx1_ASAP7_75t_R FILLER_30_206 ();
 DECAPx4_ASAP7_75t_R FILLER_30_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_223 ();
 DECAPx10_ASAP7_75t_R FILLER_30_227 ();
 DECAPx10_ASAP7_75t_R FILLER_30_249 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_271 ();
 DECAPx2_ASAP7_75t_R FILLER_30_300 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_306 ();
 DECAPx4_ASAP7_75t_R FILLER_30_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_345 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_352 ();
 DECAPx4_ASAP7_75t_R FILLER_30_358 ();
 FILLER_ASAP7_75t_R FILLER_30_368 ();
 DECAPx6_ASAP7_75t_R FILLER_30_373 ();
 FILLER_ASAP7_75t_R FILLER_30_387 ();
 FILLER_ASAP7_75t_R FILLER_30_395 ();
 FILLER_ASAP7_75t_R FILLER_30_403 ();
 FILLER_ASAP7_75t_R FILLER_30_411 ();
 DECAPx2_ASAP7_75t_R FILLER_30_419 ();
 FILLER_ASAP7_75t_R FILLER_30_431 ();
 FILLER_ASAP7_75t_R FILLER_30_436 ();
 DECAPx6_ASAP7_75t_R FILLER_30_441 ();
 DECAPx2_ASAP7_75t_R FILLER_30_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_461 ();
 FILLER_ASAP7_75t_R FILLER_30_464 ();
 DECAPx1_ASAP7_75t_R FILLER_30_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_482 ();
 DECAPx1_ASAP7_75t_R FILLER_30_490 ();
 FILLER_ASAP7_75t_R FILLER_30_500 ();
 DECAPx2_ASAP7_75t_R FILLER_30_510 ();
 DECAPx2_ASAP7_75t_R FILLER_30_528 ();
 DECAPx10_ASAP7_75t_R FILLER_30_540 ();
 DECAPx6_ASAP7_75t_R FILLER_30_562 ();
 DECAPx1_ASAP7_75t_R FILLER_30_576 ();
 FILLER_ASAP7_75t_R FILLER_30_588 ();
 DECAPx10_ASAP7_75t_R FILLER_30_597 ();
 DECAPx4_ASAP7_75t_R FILLER_30_619 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_629 ();
 FILLER_ASAP7_75t_R FILLER_30_640 ();
 DECAPx1_ASAP7_75t_R FILLER_30_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_653 ();
 DECAPx10_ASAP7_75t_R FILLER_30_661 ();
 DECAPx2_ASAP7_75t_R FILLER_30_683 ();
 FILLER_ASAP7_75t_R FILLER_30_711 ();
 FILLER_ASAP7_75t_R FILLER_30_719 ();
 DECAPx6_ASAP7_75t_R FILLER_30_724 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_738 ();
 FILLER_ASAP7_75t_R FILLER_30_757 ();
 DECAPx10_ASAP7_75t_R FILLER_30_767 ();
 FILLER_ASAP7_75t_R FILLER_30_789 ();
 DECAPx1_ASAP7_75t_R FILLER_30_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_821 ();
 DECAPx10_ASAP7_75t_R FILLER_30_825 ();
 DECAPx4_ASAP7_75t_R FILLER_30_847 ();
 FILLER_ASAP7_75t_R FILLER_30_857 ();
 DECAPx10_ASAP7_75t_R FILLER_30_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_901 ();
 FILLER_ASAP7_75t_R FILLER_30_908 ();
 FILLER_ASAP7_75t_R FILLER_30_916 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_924 ();
 DECAPx2_ASAP7_75t_R FILLER_30_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_939 ();
 DECAPx6_ASAP7_75t_R FILLER_30_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_957 ();
 DECAPx6_ASAP7_75t_R FILLER_30_968 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_982 ();
 FILLER_ASAP7_75t_R FILLER_30_991 ();
 FILLER_ASAP7_75t_R FILLER_30_1002 ();
 DECAPx6_ASAP7_75t_R FILLER_30_1010 ();
 DECAPx6_ASAP7_75t_R FILLER_30_1034 ();
 FILLER_ASAP7_75t_R FILLER_30_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_30_1056 ();
 FILLER_ASAP7_75t_R FILLER_30_1062 ();
 DECAPx2_ASAP7_75t_R FILLER_30_1090 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1102 ();
 DECAPx1_ASAP7_75t_R FILLER_30_1124 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1182 ();
 DECAPx6_ASAP7_75t_R FILLER_30_1204 ();
 FILLER_ASAP7_75t_R FILLER_30_1218 ();
 DECAPx1_ASAP7_75t_R FILLER_30_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1230 ();
 DECAPx6_ASAP7_75t_R FILLER_30_1241 ();
 FILLER_ASAP7_75t_R FILLER_30_1255 ();
 DECAPx4_ASAP7_75t_R FILLER_30_1263 ();
 DECAPx6_ASAP7_75t_R FILLER_30_1279 ();
 DECAPx2_ASAP7_75t_R FILLER_30_1293 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_1299 ();
 FILLER_ASAP7_75t_R FILLER_30_1310 ();
 FILLER_ASAP7_75t_R FILLER_30_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_30_1343 ();
 DECAPx4_ASAP7_75t_R FILLER_30_1365 ();
 FILLER_ASAP7_75t_R FILLER_30_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_31_2 ();
 DECAPx2_ASAP7_75t_R FILLER_31_24 ();
 DECAPx1_ASAP7_75t_R FILLER_31_36 ();
 FILLER_ASAP7_75t_R FILLER_31_47 ();
 FILLER_ASAP7_75t_R FILLER_31_56 ();
 FILLER_ASAP7_75t_R FILLER_31_65 ();
 FILLER_ASAP7_75t_R FILLER_31_74 ();
 DECAPx2_ASAP7_75t_R FILLER_31_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_88 ();
 DECAPx4_ASAP7_75t_R FILLER_31_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_105 ();
 DECAPx4_ASAP7_75t_R FILLER_31_132 ();
 FILLER_ASAP7_75t_R FILLER_31_142 ();
 DECAPx1_ASAP7_75t_R FILLER_31_170 ();
 DECAPx6_ASAP7_75t_R FILLER_31_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_214 ();
 FILLER_ASAP7_75t_R FILLER_31_221 ();
 DECAPx2_ASAP7_75t_R FILLER_31_226 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_232 ();
 DECAPx2_ASAP7_75t_R FILLER_31_261 ();
 DECAPx2_ASAP7_75t_R FILLER_31_273 ();
 FILLER_ASAP7_75t_R FILLER_31_279 ();
 FILLER_ASAP7_75t_R FILLER_31_287 ();
 DECAPx1_ASAP7_75t_R FILLER_31_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_296 ();
 DECAPx4_ASAP7_75t_R FILLER_31_300 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_310 ();
 DECAPx2_ASAP7_75t_R FILLER_31_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_322 ();
 DECAPx2_ASAP7_75t_R FILLER_31_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_332 ();
 DECAPx6_ASAP7_75t_R FILLER_31_336 ();
 DECAPx2_ASAP7_75t_R FILLER_31_350 ();
 DECAPx6_ASAP7_75t_R FILLER_31_362 ();
 DECAPx1_ASAP7_75t_R FILLER_31_376 ();
 DECAPx2_ASAP7_75t_R FILLER_31_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_392 ();
 DECAPx4_ASAP7_75t_R FILLER_31_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_409 ();
 DECAPx6_ASAP7_75t_R FILLER_31_413 ();
 DECAPx2_ASAP7_75t_R FILLER_31_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_433 ();
 DECAPx2_ASAP7_75t_R FILLER_31_440 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_446 ();
 FILLER_ASAP7_75t_R FILLER_31_475 ();
 FILLER_ASAP7_75t_R FILLER_31_497 ();
 FILLER_ASAP7_75t_R FILLER_31_505 ();
 DECAPx1_ASAP7_75t_R FILLER_31_514 ();
 FILLER_ASAP7_75t_R FILLER_31_538 ();
 DECAPx2_ASAP7_75t_R FILLER_31_548 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_554 ();
 FILLER_ASAP7_75t_R FILLER_31_563 ();
 DECAPx4_ASAP7_75t_R FILLER_31_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_581 ();
 FILLER_ASAP7_75t_R FILLER_31_588 ();
 FILLER_ASAP7_75t_R FILLER_31_596 ();
 DECAPx4_ASAP7_75t_R FILLER_31_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_618 ();
 DECAPx10_ASAP7_75t_R FILLER_31_633 ();
 FILLER_ASAP7_75t_R FILLER_31_655 ();
 DECAPx2_ASAP7_75t_R FILLER_31_663 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_669 ();
 FILLER_ASAP7_75t_R FILLER_31_680 ();
 DECAPx1_ASAP7_75t_R FILLER_31_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_692 ();
 DECAPx2_ASAP7_75t_R FILLER_31_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_705 ();
 FILLER_ASAP7_75t_R FILLER_31_713 ();
 DECAPx10_ASAP7_75t_R FILLER_31_721 ();
 DECAPx2_ASAP7_75t_R FILLER_31_743 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_749 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_772 ();
 DECAPx1_ASAP7_75t_R FILLER_31_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_805 ();
 DECAPx2_ASAP7_75t_R FILLER_31_809 ();
 FILLER_ASAP7_75t_R FILLER_31_815 ();
 FILLER_ASAP7_75t_R FILLER_31_825 ();
 FILLER_ASAP7_75t_R FILLER_31_833 ();
 DECAPx6_ASAP7_75t_R FILLER_31_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_852 ();
 DECAPx10_ASAP7_75t_R FILLER_31_859 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_881 ();
 FILLER_ASAP7_75t_R FILLER_31_891 ();
 FILLER_ASAP7_75t_R FILLER_31_899 ();
 DECAPx2_ASAP7_75t_R FILLER_31_907 ();
 DECAPx1_ASAP7_75t_R FILLER_31_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_924 ();
 DECAPx4_ASAP7_75t_R FILLER_31_927 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_937 ();
 DECAPx2_ASAP7_75t_R FILLER_31_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_953 ();
 FILLER_ASAP7_75t_R FILLER_31_960 ();
 DECAPx1_ASAP7_75t_R FILLER_31_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_992 ();
 DECAPx1_ASAP7_75t_R FILLER_31_1001 ();
 FILLER_ASAP7_75t_R FILLER_31_1031 ();
 FILLER_ASAP7_75t_R FILLER_31_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_31_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_31_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1076 ();
 FILLER_ASAP7_75t_R FILLER_31_1083 ();
 DECAPx4_ASAP7_75t_R FILLER_31_1111 ();
 FILLER_ASAP7_75t_R FILLER_31_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_31_1133 ();
 FILLER_ASAP7_75t_R FILLER_31_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_31_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_31_1183 ();
 FILLER_ASAP7_75t_R FILLER_31_1189 ();
 FILLER_ASAP7_75t_R FILLER_31_1217 ();
 DECAPx4_ASAP7_75t_R FILLER_31_1245 ();
 FILLER_ASAP7_75t_R FILLER_31_1255 ();
 DECAPx2_ASAP7_75t_R FILLER_31_1267 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_1273 ();
 DECAPx4_ASAP7_75t_R FILLER_31_1284 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_1294 ();
 DECAPx6_ASAP7_75t_R FILLER_31_1300 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_31_1345 ();
 DECAPx4_ASAP7_75t_R FILLER_31_1367 ();
 DECAPx6_ASAP7_75t_R FILLER_32_2 ();
 FILLER_ASAP7_75t_R FILLER_32_22 ();
 DECAPx4_ASAP7_75t_R FILLER_32_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_40 ();
 DECAPx2_ASAP7_75t_R FILLER_32_44 ();
 DECAPx1_ASAP7_75t_R FILLER_32_76 ();
 DECAPx1_ASAP7_75t_R FILLER_32_106 ();
 DECAPx10_ASAP7_75t_R FILLER_32_116 ();
 DECAPx4_ASAP7_75t_R FILLER_32_138 ();
 DECAPx1_ASAP7_75t_R FILLER_32_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_158 ();
 DECAPx10_ASAP7_75t_R FILLER_32_162 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_184 ();
 FILLER_ASAP7_75t_R FILLER_32_193 ();
 DECAPx4_ASAP7_75t_R FILLER_32_198 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_234 ();
 FILLER_ASAP7_75t_R FILLER_32_243 ();
 FILLER_ASAP7_75t_R FILLER_32_251 ();
 DECAPx1_ASAP7_75t_R FILLER_32_279 ();
 DECAPx10_ASAP7_75t_R FILLER_32_289 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_311 ();
 DECAPx6_ASAP7_75t_R FILLER_32_320 ();
 DECAPx2_ASAP7_75t_R FILLER_32_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_346 ();
 FILLER_ASAP7_75t_R FILLER_32_373 ();
 FILLER_ASAP7_75t_R FILLER_32_401 ();
 DECAPx2_ASAP7_75t_R FILLER_32_406 ();
 FILLER_ASAP7_75t_R FILLER_32_412 ();
 DECAPx1_ASAP7_75t_R FILLER_32_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_424 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_451 ();
 FILLER_ASAP7_75t_R FILLER_32_460 ();
 FILLER_ASAP7_75t_R FILLER_32_464 ();
 DECAPx4_ASAP7_75t_R FILLER_32_472 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_482 ();
 FILLER_ASAP7_75t_R FILLER_32_491 ();
 FILLER_ASAP7_75t_R FILLER_32_501 ();
 DECAPx10_ASAP7_75t_R FILLER_32_510 ();
 DECAPx6_ASAP7_75t_R FILLER_32_532 ();
 FILLER_ASAP7_75t_R FILLER_32_546 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_556 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_568 ();
 FILLER_ASAP7_75t_R FILLER_32_580 ();
 DECAPx2_ASAP7_75t_R FILLER_32_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_595 ();
 DECAPx2_ASAP7_75t_R FILLER_32_606 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_612 ();
 FILLER_ASAP7_75t_R FILLER_32_622 ();
 DECAPx2_ASAP7_75t_R FILLER_32_630 ();
 FILLER_ASAP7_75t_R FILLER_32_636 ();
 DECAPx2_ASAP7_75t_R FILLER_32_645 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_651 ();
 FILLER_ASAP7_75t_R FILLER_32_660 ();
 DECAPx10_ASAP7_75t_R FILLER_32_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_690 ();
 FILLER_ASAP7_75t_R FILLER_32_697 ();
 DECAPx4_ASAP7_75t_R FILLER_32_705 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_715 ();
 DECAPx1_ASAP7_75t_R FILLER_32_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_728 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_735 ();
 DECAPx6_ASAP7_75t_R FILLER_32_744 ();
 DECAPx2_ASAP7_75t_R FILLER_32_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_764 ();
 FILLER_ASAP7_75t_R FILLER_32_771 ();
 FILLER_ASAP7_75t_R FILLER_32_780 ();
 FILLER_ASAP7_75t_R FILLER_32_789 ();
 FILLER_ASAP7_75t_R FILLER_32_797 ();
 DECAPx4_ASAP7_75t_R FILLER_32_802 ();
 FILLER_ASAP7_75t_R FILLER_32_832 ();
 DECAPx1_ASAP7_75t_R FILLER_32_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_847 ();
 DECAPx4_ASAP7_75t_R FILLER_32_851 ();
 FILLER_ASAP7_75t_R FILLER_32_867 ();
 DECAPx2_ASAP7_75t_R FILLER_32_875 ();
 FILLER_ASAP7_75t_R FILLER_32_881 ();
 DECAPx1_ASAP7_75t_R FILLER_32_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_907 ();
 FILLER_ASAP7_75t_R FILLER_32_911 ();
 FILLER_ASAP7_75t_R FILLER_32_933 ();
 DECAPx6_ASAP7_75t_R FILLER_32_941 ();
 DECAPx1_ASAP7_75t_R FILLER_32_955 ();
 DECAPx6_ASAP7_75t_R FILLER_32_962 ();
 DECAPx10_ASAP7_75t_R FILLER_32_979 ();
 DECAPx2_ASAP7_75t_R FILLER_32_1001 ();
 DECAPx4_ASAP7_75t_R FILLER_32_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_32_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_32_1036 ();
 DECAPx2_ASAP7_75t_R FILLER_32_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_32_1067 ();
 FILLER_ASAP7_75t_R FILLER_32_1089 ();
 DECAPx4_ASAP7_75t_R FILLER_32_1101 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_1111 ();
 FILLER_ASAP7_75t_R FILLER_32_1122 ();
 DECAPx4_ASAP7_75t_R FILLER_32_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_32_1152 ();
 FILLER_ASAP7_75t_R FILLER_32_1166 ();
 FILLER_ASAP7_75t_R FILLER_32_1174 ();
 FILLER_ASAP7_75t_R FILLER_32_1202 ();
 FILLER_ASAP7_75t_R FILLER_32_1211 ();
 DECAPx4_ASAP7_75t_R FILLER_32_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_1229 ();
 FILLER_ASAP7_75t_R FILLER_32_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_32_1242 ();
 DECAPx1_ASAP7_75t_R FILLER_32_1256 ();
 FILLER_ASAP7_75t_R FILLER_32_1286 ();
 DECAPx4_ASAP7_75t_R FILLER_32_1314 ();
 FILLER_ASAP7_75t_R FILLER_32_1324 ();
 FILLER_ASAP7_75t_R FILLER_32_1333 ();
 FILLER_ASAP7_75t_R FILLER_32_1341 ();
 FILLER_ASAP7_75t_R FILLER_32_1346 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_1374 ();
 DECAPx2_ASAP7_75t_R FILLER_33_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_8 ();
 FILLER_ASAP7_75t_R FILLER_33_37 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_42 ();
 DECAPx6_ASAP7_75t_R FILLER_33_51 ();
 FILLER_ASAP7_75t_R FILLER_33_65 ();
 FILLER_ASAP7_75t_R FILLER_33_73 ();
 DECAPx1_ASAP7_75t_R FILLER_33_81 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_91 ();
 DECAPx4_ASAP7_75t_R FILLER_33_97 ();
 DECAPx6_ASAP7_75t_R FILLER_33_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_127 ();
 DECAPx1_ASAP7_75t_R FILLER_33_134 ();
 DECAPx10_ASAP7_75t_R FILLER_33_141 ();
 FILLER_ASAP7_75t_R FILLER_33_166 ();
 DECAPx2_ASAP7_75t_R FILLER_33_174 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_180 ();
 FILLER_ASAP7_75t_R FILLER_33_209 ();
 DECAPx4_ASAP7_75t_R FILLER_33_217 ();
 FILLER_ASAP7_75t_R FILLER_33_227 ();
 FILLER_ASAP7_75t_R FILLER_33_235 ();
 DECAPx2_ASAP7_75t_R FILLER_33_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_249 ();
 DECAPx2_ASAP7_75t_R FILLER_33_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_259 ();
 FILLER_ASAP7_75t_R FILLER_33_266 ();
 DECAPx2_ASAP7_75t_R FILLER_33_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_277 ();
 DECAPx1_ASAP7_75t_R FILLER_33_304 ();
 FILLER_ASAP7_75t_R FILLER_33_334 ();
 DECAPx4_ASAP7_75t_R FILLER_33_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_352 ();
 DECAPx1_ASAP7_75t_R FILLER_33_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_363 ();
 DECAPx4_ASAP7_75t_R FILLER_33_367 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_377 ();
 DECAPx1_ASAP7_75t_R FILLER_33_386 ();
 DECAPx2_ASAP7_75t_R FILLER_33_393 ();
 DECAPx2_ASAP7_75t_R FILLER_33_402 ();
 FILLER_ASAP7_75t_R FILLER_33_414 ();
 DECAPx2_ASAP7_75t_R FILLER_33_423 ();
 DECAPx1_ASAP7_75t_R FILLER_33_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_439 ();
 DECAPx6_ASAP7_75t_R FILLER_33_443 ();
 DECAPx2_ASAP7_75t_R FILLER_33_457 ();
 DECAPx10_ASAP7_75t_R FILLER_33_466 ();
 DECAPx10_ASAP7_75t_R FILLER_33_488 ();
 FILLER_ASAP7_75t_R FILLER_33_510 ();
 DECAPx2_ASAP7_75t_R FILLER_33_540 ();
 FILLER_ASAP7_75t_R FILLER_33_546 ();
 DECAPx2_ASAP7_75t_R FILLER_33_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_561 ();
 DECAPx2_ASAP7_75t_R FILLER_33_568 ();
 FILLER_ASAP7_75t_R FILLER_33_574 ();
 FILLER_ASAP7_75t_R FILLER_33_582 ();
 FILLER_ASAP7_75t_R FILLER_33_606 ();
 DECAPx2_ASAP7_75t_R FILLER_33_614 ();
 FILLER_ASAP7_75t_R FILLER_33_626 ();
 FILLER_ASAP7_75t_R FILLER_33_634 ();
 FILLER_ASAP7_75t_R FILLER_33_650 ();
 DECAPx1_ASAP7_75t_R FILLER_33_662 ();
 DECAPx6_ASAP7_75t_R FILLER_33_672 ();
 DECAPx1_ASAP7_75t_R FILLER_33_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_690 ();
 DECAPx6_ASAP7_75t_R FILLER_33_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_713 ();
 FILLER_ASAP7_75t_R FILLER_33_722 ();
 DECAPx2_ASAP7_75t_R FILLER_33_730 ();
 FILLER_ASAP7_75t_R FILLER_33_736 ();
 DECAPx10_ASAP7_75t_R FILLER_33_746 ();
 DECAPx10_ASAP7_75t_R FILLER_33_768 ();
 DECAPx10_ASAP7_75t_R FILLER_33_796 ();
 DECAPx4_ASAP7_75t_R FILLER_33_818 ();
 FILLER_ASAP7_75t_R FILLER_33_828 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_836 ();
 FILLER_ASAP7_75t_R FILLER_33_845 ();
 FILLER_ASAP7_75t_R FILLER_33_856 ();
 FILLER_ASAP7_75t_R FILLER_33_867 ();
 DECAPx4_ASAP7_75t_R FILLER_33_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_887 ();
 DECAPx10_ASAP7_75t_R FILLER_33_892 ();
 DECAPx4_ASAP7_75t_R FILLER_33_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_924 ();
 DECAPx6_ASAP7_75t_R FILLER_33_927 ();
 FILLER_ASAP7_75t_R FILLER_33_941 ();
 FILLER_ASAP7_75t_R FILLER_33_951 ();
 DECAPx4_ASAP7_75t_R FILLER_33_956 ();
 DECAPx2_ASAP7_75t_R FILLER_33_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_979 ();
 FILLER_ASAP7_75t_R FILLER_33_983 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_995 ();
 FILLER_ASAP7_75t_R FILLER_33_1010 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1073 ();
 DECAPx6_ASAP7_75t_R FILLER_33_1081 ();
 DECAPx1_ASAP7_75t_R FILLER_33_1095 ();
 FILLER_ASAP7_75t_R FILLER_33_1106 ();
 FILLER_ASAP7_75t_R FILLER_33_1114 ();
 DECAPx6_ASAP7_75t_R FILLER_33_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1142 ();
 FILLER_ASAP7_75t_R FILLER_33_1149 ();
 FILLER_ASAP7_75t_R FILLER_33_1163 ();
 FILLER_ASAP7_75t_R FILLER_33_1172 ();
 DECAPx4_ASAP7_75t_R FILLER_33_1181 ();
 DECAPx4_ASAP7_75t_R FILLER_33_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1204 ();
 DECAPx4_ASAP7_75t_R FILLER_33_1208 ();
 DECAPx6_ASAP7_75t_R FILLER_33_1226 ();
 FILLER_ASAP7_75t_R FILLER_33_1240 ();
 DECAPx2_ASAP7_75t_R FILLER_33_1254 ();
 DECAPx4_ASAP7_75t_R FILLER_33_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1273 ();
 FILLER_ASAP7_75t_R FILLER_33_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_33_1282 ();
 DECAPx1_ASAP7_75t_R FILLER_33_1304 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1308 ();
 FILLER_ASAP7_75t_R FILLER_33_1321 ();
 FILLER_ASAP7_75t_R FILLER_33_1349 ();
 FILLER_ASAP7_75t_R FILLER_33_1358 ();
 DECAPx4_ASAP7_75t_R FILLER_33_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_34_2 ();
 FILLER_ASAP7_75t_R FILLER_34_24 ();
 DECAPx2_ASAP7_75t_R FILLER_34_29 ();
 FILLER_ASAP7_75t_R FILLER_34_35 ();
 FILLER_ASAP7_75t_R FILLER_34_43 ();
 DECAPx6_ASAP7_75t_R FILLER_34_53 ();
 FILLER_ASAP7_75t_R FILLER_34_75 ();
 DECAPx10_ASAP7_75t_R FILLER_34_83 ();
 FILLER_ASAP7_75t_R FILLER_34_113 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_121 ();
 DECAPx6_ASAP7_75t_R FILLER_34_150 ();
 DECAPx1_ASAP7_75t_R FILLER_34_164 ();
 FILLER_ASAP7_75t_R FILLER_34_176 ();
 DECAPx2_ASAP7_75t_R FILLER_34_184 ();
 FILLER_ASAP7_75t_R FILLER_34_196 ();
 DECAPx10_ASAP7_75t_R FILLER_34_201 ();
 DECAPx2_ASAP7_75t_R FILLER_34_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_229 ();
 DECAPx10_ASAP7_75t_R FILLER_34_238 ();
 DECAPx2_ASAP7_75t_R FILLER_34_260 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_266 ();
 DECAPx2_ASAP7_75t_R FILLER_34_275 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_281 ();
 FILLER_ASAP7_75t_R FILLER_34_290 ();
 FILLER_ASAP7_75t_R FILLER_34_298 ();
 FILLER_ASAP7_75t_R FILLER_34_307 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_315 ();
 FILLER_ASAP7_75t_R FILLER_34_324 ();
 DECAPx2_ASAP7_75t_R FILLER_34_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_335 ();
 DECAPx10_ASAP7_75t_R FILLER_34_344 ();
 DECAPx2_ASAP7_75t_R FILLER_34_366 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_372 ();
 DECAPx6_ASAP7_75t_R FILLER_34_401 ();
 DECAPx4_ASAP7_75t_R FILLER_34_423 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_439 ();
 FILLER_ASAP7_75t_R FILLER_34_449 ();
 DECAPx1_ASAP7_75t_R FILLER_34_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_461 ();
 FILLER_ASAP7_75t_R FILLER_34_464 ();
 FILLER_ASAP7_75t_R FILLER_34_472 ();
 DECAPx1_ASAP7_75t_R FILLER_34_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_481 ();
 DECAPx10_ASAP7_75t_R FILLER_34_488 ();
 FILLER_ASAP7_75t_R FILLER_34_548 ();
 DECAPx2_ASAP7_75t_R FILLER_34_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_563 ();
 DECAPx6_ASAP7_75t_R FILLER_34_573 ();
 DECAPx1_ASAP7_75t_R FILLER_34_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_591 ();
 DECAPx6_ASAP7_75t_R FILLER_34_598 ();
 DECAPx2_ASAP7_75t_R FILLER_34_612 ();
 DECAPx2_ASAP7_75t_R FILLER_34_627 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_633 ();
 DECAPx2_ASAP7_75t_R FILLER_34_650 ();
 DECAPx2_ASAP7_75t_R FILLER_34_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_671 ();
 FILLER_ASAP7_75t_R FILLER_34_681 ();
 DECAPx2_ASAP7_75t_R FILLER_34_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_695 ();
 DECAPx1_ASAP7_75t_R FILLER_34_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_722 ();
 FILLER_ASAP7_75t_R FILLER_34_739 ();
 FILLER_ASAP7_75t_R FILLER_34_750 ();
 FILLER_ASAP7_75t_R FILLER_34_755 ();
 DECAPx6_ASAP7_75t_R FILLER_34_763 ();
 DECAPx2_ASAP7_75t_R FILLER_34_777 ();
 FILLER_ASAP7_75t_R FILLER_34_789 ();
 DECAPx2_ASAP7_75t_R FILLER_34_797 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_803 ();
 DECAPx6_ASAP7_75t_R FILLER_34_820 ();
 DECAPx1_ASAP7_75t_R FILLER_34_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_838 ();
 DECAPx2_ASAP7_75t_R FILLER_34_842 ();
 FILLER_ASAP7_75t_R FILLER_34_848 ();
 DECAPx4_ASAP7_75t_R FILLER_34_853 ();
 FILLER_ASAP7_75t_R FILLER_34_863 ();
 DECAPx6_ASAP7_75t_R FILLER_34_885 ();
 DECAPx2_ASAP7_75t_R FILLER_34_899 ();
 FILLER_ASAP7_75t_R FILLER_34_911 ();
 DECAPx4_ASAP7_75t_R FILLER_34_919 ();
 DECAPx1_ASAP7_75t_R FILLER_34_955 ();
 FILLER_ASAP7_75t_R FILLER_34_965 ();
 FILLER_ASAP7_75t_R FILLER_34_993 ();
 FILLER_ASAP7_75t_R FILLER_34_1021 ();
 FILLER_ASAP7_75t_R FILLER_34_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_34_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1059 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_1065 ();
 DECAPx4_ASAP7_75t_R FILLER_34_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_34_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1129 ();
 DECAPx4_ASAP7_75t_R FILLER_34_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1155 ();
 DECAPx1_ASAP7_75t_R FILLER_34_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_34_1187 ();
 FILLER_ASAP7_75t_R FILLER_34_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1223 ();
 DECAPx6_ASAP7_75t_R FILLER_34_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_1261 ();
 DECAPx6_ASAP7_75t_R FILLER_34_1272 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_1286 ();
 DECAPx6_ASAP7_75t_R FILLER_34_1315 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_1329 ();
 DECAPx2_ASAP7_75t_R FILLER_34_1354 ();
 FILLER_ASAP7_75t_R FILLER_34_1360 ();
 DECAPx4_ASAP7_75t_R FILLER_34_1365 ();
 FILLER_ASAP7_75t_R FILLER_34_1375 ();
 DECAPx4_ASAP7_75t_R FILLER_35_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_12 ();
 FILLER_ASAP7_75t_R FILLER_35_19 ();
 DECAPx1_ASAP7_75t_R FILLER_35_27 ();
 DECAPx4_ASAP7_75t_R FILLER_35_34 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_44 ();
 DECAPx6_ASAP7_75t_R FILLER_35_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_69 ();
 DECAPx4_ASAP7_75t_R FILLER_35_78 ();
 FILLER_ASAP7_75t_R FILLER_35_94 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_102 ();
 DECAPx4_ASAP7_75t_R FILLER_35_113 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_123 ();
 DECAPx2_ASAP7_75t_R FILLER_35_132 ();
 FILLER_ASAP7_75t_R FILLER_35_144 ();
 FILLER_ASAP7_75t_R FILLER_35_152 ();
 DECAPx2_ASAP7_75t_R FILLER_35_160 ();
 FILLER_ASAP7_75t_R FILLER_35_166 ();
 DECAPx6_ASAP7_75t_R FILLER_35_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_190 ();
 FILLER_ASAP7_75t_R FILLER_35_194 ();
 DECAPx4_ASAP7_75t_R FILLER_35_202 ();
 FILLER_ASAP7_75t_R FILLER_35_212 ();
 DECAPx4_ASAP7_75t_R FILLER_35_220 ();
 FILLER_ASAP7_75t_R FILLER_35_230 ();
 DECAPx4_ASAP7_75t_R FILLER_35_240 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_250 ();
 DECAPx2_ASAP7_75t_R FILLER_35_261 ();
 FILLER_ASAP7_75t_R FILLER_35_275 ();
 DECAPx4_ASAP7_75t_R FILLER_35_283 ();
 DECAPx1_ASAP7_75t_R FILLER_35_296 ();
 DECAPx10_ASAP7_75t_R FILLER_35_308 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_330 ();
 DECAPx2_ASAP7_75t_R FILLER_35_340 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_346 ();
 FILLER_ASAP7_75t_R FILLER_35_355 ();
 FILLER_ASAP7_75t_R FILLER_35_365 ();
 DECAPx1_ASAP7_75t_R FILLER_35_373 ();
 DECAPx4_ASAP7_75t_R FILLER_35_383 ();
 FILLER_ASAP7_75t_R FILLER_35_393 ();
 FILLER_ASAP7_75t_R FILLER_35_401 ();
 DECAPx10_ASAP7_75t_R FILLER_35_411 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_441 ();
 DECAPx4_ASAP7_75t_R FILLER_35_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_464 ();
 DECAPx2_ASAP7_75t_R FILLER_35_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_479 ();
 FILLER_ASAP7_75t_R FILLER_35_506 ();
 FILLER_ASAP7_75t_R FILLER_35_515 ();
 FILLER_ASAP7_75t_R FILLER_35_524 ();
 FILLER_ASAP7_75t_R FILLER_35_546 ();
 FILLER_ASAP7_75t_R FILLER_35_557 ();
 DECAPx4_ASAP7_75t_R FILLER_35_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_579 ();
 FILLER_ASAP7_75t_R FILLER_35_589 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_599 ();
 FILLER_ASAP7_75t_R FILLER_35_612 ();
 DECAPx2_ASAP7_75t_R FILLER_35_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_627 ();
 FILLER_ASAP7_75t_R FILLER_35_636 ();
 DECAPx2_ASAP7_75t_R FILLER_35_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_650 ();
 DECAPx6_ASAP7_75t_R FILLER_35_657 ();
 DECAPx2_ASAP7_75t_R FILLER_35_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_677 ();
 DECAPx2_ASAP7_75t_R FILLER_35_688 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_694 ();
 FILLER_ASAP7_75t_R FILLER_35_703 ();
 FILLER_ASAP7_75t_R FILLER_35_711 ();
 DECAPx6_ASAP7_75t_R FILLER_35_719 ();
 DECAPx1_ASAP7_75t_R FILLER_35_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_737 ();
 FILLER_ASAP7_75t_R FILLER_35_744 ();
 FILLER_ASAP7_75t_R FILLER_35_754 ();
 FILLER_ASAP7_75t_R FILLER_35_764 ();
 DECAPx2_ASAP7_75t_R FILLER_35_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_779 ();
 FILLER_ASAP7_75t_R FILLER_35_787 ();
 DECAPx2_ASAP7_75t_R FILLER_35_797 ();
 FILLER_ASAP7_75t_R FILLER_35_803 ();
 DECAPx2_ASAP7_75t_R FILLER_35_811 ();
 FILLER_ASAP7_75t_R FILLER_35_823 ();
 DECAPx6_ASAP7_75t_R FILLER_35_828 ();
 DECAPx1_ASAP7_75t_R FILLER_35_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_846 ();
 DECAPx10_ASAP7_75t_R FILLER_35_853 ();
 DECAPx6_ASAP7_75t_R FILLER_35_875 ();
 FILLER_ASAP7_75t_R FILLER_35_889 ();
 FILLER_ASAP7_75t_R FILLER_35_898 ();
 DECAPx2_ASAP7_75t_R FILLER_35_906 ();
 FILLER_ASAP7_75t_R FILLER_35_912 ();
 FILLER_ASAP7_75t_R FILLER_35_923 ();
 FILLER_ASAP7_75t_R FILLER_35_927 ();
 DECAPx2_ASAP7_75t_R FILLER_35_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_941 ();
 DECAPx1_ASAP7_75t_R FILLER_35_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_952 ();
 FILLER_ASAP7_75t_R FILLER_35_963 ();
 DECAPx4_ASAP7_75t_R FILLER_35_971 ();
 FILLER_ASAP7_75t_R FILLER_35_981 ();
 DECAPx6_ASAP7_75t_R FILLER_35_989 ();
 FILLER_ASAP7_75t_R FILLER_35_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_35_1011 ();
 FILLER_ASAP7_75t_R FILLER_35_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_35_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_35_1062 ();
 FILLER_ASAP7_75t_R FILLER_35_1074 ();
 FILLER_ASAP7_75t_R FILLER_35_1082 ();
 FILLER_ASAP7_75t_R FILLER_35_1094 ();
 FILLER_ASAP7_75t_R FILLER_35_1106 ();
 DECAPx4_ASAP7_75t_R FILLER_35_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_35_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_1153 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_35_1176 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_1182 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_1192 ();
 FILLER_ASAP7_75t_R FILLER_35_1207 ();
 DECAPx6_ASAP7_75t_R FILLER_35_1215 ();
 DECAPx1_ASAP7_75t_R FILLER_35_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_35_1243 ();
 DECAPx2_ASAP7_75t_R FILLER_35_1256 ();
 FILLER_ASAP7_75t_R FILLER_35_1288 ();
 FILLER_ASAP7_75t_R FILLER_35_1298 ();
 FILLER_ASAP7_75t_R FILLER_35_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_35_1315 ();
 DECAPx4_ASAP7_75t_R FILLER_35_1337 ();
 FILLER_ASAP7_75t_R FILLER_35_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_35_1371 ();
 DECAPx1_ASAP7_75t_R FILLER_36_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_6 ();
 DECAPx2_ASAP7_75t_R FILLER_36_33 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_47 ();
 DECAPx10_ASAP7_75t_R FILLER_36_56 ();
 DECAPx4_ASAP7_75t_R FILLER_36_78 ();
 FILLER_ASAP7_75t_R FILLER_36_96 ();
 DECAPx10_ASAP7_75t_R FILLER_36_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_128 ();
 DECAPx4_ASAP7_75t_R FILLER_36_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_145 ();
 DECAPx10_ASAP7_75t_R FILLER_36_154 ();
 DECAPx4_ASAP7_75t_R FILLER_36_176 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_186 ();
 FILLER_ASAP7_75t_R FILLER_36_195 ();
 FILLER_ASAP7_75t_R FILLER_36_203 ();
 DECAPx6_ASAP7_75t_R FILLER_36_231 ();
 FILLER_ASAP7_75t_R FILLER_36_251 ();
 DECAPx2_ASAP7_75t_R FILLER_36_261 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_267 ();
 DECAPx10_ASAP7_75t_R FILLER_36_292 ();
 DECAPx1_ASAP7_75t_R FILLER_36_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_318 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_322 ();
 DECAPx2_ASAP7_75t_R FILLER_36_331 ();
 DECAPx2_ASAP7_75t_R FILLER_36_347 ();
 DECAPx10_ASAP7_75t_R FILLER_36_361 ();
 DECAPx6_ASAP7_75t_R FILLER_36_383 ();
 DECAPx2_ASAP7_75t_R FILLER_36_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_403 ();
 DECAPx4_ASAP7_75t_R FILLER_36_407 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_417 ();
 DECAPx4_ASAP7_75t_R FILLER_36_426 ();
 FILLER_ASAP7_75t_R FILLER_36_436 ();
 FILLER_ASAP7_75t_R FILLER_36_460 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_464 ();
 DECAPx2_ASAP7_75t_R FILLER_36_475 ();
 DECAPx2_ASAP7_75t_R FILLER_36_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_493 ();
 DECAPx2_ASAP7_75t_R FILLER_36_497 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_503 ();
 FILLER_ASAP7_75t_R FILLER_36_526 ();
 FILLER_ASAP7_75t_R FILLER_36_548 ();
 DECAPx10_ASAP7_75t_R FILLER_36_556 ();
 DECAPx2_ASAP7_75t_R FILLER_36_578 ();
 DECAPx1_ASAP7_75t_R FILLER_36_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_594 ();
 FILLER_ASAP7_75t_R FILLER_36_598 ();
 FILLER_ASAP7_75t_R FILLER_36_606 ();
 DECAPx6_ASAP7_75t_R FILLER_36_615 ();
 DECAPx2_ASAP7_75t_R FILLER_36_629 ();
 DECAPx6_ASAP7_75t_R FILLER_36_641 ();
 DECAPx1_ASAP7_75t_R FILLER_36_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_665 ();
 DECAPx2_ASAP7_75t_R FILLER_36_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_675 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_682 ();
 DECAPx6_ASAP7_75t_R FILLER_36_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_705 ();
 FILLER_ASAP7_75t_R FILLER_36_712 ();
 DECAPx10_ASAP7_75t_R FILLER_36_722 ();
 DECAPx6_ASAP7_75t_R FILLER_36_744 ();
 FILLER_ASAP7_75t_R FILLER_36_765 ();
 FILLER_ASAP7_75t_R FILLER_36_775 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_780 ();
 DECAPx10_ASAP7_75t_R FILLER_36_789 ();
 DECAPx2_ASAP7_75t_R FILLER_36_811 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_817 ();
 DECAPx2_ASAP7_75t_R FILLER_36_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_834 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_845 ();
 DECAPx6_ASAP7_75t_R FILLER_36_855 ();
 FILLER_ASAP7_75t_R FILLER_36_869 ();
 FILLER_ASAP7_75t_R FILLER_36_877 ();
 DECAPx1_ASAP7_75t_R FILLER_36_885 ();
 DECAPx2_ASAP7_75t_R FILLER_36_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_915 ();
 FILLER_ASAP7_75t_R FILLER_36_919 ();
 DECAPx2_ASAP7_75t_R FILLER_36_947 ();
 FILLER_ASAP7_75t_R FILLER_36_953 ();
 DECAPx10_ASAP7_75t_R FILLER_36_961 ();
 DECAPx10_ASAP7_75t_R FILLER_36_983 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1005 ();
 DECAPx4_ASAP7_75t_R FILLER_36_1027 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_1037 ();
 FILLER_ASAP7_75t_R FILLER_36_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_36_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1139 ();
 FILLER_ASAP7_75t_R FILLER_36_1145 ();
 FILLER_ASAP7_75t_R FILLER_36_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_36_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1218 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1234 ();
 FILLER_ASAP7_75t_R FILLER_36_1240 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1254 ();
 FILLER_ASAP7_75t_R FILLER_36_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1274 ();
 FILLER_ASAP7_75t_R FILLER_36_1278 ();
 FILLER_ASAP7_75t_R FILLER_36_1290 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1298 ();
 FILLER_ASAP7_75t_R FILLER_36_1304 ();
 FILLER_ASAP7_75t_R FILLER_36_1312 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1321 ();
 FILLER_ASAP7_75t_R FILLER_36_1327 ();
 DECAPx1_ASAP7_75t_R FILLER_36_1332 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_1336 ();
 FILLER_ASAP7_75t_R FILLER_36_1343 ();
 DECAPx2_ASAP7_75t_R FILLER_36_1371 ();
 DECAPx6_ASAP7_75t_R FILLER_37_2 ();
 DECAPx2_ASAP7_75t_R FILLER_37_16 ();
 DECAPx2_ASAP7_75t_R FILLER_37_25 ();
 FILLER_ASAP7_75t_R FILLER_37_37 ();
 DECAPx1_ASAP7_75t_R FILLER_37_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_51 ();
 DECAPx2_ASAP7_75t_R FILLER_37_58 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_37_64 ();
 DECAPx2_ASAP7_75t_R FILLER_37_82 ();
 FILLER_ASAP7_75t_R FILLER_37_88 ();
 FILLER_ASAP7_75t_R FILLER_37_96 ();
 DECAPx2_ASAP7_75t_R FILLER_37_120 ();
 FILLER_ASAP7_75t_R FILLER_37_129 ();
 DECAPx2_ASAP7_75t_R FILLER_37_139 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_37_145 ();
 DECAPx6_ASAP7_75t_R FILLER_37_154 ();
 DECAPx1_ASAP7_75t_R FILLER_37_168 ();
 FILLER_ASAP7_75t_R FILLER_37_179 ();
 FILLER_ASAP7_75t_R FILLER_37_187 ();
 DECAPx4_ASAP7_75t_R FILLER_37_197 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_37_207 ();
 DECAPx1_ASAP7_75t_R FILLER_37_216 ();
 FILLER_ASAP7_75t_R FILLER_37_223 ();
 FILLER_ASAP7_75t_R FILLER_37_231 ();
 FILLER_ASAP7_75t_R FILLER_37_241 ();
 FILLER_ASAP7_75t_R FILLER_37_249 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_37_257 ();
 FILLER_ASAP7_75t_R FILLER_37_266 ();
 DECAPx10_ASAP7_75t_R FILLER_37_276 ();
 DECAPx6_ASAP7_75t_R FILLER_37_298 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_37_312 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_37_323 ();
 DECAPx1_ASAP7_75t_R FILLER_37_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_338 ();
 DECAPx6_ASAP7_75t_R FILLER_37_345 ();
 DECAPx2_ASAP7_75t_R FILLER_37_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_365 ();
 DECAPx4_ASAP7_75t_R FILLER_37_374 ();
 FILLER_ASAP7_75t_R FILLER_37_384 ();
 DECAPx4_ASAP7_75t_R FILLER_37_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_402 ();
 DECAPx6_ASAP7_75t_R FILLER_37_411 ();
 DECAPx2_ASAP7_75t_R FILLER_37_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_431 ();
 DECAPx2_ASAP7_75t_R FILLER_37_438 ();
 DECAPx6_ASAP7_75t_R FILLER_37_450 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_37_464 ();
 DECAPx10_ASAP7_75t_R FILLER_37_473 ();
 DECAPx1_ASAP7_75t_R FILLER_37_495 ();
 DECAPx2_ASAP7_75t_R FILLER_37_502 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_37_508 ();
 FILLER_ASAP7_75t_R FILLER_37_517 ();
 FILLER_ASAP7_75t_R FILLER_37_526 ();
 DECAPx2_ASAP7_75t_R FILLER_37_550 ();
 FILLER_ASAP7_75t_R FILLER_37_556 ();
 DECAPx2_ASAP7_75t_R FILLER_37_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_570 ();
 DECAPx6_ASAP7_75t_R FILLER_37_578 ();
 DECAPx1_ASAP7_75t_R FILLER_37_592 ();
 DECAPx6_ASAP7_75t_R FILLER_37_604 ();
 DECAPx2_ASAP7_75t_R FILLER_37_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_624 ();
 DECAPx2_ASAP7_75t_R FILLER_37_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_639 ();
 DECAPx2_ASAP7_75t_R FILLER_37_650 ();
 DECAPx6_ASAP7_75t_R FILLER_37_666 ();
 DECAPx1_ASAP7_75t_R FILLER_37_680 ();
 DECAPx2_ASAP7_75t_R FILLER_37_690 ();
 FILLER_ASAP7_75t_R FILLER_37_704 ();
 DECAPx6_ASAP7_75t_R FILLER_37_713 ();
 DECAPx1_ASAP7_75t_R FILLER_37_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_731 ();
 DECAPx10_ASAP7_75t_R FILLER_37_738 ();
 DECAPx6_ASAP7_75t_R FILLER_37_760 ();
 DECAPx1_ASAP7_75t_R FILLER_37_774 ();
 FILLER_ASAP7_75t_R FILLER_37_785 ();
 DECAPx4_ASAP7_75t_R FILLER_37_793 ();
 FILLER_ASAP7_75t_R FILLER_37_803 ();
 FILLER_ASAP7_75t_R FILLER_37_815 ();
 FILLER_ASAP7_75t_R FILLER_37_823 ();
 FILLER_ASAP7_75t_R FILLER_37_845 ();
 DECAPx1_ASAP7_75t_R FILLER_37_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_871 ();
 DECAPx4_ASAP7_75t_R FILLER_37_878 ();
 FILLER_ASAP7_75t_R FILLER_37_888 ();
 DECAPx6_ASAP7_75t_R FILLER_37_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_907 ();
 DECAPx6_ASAP7_75t_R FILLER_37_911 ();
 DECAPx2_ASAP7_75t_R FILLER_37_927 ();
 FILLER_ASAP7_75t_R FILLER_37_933 ();
 DECAPx6_ASAP7_75t_R FILLER_37_938 ();
 DECAPx1_ASAP7_75t_R FILLER_37_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_956 ();
 DECAPx2_ASAP7_75t_R FILLER_37_967 ();
 DECAPx2_ASAP7_75t_R FILLER_37_999 ();
 FILLER_ASAP7_75t_R FILLER_37_1005 ();
 DECAPx1_ASAP7_75t_R FILLER_37_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1021 ();
 FILLER_ASAP7_75t_R FILLER_37_1032 ();
 FILLER_ASAP7_75t_R FILLER_37_1046 ();
 DECAPx1_ASAP7_75t_R FILLER_37_1074 ();
 DECAPx6_ASAP7_75t_R FILLER_37_1084 ();
 DECAPx2_ASAP7_75t_R FILLER_37_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1104 ();
 FILLER_ASAP7_75t_R FILLER_37_1115 ();
 DECAPx4_ASAP7_75t_R FILLER_37_1125 ();
 FILLER_ASAP7_75t_R FILLER_37_1135 ();
 FILLER_ASAP7_75t_R FILLER_37_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1152 ();
 FILLER_ASAP7_75t_R FILLER_37_1174 ();
 DECAPx4_ASAP7_75t_R FILLER_37_1182 ();
 FILLER_ASAP7_75t_R FILLER_37_1198 ();
 DECAPx4_ASAP7_75t_R FILLER_37_1203 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_37_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_37_1272 ();
 DECAPx6_ASAP7_75t_R FILLER_37_1294 ();
 DECAPx2_ASAP7_75t_R FILLER_37_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_1314 ();
 DECAPx1_ASAP7_75t_R FILLER_37_1341 ();
 DECAPx2_ASAP7_75t_R FILLER_37_1352 ();
 FILLER_ASAP7_75t_R FILLER_37_1358 ();
 DECAPx6_ASAP7_75t_R FILLER_37_1363 ();
 DECAPx10_ASAP7_75t_R FILLER_38_2 ();
 DECAPx4_ASAP7_75t_R FILLER_38_24 ();
 DECAPx6_ASAP7_75t_R FILLER_38_40 ();
 DECAPx2_ASAP7_75t_R FILLER_38_54 ();
 FILLER_ASAP7_75t_R FILLER_38_66 ();
 FILLER_ASAP7_75t_R FILLER_38_74 ();
 DECAPx4_ASAP7_75t_R FILLER_38_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_92 ();
 DECAPx1_ASAP7_75t_R FILLER_38_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_103 ();
 DECAPx2_ASAP7_75t_R FILLER_38_130 ();
 FILLER_ASAP7_75t_R FILLER_38_136 ();
 FILLER_ASAP7_75t_R FILLER_38_146 ();
 DECAPx1_ASAP7_75t_R FILLER_38_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_164 ();
 DECAPx10_ASAP7_75t_R FILLER_38_173 ();
 DECAPx10_ASAP7_75t_R FILLER_38_195 ();
 DECAPx2_ASAP7_75t_R FILLER_38_217 ();
 FILLER_ASAP7_75t_R FILLER_38_229 ();
 DECAPx10_ASAP7_75t_R FILLER_38_239 ();
 DECAPx10_ASAP7_75t_R FILLER_38_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_283 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_38_290 ();
 FILLER_ASAP7_75t_R FILLER_38_296 ();
 FILLER_ASAP7_75t_R FILLER_38_304 ();
 DECAPx2_ASAP7_75t_R FILLER_38_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_318 ();
 FILLER_ASAP7_75t_R FILLER_38_327 ();
 DECAPx6_ASAP7_75t_R FILLER_38_336 ();
 FILLER_ASAP7_75t_R FILLER_38_356 ();
 FILLER_ASAP7_75t_R FILLER_38_364 ();
 DECAPx1_ASAP7_75t_R FILLER_38_374 ();
 DECAPx1_ASAP7_75t_R FILLER_38_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_408 ();
 FILLER_ASAP7_75t_R FILLER_38_417 ();
 FILLER_ASAP7_75t_R FILLER_38_426 ();
 DECAPx2_ASAP7_75t_R FILLER_38_454 ();
 FILLER_ASAP7_75t_R FILLER_38_460 ();
 DECAPx10_ASAP7_75t_R FILLER_38_464 ();
 DECAPx1_ASAP7_75t_R FILLER_38_492 ();
 DECAPx2_ASAP7_75t_R FILLER_38_522 ();
 DECAPx2_ASAP7_75t_R FILLER_38_550 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_38_556 ();
 FILLER_ASAP7_75t_R FILLER_38_571 ();
 DECAPx6_ASAP7_75t_R FILLER_38_583 ();
 FILLER_ASAP7_75t_R FILLER_38_597 ();
 FILLER_ASAP7_75t_R FILLER_38_608 ();
 FILLER_ASAP7_75t_R FILLER_38_622 ();
 DECAPx1_ASAP7_75t_R FILLER_38_630 ();
 DECAPx1_ASAP7_75t_R FILLER_38_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_645 ();
 FILLER_ASAP7_75t_R FILLER_38_656 ();
 FILLER_ASAP7_75t_R FILLER_38_664 ();
 DECAPx2_ASAP7_75t_R FILLER_38_676 ();
 DECAPx10_ASAP7_75t_R FILLER_38_692 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_38_714 ();
 DECAPx1_ASAP7_75t_R FILLER_38_725 ();
 FILLER_ASAP7_75t_R FILLER_38_749 ();
 DECAPx4_ASAP7_75t_R FILLER_38_761 ();
 DECAPx1_ASAP7_75t_R FILLER_38_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_797 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_38_804 ();
 DECAPx10_ASAP7_75t_R FILLER_38_827 ();
 DECAPx2_ASAP7_75t_R FILLER_38_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_855 ();
 DECAPx4_ASAP7_75t_R FILLER_38_860 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_38_870 ();
 DECAPx4_ASAP7_75t_R FILLER_38_881 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_38_891 ();
 DECAPx6_ASAP7_75t_R FILLER_38_900 ();
 DECAPx2_ASAP7_75t_R FILLER_38_920 ();
 DECAPx1_ASAP7_75t_R FILLER_38_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_940 ();
 DECAPx1_ASAP7_75t_R FILLER_38_951 ();
 FILLER_ASAP7_75t_R FILLER_38_958 ();
 DECAPx2_ASAP7_75t_R FILLER_38_986 ();
 FILLER_ASAP7_75t_R FILLER_38_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_38_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1024 ();
 DECAPx1_ASAP7_75t_R FILLER_38_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1049 ();
 DECAPx4_ASAP7_75t_R FILLER_38_1056 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_38_1066 ();
 FILLER_ASAP7_75t_R FILLER_38_1076 ();
 DECAPx4_ASAP7_75t_R FILLER_38_1090 ();
 FILLER_ASAP7_75t_R FILLER_38_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_38_1176 ();
 DECAPx6_ASAP7_75t_R FILLER_38_1198 ();
 DECAPx2_ASAP7_75t_R FILLER_38_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1218 ();
 FILLER_ASAP7_75t_R FILLER_38_1239 ();
 FILLER_ASAP7_75t_R FILLER_38_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_38_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_38_1284 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_38_1294 ();
 DECAPx2_ASAP7_75t_R FILLER_38_1305 ();
 FILLER_ASAP7_75t_R FILLER_38_1314 ();
 FILLER_ASAP7_75t_R FILLER_38_1322 ();
 FILLER_ASAP7_75t_R FILLER_38_1330 ();
 DECAPx6_ASAP7_75t_R FILLER_38_1358 ();
 DECAPx1_ASAP7_75t_R FILLER_38_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_39_2 ();
 FILLER_ASAP7_75t_R FILLER_39_8 ();
 DECAPx6_ASAP7_75t_R FILLER_39_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_50 ();
 DECAPx2_ASAP7_75t_R FILLER_39_57 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_63 ();
 DECAPx1_ASAP7_75t_R FILLER_39_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_78 ();
 DECAPx2_ASAP7_75t_R FILLER_39_85 ();
 FILLER_ASAP7_75t_R FILLER_39_91 ();
 DECAPx2_ASAP7_75t_R FILLER_39_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_105 ();
 FILLER_ASAP7_75t_R FILLER_39_112 ();
 FILLER_ASAP7_75t_R FILLER_39_120 ();
 DECAPx2_ASAP7_75t_R FILLER_39_125 ();
 DECAPx6_ASAP7_75t_R FILLER_39_137 ();
 DECAPx2_ASAP7_75t_R FILLER_39_151 ();
 FILLER_ASAP7_75t_R FILLER_39_163 ();
 FILLER_ASAP7_75t_R FILLER_39_173 ();
 DECAPx2_ASAP7_75t_R FILLER_39_182 ();
 FILLER_ASAP7_75t_R FILLER_39_188 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_196 ();
 FILLER_ASAP7_75t_R FILLER_39_205 ();
 DECAPx1_ASAP7_75t_R FILLER_39_213 ();
 DECAPx6_ASAP7_75t_R FILLER_39_223 ();
 DECAPx10_ASAP7_75t_R FILLER_39_243 ();
 DECAPx1_ASAP7_75t_R FILLER_39_271 ();
 FILLER_ASAP7_75t_R FILLER_39_301 ();
 FILLER_ASAP7_75t_R FILLER_39_311 ();
 DECAPx10_ASAP7_75t_R FILLER_39_319 ();
 DECAPx2_ASAP7_75t_R FILLER_39_341 ();
 DECAPx1_ASAP7_75t_R FILLER_39_355 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_365 ();
 DECAPx2_ASAP7_75t_R FILLER_39_374 ();
 FILLER_ASAP7_75t_R FILLER_39_380 ();
 DECAPx1_ASAP7_75t_R FILLER_39_388 ();
 DECAPx1_ASAP7_75t_R FILLER_39_395 ();
 FILLER_ASAP7_75t_R FILLER_39_405 ();
 DECAPx10_ASAP7_75t_R FILLER_39_410 ();
 DECAPx4_ASAP7_75t_R FILLER_39_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_442 ();
 DECAPx2_ASAP7_75t_R FILLER_39_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_452 ();
 DECAPx2_ASAP7_75t_R FILLER_39_461 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_482 ();
 FILLER_ASAP7_75t_R FILLER_39_511 ();
 FILLER_ASAP7_75t_R FILLER_39_516 ();
 FILLER_ASAP7_75t_R FILLER_39_524 ();
 DECAPx2_ASAP7_75t_R FILLER_39_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_552 ();
 DECAPx2_ASAP7_75t_R FILLER_39_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_565 ();
 DECAPx4_ASAP7_75t_R FILLER_39_572 ();
 DECAPx4_ASAP7_75t_R FILLER_39_589 ();
 DECAPx1_ASAP7_75t_R FILLER_39_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_609 ();
 DECAPx10_ASAP7_75t_R FILLER_39_616 ();
 DECAPx1_ASAP7_75t_R FILLER_39_638 ();
 DECAPx4_ASAP7_75t_R FILLER_39_648 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_658 ();
 FILLER_ASAP7_75t_R FILLER_39_668 ();
 DECAPx10_ASAP7_75t_R FILLER_39_678 ();
 DECAPx1_ASAP7_75t_R FILLER_39_700 ();
 FILLER_ASAP7_75t_R FILLER_39_714 ();
 DECAPx10_ASAP7_75t_R FILLER_39_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_746 ();
 FILLER_ASAP7_75t_R FILLER_39_753 ();
 DECAPx1_ASAP7_75t_R FILLER_39_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_767 ();
 FILLER_ASAP7_75t_R FILLER_39_774 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_783 ();
 DECAPx2_ASAP7_75t_R FILLER_39_794 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_800 ();
 DECAPx10_ASAP7_75t_R FILLER_39_811 ();
 DECAPx10_ASAP7_75t_R FILLER_39_833 ();
 DECAPx6_ASAP7_75t_R FILLER_39_855 ();
 DECAPx1_ASAP7_75t_R FILLER_39_869 ();
 FILLER_ASAP7_75t_R FILLER_39_893 ();
 DECAPx2_ASAP7_75t_R FILLER_39_901 ();
 FILLER_ASAP7_75t_R FILLER_39_907 ();
 DECAPx2_ASAP7_75t_R FILLER_39_917 ();
 FILLER_ASAP7_75t_R FILLER_39_923 ();
 DECAPx2_ASAP7_75t_R FILLER_39_927 ();
 FILLER_ASAP7_75t_R FILLER_39_945 ();
 DECAPx6_ASAP7_75t_R FILLER_39_957 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_971 ();
 DECAPx1_ASAP7_75t_R FILLER_39_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_981 ();
 FILLER_ASAP7_75t_R FILLER_39_989 ();
 DECAPx2_ASAP7_75t_R FILLER_39_997 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_39_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1038 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_1044 ();
 DECAPx4_ASAP7_75t_R FILLER_39_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1091 ();
 FILLER_ASAP7_75t_R FILLER_39_1097 ();
 FILLER_ASAP7_75t_R FILLER_39_1107 ();
 FILLER_ASAP7_75t_R FILLER_39_1117 ();
 DECAPx1_ASAP7_75t_R FILLER_39_1122 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_1134 ();
 DECAPx4_ASAP7_75t_R FILLER_39_1140 ();
 FILLER_ASAP7_75t_R FILLER_39_1150 ();
 FILLER_ASAP7_75t_R FILLER_39_1178 ();
 FILLER_ASAP7_75t_R FILLER_39_1186 ();
 FILLER_ASAP7_75t_R FILLER_39_1208 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_1216 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1229 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_1235 ();
 DECAPx1_ASAP7_75t_R FILLER_39_1264 ();
 FILLER_ASAP7_75t_R FILLER_39_1271 ();
 FILLER_ASAP7_75t_R FILLER_39_1299 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1327 ();
 DECAPx1_ASAP7_75t_R FILLER_39_1340 ();
 FILLER_ASAP7_75t_R FILLER_39_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_39_1371 ();
 DECAPx2_ASAP7_75t_R FILLER_40_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_40_8 ();
 FILLER_ASAP7_75t_R FILLER_40_17 ();
 DECAPx1_ASAP7_75t_R FILLER_40_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_29 ();
 FILLER_ASAP7_75t_R FILLER_40_56 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_40_61 ();
 FILLER_ASAP7_75t_R FILLER_40_70 ();
 DECAPx2_ASAP7_75t_R FILLER_40_80 ();
 FILLER_ASAP7_75t_R FILLER_40_92 ();
 DECAPx6_ASAP7_75t_R FILLER_40_102 ();
 DECAPx1_ASAP7_75t_R FILLER_40_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_120 ();
 FILLER_ASAP7_75t_R FILLER_40_127 ();
 DECAPx10_ASAP7_75t_R FILLER_40_132 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_40_154 ();
 DECAPx2_ASAP7_75t_R FILLER_40_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_166 ();
 DECAPx6_ASAP7_75t_R FILLER_40_173 ();
 FILLER_ASAP7_75t_R FILLER_40_195 ();
 DECAPx2_ASAP7_75t_R FILLER_40_207 ();
 DECAPx1_ASAP7_75t_R FILLER_40_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_243 ();
 FILLER_ASAP7_75t_R FILLER_40_250 ();
 DECAPx1_ASAP7_75t_R FILLER_40_258 ();
 FILLER_ASAP7_75t_R FILLER_40_268 ();
 DECAPx1_ASAP7_75t_R FILLER_40_276 ();
 DECAPx1_ASAP7_75t_R FILLER_40_286 ();
 DECAPx2_ASAP7_75t_R FILLER_40_293 ();
 DECAPx10_ASAP7_75t_R FILLER_40_305 ();
 DECAPx2_ASAP7_75t_R FILLER_40_327 ();
 DECAPx4_ASAP7_75t_R FILLER_40_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_349 ();
 DECAPx10_ASAP7_75t_R FILLER_40_357 ();
 DECAPx4_ASAP7_75t_R FILLER_40_379 ();
 DECAPx2_ASAP7_75t_R FILLER_40_395 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_40_401 ();
 FILLER_ASAP7_75t_R FILLER_40_410 ();
 DECAPx2_ASAP7_75t_R FILLER_40_420 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_40_426 ();
 FILLER_ASAP7_75t_R FILLER_40_435 ();
 DECAPx4_ASAP7_75t_R FILLER_40_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_453 ();
 DECAPx1_ASAP7_75t_R FILLER_40_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_461 ();
 FILLER_ASAP7_75t_R FILLER_40_464 ();
 FILLER_ASAP7_75t_R FILLER_40_474 ();
 DECAPx2_ASAP7_75t_R FILLER_40_482 ();
 FILLER_ASAP7_75t_R FILLER_40_488 ();
 FILLER_ASAP7_75t_R FILLER_40_496 ();
 FILLER_ASAP7_75t_R FILLER_40_504 ();
 FILLER_ASAP7_75t_R FILLER_40_509 ();
 FILLER_ASAP7_75t_R FILLER_40_517 ();
 DECAPx2_ASAP7_75t_R FILLER_40_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_547 ();
 DECAPx2_ASAP7_75t_R FILLER_40_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_562 ();
 DECAPx2_ASAP7_75t_R FILLER_40_575 ();
 FILLER_ASAP7_75t_R FILLER_40_588 ();
 FILLER_ASAP7_75t_R FILLER_40_596 ();
 DECAPx6_ASAP7_75t_R FILLER_40_605 ();
 FILLER_ASAP7_75t_R FILLER_40_619 ();
 DECAPx10_ASAP7_75t_R FILLER_40_627 ();
 DECAPx4_ASAP7_75t_R FILLER_40_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_659 ();
 FILLER_ASAP7_75t_R FILLER_40_667 ();
 DECAPx2_ASAP7_75t_R FILLER_40_679 ();
 DECAPx2_ASAP7_75t_R FILLER_40_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_700 ();
 FILLER_ASAP7_75t_R FILLER_40_713 ();
 DECAPx4_ASAP7_75t_R FILLER_40_722 ();
 FILLER_ASAP7_75t_R FILLER_40_738 ();
 DECAPx6_ASAP7_75t_R FILLER_40_743 ();
 FILLER_ASAP7_75t_R FILLER_40_757 ();
 FILLER_ASAP7_75t_R FILLER_40_762 ();
 DECAPx4_ASAP7_75t_R FILLER_40_773 ();
 FILLER_ASAP7_75t_R FILLER_40_783 ();
 DECAPx4_ASAP7_75t_R FILLER_40_805 ();
 FILLER_ASAP7_75t_R FILLER_40_815 ();
 DECAPx2_ASAP7_75t_R FILLER_40_843 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_40_849 ();
 FILLER_ASAP7_75t_R FILLER_40_859 ();
 DECAPx2_ASAP7_75t_R FILLER_40_867 ();
 FILLER_ASAP7_75t_R FILLER_40_873 ();
 DECAPx4_ASAP7_75t_R FILLER_40_881 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_40_891 ();
 DECAPx4_ASAP7_75t_R FILLER_40_902 ();
 FILLER_ASAP7_75t_R FILLER_40_918 ();
 DECAPx10_ASAP7_75t_R FILLER_40_926 ();
 DECAPx6_ASAP7_75t_R FILLER_40_948 ();
 DECAPx1_ASAP7_75t_R FILLER_40_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_966 ();
 FILLER_ASAP7_75t_R FILLER_40_973 ();
 DECAPx2_ASAP7_75t_R FILLER_40_982 ();
 DECAPx10_ASAP7_75t_R FILLER_40_991 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_40_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_40_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1029 ();
 FILLER_ASAP7_75t_R FILLER_40_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_40_1070 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_40_1076 ();
 DECAPx6_ASAP7_75t_R FILLER_40_1082 ();
 FILLER_ASAP7_75t_R FILLER_40_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1101 ();
 FILLER_ASAP7_75t_R FILLER_40_1123 ();
 DECAPx4_ASAP7_75t_R FILLER_40_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_40_1152 ();
 FILLER_ASAP7_75t_R FILLER_40_1168 ();
 FILLER_ASAP7_75t_R FILLER_40_1196 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_40_1204 ();
 DECAPx4_ASAP7_75t_R FILLER_40_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1226 ();
 FILLER_ASAP7_75t_R FILLER_40_1239 ();
 DECAPx2_ASAP7_75t_R FILLER_40_1247 ();
 DECAPx4_ASAP7_75t_R FILLER_40_1256 ();
 FILLER_ASAP7_75t_R FILLER_40_1266 ();
 FILLER_ASAP7_75t_R FILLER_40_1276 ();
 FILLER_ASAP7_75t_R FILLER_40_1286 ();
 DECAPx1_ASAP7_75t_R FILLER_40_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1301 ();
 DECAPx6_ASAP7_75t_R FILLER_40_1323 ();
 DECAPx2_ASAP7_75t_R FILLER_40_1337 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_1343 ();
 DECAPx10_ASAP7_75t_R FILLER_40_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_40_1369 ();
 FILLER_ASAP7_75t_R FILLER_40_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_41_2 ();
 DECAPx6_ASAP7_75t_R FILLER_41_27 ();
 FILLER_ASAP7_75t_R FILLER_41_41 ();
 FILLER_ASAP7_75t_R FILLER_41_46 ();
 FILLER_ASAP7_75t_R FILLER_41_54 ();
 FILLER_ASAP7_75t_R FILLER_41_68 ();
 DECAPx10_ASAP7_75t_R FILLER_41_76 ();
 DECAPx4_ASAP7_75t_R FILLER_41_98 ();
 FILLER_ASAP7_75t_R FILLER_41_108 ();
 DECAPx2_ASAP7_75t_R FILLER_41_136 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_142 ();
 DECAPx6_ASAP7_75t_R FILLER_41_151 ();
 FILLER_ASAP7_75t_R FILLER_41_165 ();
 DECAPx6_ASAP7_75t_R FILLER_41_173 ();
 FILLER_ASAP7_75t_R FILLER_41_187 ();
 DECAPx4_ASAP7_75t_R FILLER_41_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_202 ();
 DECAPx2_ASAP7_75t_R FILLER_41_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_215 ();
 DECAPx1_ASAP7_75t_R FILLER_41_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_226 ();
 DECAPx2_ASAP7_75t_R FILLER_41_230 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_236 ();
 FILLER_ASAP7_75t_R FILLER_41_265 ();
 FILLER_ASAP7_75t_R FILLER_41_270 ();
 FILLER_ASAP7_75t_R FILLER_41_282 ();
 FILLER_ASAP7_75t_R FILLER_41_290 ();
 DECAPx10_ASAP7_75t_R FILLER_41_298 ();
 DECAPx2_ASAP7_75t_R FILLER_41_326 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_332 ();
 FILLER_ASAP7_75t_R FILLER_41_343 ();
 DECAPx6_ASAP7_75t_R FILLER_41_352 ();
 FILLER_ASAP7_75t_R FILLER_41_366 ();
 DECAPx4_ASAP7_75t_R FILLER_41_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_384 ();
 FILLER_ASAP7_75t_R FILLER_41_411 ();
 DECAPx2_ASAP7_75t_R FILLER_41_419 ();
 DECAPx4_ASAP7_75t_R FILLER_41_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_461 ();
 FILLER_ASAP7_75t_R FILLER_41_470 ();
 DECAPx10_ASAP7_75t_R FILLER_41_478 ();
 DECAPx4_ASAP7_75t_R FILLER_41_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_510 ();
 FILLER_ASAP7_75t_R FILLER_41_517 ();
 DECAPx2_ASAP7_75t_R FILLER_41_541 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_547 ();
 FILLER_ASAP7_75t_R FILLER_41_556 ();
 DECAPx2_ASAP7_75t_R FILLER_41_561 ();
 FILLER_ASAP7_75t_R FILLER_41_567 ();
 DECAPx2_ASAP7_75t_R FILLER_41_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_585 ();
 DECAPx10_ASAP7_75t_R FILLER_41_593 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_615 ();
 FILLER_ASAP7_75t_R FILLER_41_625 ();
 FILLER_ASAP7_75t_R FILLER_41_637 ();
 DECAPx4_ASAP7_75t_R FILLER_41_646 ();
 DECAPx10_ASAP7_75t_R FILLER_41_663 ();
 DECAPx2_ASAP7_75t_R FILLER_41_685 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_691 ();
 DECAPx6_ASAP7_75t_R FILLER_41_701 ();
 DECAPx1_ASAP7_75t_R FILLER_41_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_719 ();
 DECAPx6_ASAP7_75t_R FILLER_41_746 ();
 FILLER_ASAP7_75t_R FILLER_41_760 ();
 FILLER_ASAP7_75t_R FILLER_41_770 ();
 DECAPx10_ASAP7_75t_R FILLER_41_778 ();
 DECAPx6_ASAP7_75t_R FILLER_41_800 ();
 FILLER_ASAP7_75t_R FILLER_41_840 ();
 DECAPx1_ASAP7_75t_R FILLER_41_850 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_874 ();
 DECAPx10_ASAP7_75t_R FILLER_41_884 ();
 DECAPx6_ASAP7_75t_R FILLER_41_906 ();
 DECAPx1_ASAP7_75t_R FILLER_41_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_924 ();
 FILLER_ASAP7_75t_R FILLER_41_927 ();
 DECAPx2_ASAP7_75t_R FILLER_41_935 ();
 DECAPx10_ASAP7_75t_R FILLER_41_949 ();
 DECAPx6_ASAP7_75t_R FILLER_41_971 ();
 FILLER_ASAP7_75t_R FILLER_41_995 ();
 DECAPx1_ASAP7_75t_R FILLER_41_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1011 ();
 FILLER_ASAP7_75t_R FILLER_41_1038 ();
 FILLER_ASAP7_75t_R FILLER_41_1047 ();
 DECAPx1_ASAP7_75t_R FILLER_41_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1062 ();
 DECAPx6_ASAP7_75t_R FILLER_41_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1098 ();
 FILLER_ASAP7_75t_R FILLER_41_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1150 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_1164 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_41_1181 ();
 FILLER_ASAP7_75t_R FILLER_41_1188 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1198 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1210 ();
 FILLER_ASAP7_75t_R FILLER_41_1216 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1224 ();
 FILLER_ASAP7_75t_R FILLER_41_1230 ();
 DECAPx2_ASAP7_75t_R FILLER_41_1235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_41_1276 ();
 DECAPx6_ASAP7_75t_R FILLER_41_1298 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_1312 ();
 FILLER_ASAP7_75t_R FILLER_41_1320 ();
 FILLER_ASAP7_75t_R FILLER_41_1328 ();
 FILLER_ASAP7_75t_R FILLER_41_1356 ();
 DECAPx4_ASAP7_75t_R FILLER_41_1364 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_1374 ();
 DECAPx10_ASAP7_75t_R FILLER_42_2 ();
 DECAPx4_ASAP7_75t_R FILLER_42_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_34 ();
 DECAPx6_ASAP7_75t_R FILLER_42_41 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_55 ();
 DECAPx10_ASAP7_75t_R FILLER_42_84 ();
 DECAPx1_ASAP7_75t_R FILLER_42_106 ();
 FILLER_ASAP7_75t_R FILLER_42_116 ();
 DECAPx1_ASAP7_75t_R FILLER_42_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_128 ();
 FILLER_ASAP7_75t_R FILLER_42_155 ();
 DECAPx1_ASAP7_75t_R FILLER_42_183 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_193 ();
 DECAPx10_ASAP7_75t_R FILLER_42_199 ();
 DECAPx10_ASAP7_75t_R FILLER_42_221 ();
 DECAPx6_ASAP7_75t_R FILLER_42_243 ();
 DECAPx6_ASAP7_75t_R FILLER_42_263 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_277 ();
 DECAPx2_ASAP7_75t_R FILLER_42_306 ();
 DECAPx6_ASAP7_75t_R FILLER_42_338 ();
 DECAPx1_ASAP7_75t_R FILLER_42_352 ();
 DECAPx1_ASAP7_75t_R FILLER_42_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_386 ();
 DECAPx2_ASAP7_75t_R FILLER_42_393 ();
 DECAPx10_ASAP7_75t_R FILLER_42_402 ();
 DECAPx4_ASAP7_75t_R FILLER_42_424 ();
 FILLER_ASAP7_75t_R FILLER_42_440 ();
 DECAPx6_ASAP7_75t_R FILLER_42_445 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_459 ();
 FILLER_ASAP7_75t_R FILLER_42_464 ();
 DECAPx6_ASAP7_75t_R FILLER_42_472 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_486 ();
 DECAPx6_ASAP7_75t_R FILLER_42_495 ();
 DECAPx2_ASAP7_75t_R FILLER_42_509 ();
 DECAPx2_ASAP7_75t_R FILLER_42_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_529 ();
 DECAPx6_ASAP7_75t_R FILLER_42_537 ();
 DECAPx10_ASAP7_75t_R FILLER_42_557 ();
 DECAPx4_ASAP7_75t_R FILLER_42_585 ();
 FILLER_ASAP7_75t_R FILLER_42_595 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_604 ();
 DECAPx2_ASAP7_75t_R FILLER_42_613 ();
 DECAPx2_ASAP7_75t_R FILLER_42_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_631 ();
 FILLER_ASAP7_75t_R FILLER_42_638 ();
 DECAPx2_ASAP7_75t_R FILLER_42_647 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_653 ();
 FILLER_ASAP7_75t_R FILLER_42_663 ();
 DECAPx2_ASAP7_75t_R FILLER_42_672 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_678 ();
 DECAPx4_ASAP7_75t_R FILLER_42_689 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_699 ();
 DECAPx10_ASAP7_75t_R FILLER_42_709 ();
 DECAPx1_ASAP7_75t_R FILLER_42_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_735 ();
 DECAPx1_ASAP7_75t_R FILLER_42_739 ();
 DECAPx1_ASAP7_75t_R FILLER_42_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_754 ();
 DECAPx4_ASAP7_75t_R FILLER_42_771 ();
 DECAPx2_ASAP7_75t_R FILLER_42_787 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_793 ();
 DECAPx1_ASAP7_75t_R FILLER_42_799 ();
 FILLER_ASAP7_75t_R FILLER_42_829 ();
 FILLER_ASAP7_75t_R FILLER_42_834 ();
 DECAPx1_ASAP7_75t_R FILLER_42_839 ();
 DECAPx10_ASAP7_75t_R FILLER_42_851 ();
 FILLER_ASAP7_75t_R FILLER_42_873 ();
 DECAPx2_ASAP7_75t_R FILLER_42_879 ();
 FILLER_ASAP7_75t_R FILLER_42_885 ();
 DECAPx4_ASAP7_75t_R FILLER_42_894 ();
 FILLER_ASAP7_75t_R FILLER_42_911 ();
 DECAPx2_ASAP7_75t_R FILLER_42_919 ();
 FILLER_ASAP7_75t_R FILLER_42_932 ();
 FILLER_ASAP7_75t_R FILLER_42_960 ();
 DECAPx4_ASAP7_75t_R FILLER_42_972 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_982 ();
 FILLER_ASAP7_75t_R FILLER_42_1005 ();
 DECAPx4_ASAP7_75t_R FILLER_42_1013 ();
 FILLER_ASAP7_75t_R FILLER_42_1023 ();
 FILLER_ASAP7_75t_R FILLER_42_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1036 ();
 DECAPx4_ASAP7_75t_R FILLER_42_1058 ();
 FILLER_ASAP7_75t_R FILLER_42_1077 ();
 DECAPx2_ASAP7_75t_R FILLER_42_1085 ();
 FILLER_ASAP7_75t_R FILLER_42_1091 ();
 DECAPx2_ASAP7_75t_R FILLER_42_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1111 ();
 DECAPx6_ASAP7_75t_R FILLER_42_1138 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_42_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_42_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_1217 ();
 FILLER_ASAP7_75t_R FILLER_42_1244 ();
 FILLER_ASAP7_75t_R FILLER_42_1258 ();
 DECAPx6_ASAP7_75t_R FILLER_42_1270 ();
 DECAPx2_ASAP7_75t_R FILLER_42_1284 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1296 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1310 ();
 FILLER_ASAP7_75t_R FILLER_42_1340 ();
 DECAPx1_ASAP7_75t_R FILLER_42_1345 ();
 FILLER_ASAP7_75t_R FILLER_42_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_43_2 ();
 DECAPx1_ASAP7_75t_R FILLER_43_16 ();
 FILLER_ASAP7_75t_R FILLER_43_46 ();
 DECAPx4_ASAP7_75t_R FILLER_43_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_64 ();
 FILLER_ASAP7_75t_R FILLER_43_71 ();
 DECAPx6_ASAP7_75t_R FILLER_43_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_90 ();
 FILLER_ASAP7_75t_R FILLER_43_98 ();
 FILLER_ASAP7_75t_R FILLER_43_106 ();
 DECAPx1_ASAP7_75t_R FILLER_43_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_138 ();
 FILLER_ASAP7_75t_R FILLER_43_145 ();
 DECAPx4_ASAP7_75t_R FILLER_43_150 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_160 ();
 FILLER_ASAP7_75t_R FILLER_43_169 ();
 DECAPx2_ASAP7_75t_R FILLER_43_174 ();
 FILLER_ASAP7_75t_R FILLER_43_180 ();
 DECAPx2_ASAP7_75t_R FILLER_43_208 ();
 FILLER_ASAP7_75t_R FILLER_43_240 ();
 DECAPx4_ASAP7_75t_R FILLER_43_248 ();
 DECAPx2_ASAP7_75t_R FILLER_43_264 ();
 FILLER_ASAP7_75t_R FILLER_43_270 ();
 DECAPx6_ASAP7_75t_R FILLER_43_278 ();
 FILLER_ASAP7_75t_R FILLER_43_292 ();
 DECAPx1_ASAP7_75t_R FILLER_43_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_301 ();
 DECAPx2_ASAP7_75t_R FILLER_43_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_314 ();
 DECAPx2_ASAP7_75t_R FILLER_43_321 ();
 FILLER_ASAP7_75t_R FILLER_43_330 ();
 DECAPx2_ASAP7_75t_R FILLER_43_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_344 ();
 DECAPx4_ASAP7_75t_R FILLER_43_351 ();
 FILLER_ASAP7_75t_R FILLER_43_361 ();
 FILLER_ASAP7_75t_R FILLER_43_369 ();
 DECAPx10_ASAP7_75t_R FILLER_43_374 ();
 DECAPx6_ASAP7_75t_R FILLER_43_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_410 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_417 ();
 DECAPx2_ASAP7_75t_R FILLER_43_426 ();
 FILLER_ASAP7_75t_R FILLER_43_432 ();
 DECAPx4_ASAP7_75t_R FILLER_43_440 ();
 FILLER_ASAP7_75t_R FILLER_43_450 ();
 FILLER_ASAP7_75t_R FILLER_43_478 ();
 FILLER_ASAP7_75t_R FILLER_43_506 ();
 DECAPx1_ASAP7_75t_R FILLER_43_511 ();
 DECAPx2_ASAP7_75t_R FILLER_43_523 ();
 FILLER_ASAP7_75t_R FILLER_43_529 ();
 DECAPx4_ASAP7_75t_R FILLER_43_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_548 ();
 FILLER_ASAP7_75t_R FILLER_43_556 ();
 DECAPx4_ASAP7_75t_R FILLER_43_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_575 ();
 DECAPx2_ASAP7_75t_R FILLER_43_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_589 ();
 DECAPx1_ASAP7_75t_R FILLER_43_596 ();
 DECAPx2_ASAP7_75t_R FILLER_43_608 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_614 ();
 DECAPx6_ASAP7_75t_R FILLER_43_623 ();
 DECAPx1_ASAP7_75t_R FILLER_43_637 ();
 DECAPx4_ASAP7_75t_R FILLER_43_648 ();
 FILLER_ASAP7_75t_R FILLER_43_658 ();
 FILLER_ASAP7_75t_R FILLER_43_670 ();
 FILLER_ASAP7_75t_R FILLER_43_678 ();
 DECAPx1_ASAP7_75t_R FILLER_43_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_694 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_702 ();
 DECAPx2_ASAP7_75t_R FILLER_43_714 ();
 FILLER_ASAP7_75t_R FILLER_43_720 ();
 FILLER_ASAP7_75t_R FILLER_43_748 ();
 DECAPx2_ASAP7_75t_R FILLER_43_756 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_762 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_774 ();
 DECAPx2_ASAP7_75t_R FILLER_43_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_786 ();
 DECAPx1_ASAP7_75t_R FILLER_43_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_817 ();
 DECAPx10_ASAP7_75t_R FILLER_43_821 ();
 DECAPx1_ASAP7_75t_R FILLER_43_843 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_857 ();
 DECAPx4_ASAP7_75t_R FILLER_43_874 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_884 ();
 DECAPx2_ASAP7_75t_R FILLER_43_895 ();
 DECAPx1_ASAP7_75t_R FILLER_43_921 ();
 DECAPx6_ASAP7_75t_R FILLER_43_927 ();
 DECAPx2_ASAP7_75t_R FILLER_43_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_947 ();
 DECAPx1_ASAP7_75t_R FILLER_43_951 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_963 ();
 FILLER_ASAP7_75t_R FILLER_43_976 ();
 DECAPx6_ASAP7_75t_R FILLER_43_984 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1024 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1046 ();
 FILLER_ASAP7_75t_R FILLER_43_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_43_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_43_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_43_1159 ();
 DECAPx6_ASAP7_75t_R FILLER_43_1181 ();
 FILLER_ASAP7_75t_R FILLER_43_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1215 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_1221 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1227 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1241 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_1247 ();
 DECAPx1_ASAP7_75t_R FILLER_43_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1264 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_1275 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_1284 ();
 FILLER_ASAP7_75t_R FILLER_43_1313 ();
 DECAPx4_ASAP7_75t_R FILLER_43_1321 ();
 FILLER_ASAP7_75t_R FILLER_43_1338 ();
 DECAPx1_ASAP7_75t_R FILLER_43_1346 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1350 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1358 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_1364 ();
 DECAPx2_ASAP7_75t_R FILLER_43_1368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_1374 ();
 DECAPx4_ASAP7_75t_R FILLER_44_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_44_12 ();
 DECAPx4_ASAP7_75t_R FILLER_44_21 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_44_31 ();
 DECAPx2_ASAP7_75t_R FILLER_44_37 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_44_43 ();
 DECAPx10_ASAP7_75t_R FILLER_44_49 ();
 DECAPx6_ASAP7_75t_R FILLER_44_71 ();
 DECAPx2_ASAP7_75t_R FILLER_44_85 ();
 FILLER_ASAP7_75t_R FILLER_44_99 ();
 FILLER_ASAP7_75t_R FILLER_44_107 ();
 DECAPx2_ASAP7_75t_R FILLER_44_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_121 ();
 DECAPx2_ASAP7_75t_R FILLER_44_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_131 ();
 DECAPx2_ASAP7_75t_R FILLER_44_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_145 ();
 DECAPx10_ASAP7_75t_R FILLER_44_152 ();
 DECAPx4_ASAP7_75t_R FILLER_44_174 ();
 DECAPx10_ASAP7_75t_R FILLER_44_190 ();
 DECAPx2_ASAP7_75t_R FILLER_44_212 ();
 DECAPx1_ASAP7_75t_R FILLER_44_224 ();
 DECAPx1_ASAP7_75t_R FILLER_44_254 ();
 DECAPx2_ASAP7_75t_R FILLER_44_266 ();
 FILLER_ASAP7_75t_R FILLER_44_294 ();
 DECAPx1_ASAP7_75t_R FILLER_44_322 ();
 DECAPx1_ASAP7_75t_R FILLER_44_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_333 ();
 DECAPx1_ASAP7_75t_R FILLER_44_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_346 ();
 DECAPx1_ASAP7_75t_R FILLER_44_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_357 ();
 DECAPx2_ASAP7_75t_R FILLER_44_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_370 ();
 DECAPx4_ASAP7_75t_R FILLER_44_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_391 ();
 DECAPx2_ASAP7_75t_R FILLER_44_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_404 ();
 FILLER_ASAP7_75t_R FILLER_44_431 ();
 DECAPx1_ASAP7_75t_R FILLER_44_436 ();
 FILLER_ASAP7_75t_R FILLER_44_447 ();
 DECAPx2_ASAP7_75t_R FILLER_44_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_461 ();
 FILLER_ASAP7_75t_R FILLER_44_464 ();
 FILLER_ASAP7_75t_R FILLER_44_472 ();
 DECAPx2_ASAP7_75t_R FILLER_44_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_483 ();
 DECAPx1_ASAP7_75t_R FILLER_44_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_494 ();
 DECAPx4_ASAP7_75t_R FILLER_44_498 ();
 FILLER_ASAP7_75t_R FILLER_44_508 ();
 FILLER_ASAP7_75t_R FILLER_44_518 ();
 FILLER_ASAP7_75t_R FILLER_44_526 ();
 DECAPx2_ASAP7_75t_R FILLER_44_548 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_44_554 ();
 DECAPx2_ASAP7_75t_R FILLER_44_565 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_44_571 ();
 DECAPx2_ASAP7_75t_R FILLER_44_584 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_44_590 ();
 FILLER_ASAP7_75t_R FILLER_44_601 ();
 DECAPx1_ASAP7_75t_R FILLER_44_613 ();
 DECAPx6_ASAP7_75t_R FILLER_44_625 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_44_639 ();
 DECAPx10_ASAP7_75t_R FILLER_44_649 ();
 DECAPx6_ASAP7_75t_R FILLER_44_671 ();
 DECAPx1_ASAP7_75t_R FILLER_44_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_689 ();
 DECAPx2_ASAP7_75t_R FILLER_44_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_702 ();
 DECAPx2_ASAP7_75t_R FILLER_44_709 ();
 FILLER_ASAP7_75t_R FILLER_44_721 ();
 DECAPx6_ASAP7_75t_R FILLER_44_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_757 ();
 FILLER_ASAP7_75t_R FILLER_44_765 ();
 FILLER_ASAP7_75t_R FILLER_44_773 ();
 DECAPx2_ASAP7_75t_R FILLER_44_781 ();
 DECAPx2_ASAP7_75t_R FILLER_44_796 ();
 DECAPx6_ASAP7_75t_R FILLER_44_805 ();
 DECAPx10_ASAP7_75t_R FILLER_44_826 ();
 DECAPx2_ASAP7_75t_R FILLER_44_852 ();
 FILLER_ASAP7_75t_R FILLER_44_862 ();
 DECAPx1_ASAP7_75t_R FILLER_44_870 ();
 FILLER_ASAP7_75t_R FILLER_44_884 ();
 DECAPx6_ASAP7_75t_R FILLER_44_892 ();
 DECAPx4_ASAP7_75t_R FILLER_44_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_921 ();
 DECAPx2_ASAP7_75t_R FILLER_44_931 ();
 FILLER_ASAP7_75t_R FILLER_44_937 ();
 DECAPx2_ASAP7_75t_R FILLER_44_945 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_44_951 ();
 DECAPx4_ASAP7_75t_R FILLER_44_957 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_44_967 ();
 DECAPx1_ASAP7_75t_R FILLER_44_996 ();
 DECAPx2_ASAP7_75t_R FILLER_44_1007 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1016 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_44_1038 ();
 FILLER_ASAP7_75t_R FILLER_44_1048 ();
 FILLER_ASAP7_75t_R FILLER_44_1056 ();
 FILLER_ASAP7_75t_R FILLER_44_1064 ();
 FILLER_ASAP7_75t_R FILLER_44_1069 ();
 DECAPx4_ASAP7_75t_R FILLER_44_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_44_1087 ();
 FILLER_ASAP7_75t_R FILLER_44_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1102 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_44_1124 ();
 DECAPx4_ASAP7_75t_R FILLER_44_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1140 ();
 FILLER_ASAP7_75t_R FILLER_44_1167 ();
 FILLER_ASAP7_75t_R FILLER_44_1181 ();
 FILLER_ASAP7_75t_R FILLER_44_1189 ();
 FILLER_ASAP7_75t_R FILLER_44_1198 ();
 FILLER_ASAP7_75t_R FILLER_44_1226 ();
 DECAPx6_ASAP7_75t_R FILLER_44_1234 ();
 DECAPx1_ASAP7_75t_R FILLER_44_1248 ();
 FILLER_ASAP7_75t_R FILLER_44_1260 ();
 DECAPx1_ASAP7_75t_R FILLER_44_1288 ();
 DECAPx1_ASAP7_75t_R FILLER_44_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1304 ();
 DECAPx4_ASAP7_75t_R FILLER_44_1312 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1322 ();
 DECAPx1_ASAP7_75t_R FILLER_44_1330 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_44_1341 ();
 DECAPx6_ASAP7_75t_R FILLER_44_1363 ();
 FILLER_ASAP7_75t_R FILLER_45_2 ();
 DECAPx10_ASAP7_75t_R FILLER_45_30 ();
 DECAPx6_ASAP7_75t_R FILLER_45_60 ();
 DECAPx1_ASAP7_75t_R FILLER_45_74 ();
 DECAPx1_ASAP7_75t_R FILLER_45_84 ();
 DECAPx1_ASAP7_75t_R FILLER_45_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_95 ();
 DECAPx6_ASAP7_75t_R FILLER_45_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_120 ();
 FILLER_ASAP7_75t_R FILLER_45_127 ();
 FILLER_ASAP7_75t_R FILLER_45_136 ();
 FILLER_ASAP7_75t_R FILLER_45_164 ();
 DECAPx10_ASAP7_75t_R FILLER_45_172 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_194 ();
 FILLER_ASAP7_75t_R FILLER_45_223 ();
 DECAPx1_ASAP7_75t_R FILLER_45_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_235 ();
 FILLER_ASAP7_75t_R FILLER_45_239 ();
 DECAPx1_ASAP7_75t_R FILLER_45_247 ();
 FILLER_ASAP7_75t_R FILLER_45_254 ();
 FILLER_ASAP7_75t_R FILLER_45_264 ();
 FILLER_ASAP7_75t_R FILLER_45_292 ();
 FILLER_ASAP7_75t_R FILLER_45_300 ();
 FILLER_ASAP7_75t_R FILLER_45_309 ();
 FILLER_ASAP7_75t_R FILLER_45_318 ();
 DECAPx10_ASAP7_75t_R FILLER_45_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_345 ();
 FILLER_ASAP7_75t_R FILLER_45_349 ();
 FILLER_ASAP7_75t_R FILLER_45_377 ();
 FILLER_ASAP7_75t_R FILLER_45_405 ();
 DECAPx4_ASAP7_75t_R FILLER_45_410 ();
 DECAPx4_ASAP7_75t_R FILLER_45_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_433 ();
 DECAPx1_ASAP7_75t_R FILLER_45_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_446 ();
 DECAPx1_ASAP7_75t_R FILLER_45_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_461 ();
 DECAPx6_ASAP7_75t_R FILLER_45_468 ();
 DECAPx2_ASAP7_75t_R FILLER_45_482 ();
 DECAPx2_ASAP7_75t_R FILLER_45_494 ();
 FILLER_ASAP7_75t_R FILLER_45_500 ();
 FILLER_ASAP7_75t_R FILLER_45_508 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_518 ();
 DECAPx2_ASAP7_75t_R FILLER_45_543 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_549 ();
 FILLER_ASAP7_75t_R FILLER_45_559 ();
 DECAPx2_ASAP7_75t_R FILLER_45_567 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_573 ();
 DECAPx6_ASAP7_75t_R FILLER_45_585 ();
 DECAPx1_ASAP7_75t_R FILLER_45_599 ();
 DECAPx10_ASAP7_75t_R FILLER_45_610 ();
 DECAPx2_ASAP7_75t_R FILLER_45_639 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_645 ();
 DECAPx1_ASAP7_75t_R FILLER_45_654 ();
 FILLER_ASAP7_75t_R FILLER_45_665 ();
 DECAPx2_ASAP7_75t_R FILLER_45_677 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_683 ();
 DECAPx6_ASAP7_75t_R FILLER_45_692 ();
 FILLER_ASAP7_75t_R FILLER_45_706 ();
 DECAPx2_ASAP7_75t_R FILLER_45_711 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_717 ();
 DECAPx10_ASAP7_75t_R FILLER_45_727 ();
 DECAPx2_ASAP7_75t_R FILLER_45_749 ();
 FILLER_ASAP7_75t_R FILLER_45_761 ();
 DECAPx2_ASAP7_75t_R FILLER_45_777 ();
 FILLER_ASAP7_75t_R FILLER_45_790 ();
 DECAPx6_ASAP7_75t_R FILLER_45_800 ();
 DECAPx2_ASAP7_75t_R FILLER_45_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_820 ();
 DECAPx2_ASAP7_75t_R FILLER_45_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_837 ();
 DECAPx4_ASAP7_75t_R FILLER_45_852 ();
 DECAPx2_ASAP7_75t_R FILLER_45_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_876 ();
 DECAPx6_ASAP7_75t_R FILLER_45_883 ();
 DECAPx1_ASAP7_75t_R FILLER_45_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_901 ();
 DECAPx2_ASAP7_75t_R FILLER_45_911 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_917 ();
 FILLER_ASAP7_75t_R FILLER_45_923 ();
 FILLER_ASAP7_75t_R FILLER_45_927 ();
 DECAPx1_ASAP7_75t_R FILLER_45_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_939 ();
 DECAPx4_ASAP7_75t_R FILLER_45_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_953 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_962 ();
 DECAPx6_ASAP7_75t_R FILLER_45_968 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_982 ();
 DECAPx10_ASAP7_75t_R FILLER_45_988 ();
 DECAPx1_ASAP7_75t_R FILLER_45_1010 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_45_1027 ();
 FILLER_ASAP7_75t_R FILLER_45_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1083 ();
 FILLER_ASAP7_75t_R FILLER_45_1105 ();
 FILLER_ASAP7_75t_R FILLER_45_1133 ();
 FILLER_ASAP7_75t_R FILLER_45_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_45_1166 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_1172 ();
 DECAPx1_ASAP7_75t_R FILLER_45_1201 ();
 FILLER_ASAP7_75t_R FILLER_45_1208 ();
 FILLER_ASAP7_75t_R FILLER_45_1232 ();
 DECAPx2_ASAP7_75t_R FILLER_45_1256 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_45_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_45_1280 ();
 DECAPx6_ASAP7_75t_R FILLER_45_1305 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_1319 ();
 DECAPx1_ASAP7_75t_R FILLER_45_1348 ();
 DECAPx2_ASAP7_75t_R FILLER_45_1359 ();
 DECAPx2_ASAP7_75t_R FILLER_45_1368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_1374 ();
 DECAPx2_ASAP7_75t_R FILLER_46_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_8 ();
 FILLER_ASAP7_75t_R FILLER_46_15 ();
 DECAPx2_ASAP7_75t_R FILLER_46_20 ();
 FILLER_ASAP7_75t_R FILLER_46_26 ();
 DECAPx1_ASAP7_75t_R FILLER_46_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_35 ();
 DECAPx2_ASAP7_75t_R FILLER_46_44 ();
 FILLER_ASAP7_75t_R FILLER_46_50 ();
 DECAPx2_ASAP7_75t_R FILLER_46_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_66 ();
 DECAPx6_ASAP7_75t_R FILLER_46_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_107 ();
 DECAPx1_ASAP7_75t_R FILLER_46_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_118 ();
 FILLER_ASAP7_75t_R FILLER_46_145 ();
 DECAPx1_ASAP7_75t_R FILLER_46_154 ();
 FILLER_ASAP7_75t_R FILLER_46_164 ();
 DECAPx2_ASAP7_75t_R FILLER_46_173 ();
 FILLER_ASAP7_75t_R FILLER_46_189 ();
 FILLER_ASAP7_75t_R FILLER_46_199 ();
 FILLER_ASAP7_75t_R FILLER_46_207 ();
 FILLER_ASAP7_75t_R FILLER_46_215 ();
 DECAPx2_ASAP7_75t_R FILLER_46_220 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_46_226 ();
 DECAPx2_ASAP7_75t_R FILLER_46_232 ();
 FILLER_ASAP7_75t_R FILLER_46_238 ();
 DECAPx10_ASAP7_75t_R FILLER_46_243 ();
 DECAPx2_ASAP7_75t_R FILLER_46_265 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_46_271 ();
 DECAPx1_ASAP7_75t_R FILLER_46_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_284 ();
 FILLER_ASAP7_75t_R FILLER_46_291 ();
 FILLER_ASAP7_75t_R FILLER_46_300 ();
 FILLER_ASAP7_75t_R FILLER_46_309 ();
 DECAPx2_ASAP7_75t_R FILLER_46_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_324 ();
 DECAPx6_ASAP7_75t_R FILLER_46_331 ();
 DECAPx2_ASAP7_75t_R FILLER_46_351 ();
 DECAPx1_ASAP7_75t_R FILLER_46_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_367 ();
 DECAPx6_ASAP7_75t_R FILLER_46_371 ();
 FILLER_ASAP7_75t_R FILLER_46_391 ();
 FILLER_ASAP7_75t_R FILLER_46_399 ();
 DECAPx2_ASAP7_75t_R FILLER_46_404 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_46_410 ();
 DECAPx10_ASAP7_75t_R FILLER_46_421 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_46_443 ();
 DECAPx4_ASAP7_75t_R FILLER_46_452 ();
 FILLER_ASAP7_75t_R FILLER_46_464 ();
 DECAPx2_ASAP7_75t_R FILLER_46_472 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_46_478 ();
 FILLER_ASAP7_75t_R FILLER_46_507 ();
 DECAPx1_ASAP7_75t_R FILLER_46_515 ();
 DECAPx2_ASAP7_75t_R FILLER_46_525 ();
 FILLER_ASAP7_75t_R FILLER_46_531 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_46_540 ();
 DECAPx4_ASAP7_75t_R FILLER_46_549 ();
 DECAPx2_ASAP7_75t_R FILLER_46_569 ();
 FILLER_ASAP7_75t_R FILLER_46_575 ();
 DECAPx4_ASAP7_75t_R FILLER_46_585 ();
 FILLER_ASAP7_75t_R FILLER_46_595 ();
 DECAPx6_ASAP7_75t_R FILLER_46_607 ();
 DECAPx1_ASAP7_75t_R FILLER_46_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_625 ();
 FILLER_ASAP7_75t_R FILLER_46_632 ();
 FILLER_ASAP7_75t_R FILLER_46_644 ();
 DECAPx1_ASAP7_75t_R FILLER_46_654 ();
 FILLER_ASAP7_75t_R FILLER_46_664 ();
 FILLER_ASAP7_75t_R FILLER_46_672 ();
 DECAPx1_ASAP7_75t_R FILLER_46_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_686 ();
 DECAPx1_ASAP7_75t_R FILLER_46_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_699 ();
 FILLER_ASAP7_75t_R FILLER_46_706 ();
 DECAPx10_ASAP7_75t_R FILLER_46_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_736 ();
 DECAPx10_ASAP7_75t_R FILLER_46_744 ();
 DECAPx6_ASAP7_75t_R FILLER_46_766 ();
 DECAPx1_ASAP7_75t_R FILLER_46_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_784 ();
 FILLER_ASAP7_75t_R FILLER_46_791 ();
 DECAPx1_ASAP7_75t_R FILLER_46_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_803 ();
 DECAPx2_ASAP7_75t_R FILLER_46_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_818 ();
 FILLER_ASAP7_75t_R FILLER_46_829 ();
 FILLER_ASAP7_75t_R FILLER_46_837 ();
 FILLER_ASAP7_75t_R FILLER_46_848 ();
 DECAPx2_ASAP7_75t_R FILLER_46_856 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_46_862 ();
 FILLER_ASAP7_75t_R FILLER_46_872 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_46_880 ();
 FILLER_ASAP7_75t_R FILLER_46_886 ();
 FILLER_ASAP7_75t_R FILLER_46_897 ();
 FILLER_ASAP7_75t_R FILLER_46_905 ();
 DECAPx4_ASAP7_75t_R FILLER_46_913 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_46_923 ();
 FILLER_ASAP7_75t_R FILLER_46_952 ();
 FILLER_ASAP7_75t_R FILLER_46_980 ();
 DECAPx4_ASAP7_75t_R FILLER_46_985 ();
 DECAPx1_ASAP7_75t_R FILLER_46_1001 ();
 FILLER_ASAP7_75t_R FILLER_46_1008 ();
 FILLER_ASAP7_75t_R FILLER_46_1036 ();
 FILLER_ASAP7_75t_R FILLER_46_1048 ();
 DECAPx6_ASAP7_75t_R FILLER_46_1053 ();
 FILLER_ASAP7_75t_R FILLER_46_1075 ();
 FILLER_ASAP7_75t_R FILLER_46_1087 ();
 DECAPx4_ASAP7_75t_R FILLER_46_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_46_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1117 ();
 FILLER_ASAP7_75t_R FILLER_46_1121 ();
 FILLER_ASAP7_75t_R FILLER_46_1145 ();
 FILLER_ASAP7_75t_R FILLER_46_1154 ();
 FILLER_ASAP7_75t_R FILLER_46_1162 ();
 DECAPx4_ASAP7_75t_R FILLER_46_1167 ();
 FILLER_ASAP7_75t_R FILLER_46_1183 ();
 FILLER_ASAP7_75t_R FILLER_46_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_46_1193 ();
 FILLER_ASAP7_75t_R FILLER_46_1215 ();
 DECAPx4_ASAP7_75t_R FILLER_46_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1233 ();
 FILLER_ASAP7_75t_R FILLER_46_1246 ();
 FILLER_ASAP7_75t_R FILLER_46_1256 ();
 FILLER_ASAP7_75t_R FILLER_46_1264 ();
 DECAPx1_ASAP7_75t_R FILLER_46_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_46_1286 ();
 DECAPx1_ASAP7_75t_R FILLER_46_1299 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_1303 ();
 DECAPx1_ASAP7_75t_R FILLER_46_1307 ();
 DECAPx4_ASAP7_75t_R FILLER_46_1318 ();
 FILLER_ASAP7_75t_R FILLER_46_1328 ();
 FILLER_ASAP7_75t_R FILLER_46_1340 ();
 DECAPx1_ASAP7_75t_R FILLER_46_1345 ();
 FILLER_ASAP7_75t_R FILLER_46_1375 ();
 FILLER_ASAP7_75t_R FILLER_47_2 ();
 DECAPx2_ASAP7_75t_R FILLER_47_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_36 ();
 FILLER_ASAP7_75t_R FILLER_47_45 ();
 FILLER_ASAP7_75t_R FILLER_47_53 ();
 FILLER_ASAP7_75t_R FILLER_47_61 ();
 DECAPx2_ASAP7_75t_R FILLER_47_69 ();
 FILLER_ASAP7_75t_R FILLER_47_81 ();
 DECAPx6_ASAP7_75t_R FILLER_47_86 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_100 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_106 ();
 DECAPx2_ASAP7_75t_R FILLER_47_115 ();
 FILLER_ASAP7_75t_R FILLER_47_121 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_129 ();
 FILLER_ASAP7_75t_R FILLER_47_139 ();
 FILLER_ASAP7_75t_R FILLER_47_148 ();
 FILLER_ASAP7_75t_R FILLER_47_156 ();
 FILLER_ASAP7_75t_R FILLER_47_161 ();
 FILLER_ASAP7_75t_R FILLER_47_166 ();
 DECAPx2_ASAP7_75t_R FILLER_47_176 ();
 DECAPx2_ASAP7_75t_R FILLER_47_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_194 ();
 DECAPx4_ASAP7_75t_R FILLER_47_198 ();
 DECAPx2_ASAP7_75t_R FILLER_47_214 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_220 ();
 DECAPx10_ASAP7_75t_R FILLER_47_229 ();
 DECAPx10_ASAP7_75t_R FILLER_47_251 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_273 ();
 FILLER_ASAP7_75t_R FILLER_47_279 ();
 DECAPx1_ASAP7_75t_R FILLER_47_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_311 ();
 DECAPx1_ASAP7_75t_R FILLER_47_338 ();
 DECAPx6_ASAP7_75t_R FILLER_47_357 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_371 ();
 DECAPx2_ASAP7_75t_R FILLER_47_380 ();
 FILLER_ASAP7_75t_R FILLER_47_386 ();
 FILLER_ASAP7_75t_R FILLER_47_391 ();
 DECAPx1_ASAP7_75t_R FILLER_47_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_404 ();
 FILLER_ASAP7_75t_R FILLER_47_411 ();
 FILLER_ASAP7_75t_R FILLER_47_421 ();
 DECAPx2_ASAP7_75t_R FILLER_47_429 ();
 FILLER_ASAP7_75t_R FILLER_47_435 ();
 FILLER_ASAP7_75t_R FILLER_47_452 ();
 FILLER_ASAP7_75t_R FILLER_47_457 ();
 FILLER_ASAP7_75t_R FILLER_47_485 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_493 ();
 DECAPx2_ASAP7_75t_R FILLER_47_499 ();
 DECAPx2_ASAP7_75t_R FILLER_47_511 ();
 DECAPx2_ASAP7_75t_R FILLER_47_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_529 ();
 DECAPx1_ASAP7_75t_R FILLER_47_550 ();
 FILLER_ASAP7_75t_R FILLER_47_561 ();
 DECAPx10_ASAP7_75t_R FILLER_47_571 ();
 DECAPx2_ASAP7_75t_R FILLER_47_593 ();
 DECAPx6_ASAP7_75t_R FILLER_47_605 ();
 DECAPx1_ASAP7_75t_R FILLER_47_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_623 ();
 FILLER_ASAP7_75t_R FILLER_47_632 ();
 DECAPx10_ASAP7_75t_R FILLER_47_640 ();
 DECAPx2_ASAP7_75t_R FILLER_47_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_668 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_675 ();
 DECAPx6_ASAP7_75t_R FILLER_47_686 ();
 DECAPx2_ASAP7_75t_R FILLER_47_708 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_714 ();
 FILLER_ASAP7_75t_R FILLER_47_737 ();
 DECAPx2_ASAP7_75t_R FILLER_47_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_765 ();
 DECAPx2_ASAP7_75t_R FILLER_47_773 ();
 FILLER_ASAP7_75t_R FILLER_47_779 ();
 FILLER_ASAP7_75t_R FILLER_47_787 ();
 DECAPx4_ASAP7_75t_R FILLER_47_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_805 ();
 FILLER_ASAP7_75t_R FILLER_47_812 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_817 ();
 FILLER_ASAP7_75t_R FILLER_47_826 ();
 DECAPx2_ASAP7_75t_R FILLER_47_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_840 ();
 DECAPx4_ASAP7_75t_R FILLER_47_848 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_858 ();
 DECAPx6_ASAP7_75t_R FILLER_47_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_889 ();
 DECAPx2_ASAP7_75t_R FILLER_47_896 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_902 ();
 DECAPx1_ASAP7_75t_R FILLER_47_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_912 ();
 FILLER_ASAP7_75t_R FILLER_47_923 ();
 DECAPx10_ASAP7_75t_R FILLER_47_927 ();
 DECAPx6_ASAP7_75t_R FILLER_47_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_963 ();
 FILLER_ASAP7_75t_R FILLER_47_990 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1027 ();
 DECAPx4_ASAP7_75t_R FILLER_47_1049 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1114 ();
 FILLER_ASAP7_75t_R FILLER_47_1120 ();
 DECAPx6_ASAP7_75t_R FILLER_47_1128 ();
 DECAPx1_ASAP7_75t_R FILLER_47_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_47_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1190 ();
 DECAPx6_ASAP7_75t_R FILLER_47_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1243 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_1249 ();
 DECAPx4_ASAP7_75t_R FILLER_47_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1288 ();
 FILLER_ASAP7_75t_R FILLER_47_1315 ();
 DECAPx2_ASAP7_75t_R FILLER_47_1343 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_1349 ();
 DECAPx6_ASAP7_75t_R FILLER_47_1358 ();
 DECAPx1_ASAP7_75t_R FILLER_47_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_1376 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_2 ();
 FILLER_ASAP7_75t_R FILLER_48_11 ();
 FILLER_ASAP7_75t_R FILLER_48_19 ();
 DECAPx4_ASAP7_75t_R FILLER_48_24 ();
 FILLER_ASAP7_75t_R FILLER_48_40 ();
 DECAPx2_ASAP7_75t_R FILLER_48_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_54 ();
 DECAPx6_ASAP7_75t_R FILLER_48_61 ();
 FILLER_ASAP7_75t_R FILLER_48_83 ();
 DECAPx1_ASAP7_75t_R FILLER_48_91 ();
 DECAPx1_ASAP7_75t_R FILLER_48_101 ();
 FILLER_ASAP7_75t_R FILLER_48_131 ();
 FILLER_ASAP7_75t_R FILLER_48_136 ();
 DECAPx2_ASAP7_75t_R FILLER_48_141 ();
 FILLER_ASAP7_75t_R FILLER_48_147 ();
 DECAPx2_ASAP7_75t_R FILLER_48_155 ();
 DECAPx4_ASAP7_75t_R FILLER_48_167 ();
 DECAPx4_ASAP7_75t_R FILLER_48_192 ();
 FILLER_ASAP7_75t_R FILLER_48_202 ();
 DECAPx2_ASAP7_75t_R FILLER_48_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_236 ();
 FILLER_ASAP7_75t_R FILLER_48_263 ();
 DECAPx4_ASAP7_75t_R FILLER_48_273 ();
 FILLER_ASAP7_75t_R FILLER_48_283 ();
 DECAPx1_ASAP7_75t_R FILLER_48_291 ();
 DECAPx2_ASAP7_75t_R FILLER_48_298 ();
 DECAPx4_ASAP7_75t_R FILLER_48_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_317 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_324 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_330 ();
 DECAPx2_ASAP7_75t_R FILLER_48_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_342 ();
 DECAPx6_ASAP7_75t_R FILLER_48_349 ();
 FILLER_ASAP7_75t_R FILLER_48_363 ();
 FILLER_ASAP7_75t_R FILLER_48_371 ();
 FILLER_ASAP7_75t_R FILLER_48_399 ();
 DECAPx6_ASAP7_75t_R FILLER_48_423 ();
 DECAPx6_ASAP7_75t_R FILLER_48_444 ();
 DECAPx1_ASAP7_75t_R FILLER_48_458 ();
 FILLER_ASAP7_75t_R FILLER_48_464 ();
 FILLER_ASAP7_75t_R FILLER_48_472 ();
 DECAPx10_ASAP7_75t_R FILLER_48_477 ();
 DECAPx1_ASAP7_75t_R FILLER_48_499 ();
 DECAPx10_ASAP7_75t_R FILLER_48_529 ();
 DECAPx1_ASAP7_75t_R FILLER_48_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_555 ();
 DECAPx1_ASAP7_75t_R FILLER_48_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_566 ();
 FILLER_ASAP7_75t_R FILLER_48_573 ();
 FILLER_ASAP7_75t_R FILLER_48_583 ();
 DECAPx4_ASAP7_75t_R FILLER_48_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_601 ();
 DECAPx2_ASAP7_75t_R FILLER_48_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_614 ();
 DECAPx10_ASAP7_75t_R FILLER_48_621 ();
 DECAPx1_ASAP7_75t_R FILLER_48_643 ();
 FILLER_ASAP7_75t_R FILLER_48_655 ();
 DECAPx2_ASAP7_75t_R FILLER_48_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_669 ();
 DECAPx6_ASAP7_75t_R FILLER_48_678 ();
 DECAPx2_ASAP7_75t_R FILLER_48_692 ();
 FILLER_ASAP7_75t_R FILLER_48_707 ();
 FILLER_ASAP7_75t_R FILLER_48_719 ();
 DECAPx4_ASAP7_75t_R FILLER_48_728 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_738 ();
 DECAPx2_ASAP7_75t_R FILLER_48_747 ();
 FILLER_ASAP7_75t_R FILLER_48_753 ();
 DECAPx1_ASAP7_75t_R FILLER_48_759 ();
 FILLER_ASAP7_75t_R FILLER_48_783 ();
 DECAPx10_ASAP7_75t_R FILLER_48_793 ();
 DECAPx2_ASAP7_75t_R FILLER_48_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_821 ();
 DECAPx4_ASAP7_75t_R FILLER_48_832 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_842 ();
 DECAPx6_ASAP7_75t_R FILLER_48_851 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_872 ();
 DECAPx2_ASAP7_75t_R FILLER_48_881 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_887 ();
 DECAPx10_ASAP7_75t_R FILLER_48_896 ();
 FILLER_ASAP7_75t_R FILLER_48_918 ();
 FILLER_ASAP7_75t_R FILLER_48_927 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_935 ();
 DECAPx4_ASAP7_75t_R FILLER_48_948 ();
 FILLER_ASAP7_75t_R FILLER_48_958 ();
 DECAPx2_ASAP7_75t_R FILLER_48_970 ();
 FILLER_ASAP7_75t_R FILLER_48_979 ();
 DECAPx2_ASAP7_75t_R FILLER_48_991 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_997 ();
 DECAPx6_ASAP7_75t_R FILLER_48_1003 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1017 ();
 DECAPx4_ASAP7_75t_R FILLER_48_1028 ();
 FILLER_ASAP7_75t_R FILLER_48_1038 ();
 DECAPx6_ASAP7_75t_R FILLER_48_1049 ();
 FILLER_ASAP7_75t_R FILLER_48_1063 ();
 FILLER_ASAP7_75t_R FILLER_48_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1080 ();
 FILLER_ASAP7_75t_R FILLER_48_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1098 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_1105 ();
 DECAPx4_ASAP7_75t_R FILLER_48_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1144 ();
 FILLER_ASAP7_75t_R FILLER_48_1148 ();
 FILLER_ASAP7_75t_R FILLER_48_1176 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1193 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_1220 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1230 ();
 DECAPx1_ASAP7_75t_R FILLER_48_1234 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1248 ();
 DECAPx6_ASAP7_75t_R FILLER_48_1261 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1275 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1289 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_1295 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1304 ();
 FILLER_ASAP7_75t_R FILLER_48_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1318 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_48_1328 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_1350 ();
 FILLER_ASAP7_75t_R FILLER_48_1360 ();
 DECAPx2_ASAP7_75t_R FILLER_48_1368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_1374 ();
 DECAPx6_ASAP7_75t_R FILLER_49_2 ();
 DECAPx2_ASAP7_75t_R FILLER_49_16 ();
 DECAPx10_ASAP7_75t_R FILLER_49_28 ();
 DECAPx4_ASAP7_75t_R FILLER_49_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_60 ();
 DECAPx2_ASAP7_75t_R FILLER_49_67 ();
 FILLER_ASAP7_75t_R FILLER_49_73 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_89 ();
 DECAPx2_ASAP7_75t_R FILLER_49_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_113 ();
 DECAPx1_ASAP7_75t_R FILLER_49_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_124 ();
 DECAPx6_ASAP7_75t_R FILLER_49_128 ();
 FILLER_ASAP7_75t_R FILLER_49_142 ();
 DECAPx6_ASAP7_75t_R FILLER_49_170 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_184 ();
 DECAPx2_ASAP7_75t_R FILLER_49_193 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_199 ();
 DECAPx4_ASAP7_75t_R FILLER_49_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_218 ();
 DECAPx2_ASAP7_75t_R FILLER_49_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_228 ();
 DECAPx2_ASAP7_75t_R FILLER_49_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_238 ();
 FILLER_ASAP7_75t_R FILLER_49_245 ();
 DECAPx1_ASAP7_75t_R FILLER_49_253 ();
 FILLER_ASAP7_75t_R FILLER_49_263 ();
 FILLER_ASAP7_75t_R FILLER_49_273 ();
 DECAPx2_ASAP7_75t_R FILLER_49_281 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_287 ();
 DECAPx6_ASAP7_75t_R FILLER_49_296 ();
 DECAPx4_ASAP7_75t_R FILLER_49_318 ();
 FILLER_ASAP7_75t_R FILLER_49_334 ();
 DECAPx2_ASAP7_75t_R FILLER_49_344 ();
 FILLER_ASAP7_75t_R FILLER_49_350 ();
 FILLER_ASAP7_75t_R FILLER_49_360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_368 ();
 FILLER_ASAP7_75t_R FILLER_49_397 ();
 FILLER_ASAP7_75t_R FILLER_49_406 ();
 FILLER_ASAP7_75t_R FILLER_49_411 ();
 FILLER_ASAP7_75t_R FILLER_49_421 ();
 FILLER_ASAP7_75t_R FILLER_49_429 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_437 ();
 DECAPx10_ASAP7_75t_R FILLER_49_451 ();
 DECAPx6_ASAP7_75t_R FILLER_49_473 ();
 DECAPx10_ASAP7_75t_R FILLER_49_493 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_515 ();
 DECAPx10_ASAP7_75t_R FILLER_49_521 ();
 DECAPx4_ASAP7_75t_R FILLER_49_543 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_553 ();
 FILLER_ASAP7_75t_R FILLER_49_562 ();
 DECAPx4_ASAP7_75t_R FILLER_49_570 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_580 ();
 DECAPx2_ASAP7_75t_R FILLER_49_591 ();
 FILLER_ASAP7_75t_R FILLER_49_604 ();
 FILLER_ASAP7_75t_R FILLER_49_613 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_621 ();
 DECAPx1_ASAP7_75t_R FILLER_49_630 ();
 DECAPx10_ASAP7_75t_R FILLER_49_640 ();
 DECAPx10_ASAP7_75t_R FILLER_49_662 ();
 DECAPx2_ASAP7_75t_R FILLER_49_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_690 ();
 FILLER_ASAP7_75t_R FILLER_49_697 ();
 DECAPx6_ASAP7_75t_R FILLER_49_705 ();
 DECAPx2_ASAP7_75t_R FILLER_49_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_725 ();
 DECAPx10_ASAP7_75t_R FILLER_49_733 ();
 DECAPx10_ASAP7_75t_R FILLER_49_755 ();
 DECAPx2_ASAP7_75t_R FILLER_49_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_783 ();
 DECAPx2_ASAP7_75t_R FILLER_49_792 ();
 FILLER_ASAP7_75t_R FILLER_49_798 ();
 DECAPx10_ASAP7_75t_R FILLER_49_806 ();
 DECAPx2_ASAP7_75t_R FILLER_49_828 ();
 FILLER_ASAP7_75t_R FILLER_49_834 ();
 DECAPx2_ASAP7_75t_R FILLER_49_846 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_852 ();
 FILLER_ASAP7_75t_R FILLER_49_863 ();
 DECAPx1_ASAP7_75t_R FILLER_49_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_872 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_879 ();
 FILLER_ASAP7_75t_R FILLER_49_892 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_902 ();
 FILLER_ASAP7_75t_R FILLER_49_914 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_922 ();
 DECAPx2_ASAP7_75t_R FILLER_49_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_933 ();
 DECAPx2_ASAP7_75t_R FILLER_49_942 ();
 DECAPx10_ASAP7_75t_R FILLER_49_974 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_996 ();
 FILLER_ASAP7_75t_R FILLER_49_1007 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_1017 ();
 FILLER_ASAP7_75t_R FILLER_49_1040 ();
 FILLER_ASAP7_75t_R FILLER_49_1048 ();
 FILLER_ASAP7_75t_R FILLER_49_1056 ();
 FILLER_ASAP7_75t_R FILLER_49_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_49_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1077 ();
 DECAPx6_ASAP7_75t_R FILLER_49_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_1113 ();
 FILLER_ASAP7_75t_R FILLER_49_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_49_1126 ();
 DECAPx4_ASAP7_75t_R FILLER_49_1156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_1166 ();
 FILLER_ASAP7_75t_R FILLER_49_1172 ();
 FILLER_ASAP7_75t_R FILLER_49_1200 ();
 FILLER_ASAP7_75t_R FILLER_49_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1213 ();
 DECAPx6_ASAP7_75t_R FILLER_49_1235 ();
 DECAPx2_ASAP7_75t_R FILLER_49_1249 ();
 DECAPx6_ASAP7_75t_R FILLER_49_1265 ();
 DECAPx1_ASAP7_75t_R FILLER_49_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_49_1313 ();
 FILLER_ASAP7_75t_R FILLER_49_1347 ();
 FILLER_ASAP7_75t_R FILLER_49_1375 ();
 DECAPx1_ASAP7_75t_R FILLER_50_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_6 ();
 DECAPx1_ASAP7_75t_R FILLER_50_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_17 ();
 DECAPx4_ASAP7_75t_R FILLER_50_44 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_54 ();
 DECAPx10_ASAP7_75t_R FILLER_50_83 ();
 DECAPx2_ASAP7_75t_R FILLER_50_105 ();
 FILLER_ASAP7_75t_R FILLER_50_137 ();
 FILLER_ASAP7_75t_R FILLER_50_145 ();
 DECAPx2_ASAP7_75t_R FILLER_50_150 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_156 ();
 DECAPx2_ASAP7_75t_R FILLER_50_162 ();
 DECAPx4_ASAP7_75t_R FILLER_50_171 ();
 FILLER_ASAP7_75t_R FILLER_50_181 ();
 DECAPx2_ASAP7_75t_R FILLER_50_191 ();
 FILLER_ASAP7_75t_R FILLER_50_197 ();
 DECAPx1_ASAP7_75t_R FILLER_50_225 ();
 DECAPx6_ASAP7_75t_R FILLER_50_235 ();
 FILLER_ASAP7_75t_R FILLER_50_249 ();
 DECAPx2_ASAP7_75t_R FILLER_50_254 ();
 DECAPx2_ASAP7_75t_R FILLER_50_263 ();
 DECAPx2_ASAP7_75t_R FILLER_50_275 ();
 FILLER_ASAP7_75t_R FILLER_50_281 ();
 FILLER_ASAP7_75t_R FILLER_50_309 ();
 DECAPx6_ASAP7_75t_R FILLER_50_318 ();
 FILLER_ASAP7_75t_R FILLER_50_332 ();
 DECAPx6_ASAP7_75t_R FILLER_50_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_354 ();
 DECAPx4_ASAP7_75t_R FILLER_50_366 ();
 DECAPx1_ASAP7_75t_R FILLER_50_382 ();
 DECAPx1_ASAP7_75t_R FILLER_50_389 ();
 FILLER_ASAP7_75t_R FILLER_50_400 ();
 DECAPx1_ASAP7_75t_R FILLER_50_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_413 ();
 DECAPx2_ASAP7_75t_R FILLER_50_422 ();
 FILLER_ASAP7_75t_R FILLER_50_428 ();
 FILLER_ASAP7_75t_R FILLER_50_436 ();
 FILLER_ASAP7_75t_R FILLER_50_460 ();
 FILLER_ASAP7_75t_R FILLER_50_464 ();
 FILLER_ASAP7_75t_R FILLER_50_469 ();
 FILLER_ASAP7_75t_R FILLER_50_477 ();
 DECAPx2_ASAP7_75t_R FILLER_50_505 ();
 FILLER_ASAP7_75t_R FILLER_50_511 ();
 FILLER_ASAP7_75t_R FILLER_50_519 ();
 DECAPx4_ASAP7_75t_R FILLER_50_539 ();
 FILLER_ASAP7_75t_R FILLER_50_549 ();
 DECAPx1_ASAP7_75t_R FILLER_50_558 ();
 DECAPx2_ASAP7_75t_R FILLER_50_570 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_576 ();
 DECAPx4_ASAP7_75t_R FILLER_50_585 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_595 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_605 ();
 DECAPx6_ASAP7_75t_R FILLER_50_615 ();
 DECAPx1_ASAP7_75t_R FILLER_50_629 ();
 DECAPx1_ASAP7_75t_R FILLER_50_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_643 ();
 FILLER_ASAP7_75t_R FILLER_50_650 ();
 DECAPx4_ASAP7_75t_R FILLER_50_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_670 ();
 DECAPx4_ASAP7_75t_R FILLER_50_677 ();
 DECAPx10_ASAP7_75t_R FILLER_50_694 ();
 DECAPx4_ASAP7_75t_R FILLER_50_716 ();
 FILLER_ASAP7_75t_R FILLER_50_746 ();
 DECAPx4_ASAP7_75t_R FILLER_50_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_764 ();
 DECAPx4_ASAP7_75t_R FILLER_50_771 ();
 FILLER_ASAP7_75t_R FILLER_50_781 ();
 DECAPx6_ASAP7_75t_R FILLER_50_789 ();
 FILLER_ASAP7_75t_R FILLER_50_810 ();
 FILLER_ASAP7_75t_R FILLER_50_818 ();
 FILLER_ASAP7_75t_R FILLER_50_826 ();
 DECAPx2_ASAP7_75t_R FILLER_50_834 ();
 DECAPx4_ASAP7_75t_R FILLER_50_862 ();
 DECAPx4_ASAP7_75t_R FILLER_50_881 ();
 FILLER_ASAP7_75t_R FILLER_50_913 ();
 DECAPx4_ASAP7_75t_R FILLER_50_921 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_931 ();
 DECAPx1_ASAP7_75t_R FILLER_50_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_941 ();
 DECAPx2_ASAP7_75t_R FILLER_50_949 ();
 FILLER_ASAP7_75t_R FILLER_50_963 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_968 ();
 DECAPx2_ASAP7_75t_R FILLER_50_981 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_987 ();
 FILLER_ASAP7_75t_R FILLER_50_993 ();
 DECAPx2_ASAP7_75t_R FILLER_50_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1016 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1025 ();
 DECAPx6_ASAP7_75t_R FILLER_50_1032 ();
 FILLER_ASAP7_75t_R FILLER_50_1046 ();
 FILLER_ASAP7_75t_R FILLER_50_1074 ();
 DECAPx4_ASAP7_75t_R FILLER_50_1082 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_1092 ();
 DECAPx6_ASAP7_75t_R FILLER_50_1121 ();
 FILLER_ASAP7_75t_R FILLER_50_1135 ();
 FILLER_ASAP7_75t_R FILLER_50_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1150 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_50_1191 ();
 FILLER_ASAP7_75t_R FILLER_50_1221 ();
 DECAPx1_ASAP7_75t_R FILLER_50_1231 ();
 FILLER_ASAP7_75t_R FILLER_50_1261 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1289 ();
 DECAPx4_ASAP7_75t_R FILLER_50_1307 ();
 DECAPx4_ASAP7_75t_R FILLER_50_1343 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1360 ();
 DECAPx2_ASAP7_75t_R FILLER_50_1369 ();
 FILLER_ASAP7_75t_R FILLER_50_1375 ();
 FILLER_ASAP7_75t_R FILLER_51_2 ();
 FILLER_ASAP7_75t_R FILLER_51_30 ();
 FILLER_ASAP7_75t_R FILLER_51_35 ();
 FILLER_ASAP7_75t_R FILLER_51_43 ();
 DECAPx2_ASAP7_75t_R FILLER_51_51 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_57 ();
 DECAPx2_ASAP7_75t_R FILLER_51_66 ();
 DECAPx10_ASAP7_75t_R FILLER_51_75 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_97 ();
 DECAPx2_ASAP7_75t_R FILLER_51_110 ();
 FILLER_ASAP7_75t_R FILLER_51_116 ();
 DECAPx2_ASAP7_75t_R FILLER_51_124 ();
 DECAPx10_ASAP7_75t_R FILLER_51_156 ();
 DECAPx2_ASAP7_75t_R FILLER_51_178 ();
 DECAPx4_ASAP7_75t_R FILLER_51_195 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_211 ();
 DECAPx2_ASAP7_75t_R FILLER_51_217 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_223 ();
 FILLER_ASAP7_75t_R FILLER_51_232 ();
 DECAPx6_ASAP7_75t_R FILLER_51_242 ();
 DECAPx2_ASAP7_75t_R FILLER_51_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_262 ();
 DECAPx6_ASAP7_75t_R FILLER_51_269 ();
 DECAPx1_ASAP7_75t_R FILLER_51_283 ();
 DECAPx1_ASAP7_75t_R FILLER_51_293 ();
 DECAPx1_ASAP7_75t_R FILLER_51_300 ();
 FILLER_ASAP7_75t_R FILLER_51_310 ();
 DECAPx2_ASAP7_75t_R FILLER_51_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_324 ();
 FILLER_ASAP7_75t_R FILLER_51_331 ();
 DECAPx10_ASAP7_75t_R FILLER_51_336 ();
 DECAPx10_ASAP7_75t_R FILLER_51_358 ();
 DECAPx1_ASAP7_75t_R FILLER_51_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_384 ();
 FILLER_ASAP7_75t_R FILLER_51_391 ();
 DECAPx2_ASAP7_75t_R FILLER_51_400 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_406 ();
 DECAPx6_ASAP7_75t_R FILLER_51_415 ();
 DECAPx2_ASAP7_75t_R FILLER_51_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_435 ();
 DECAPx2_ASAP7_75t_R FILLER_51_444 ();
 DECAPx2_ASAP7_75t_R FILLER_51_476 ();
 FILLER_ASAP7_75t_R FILLER_51_482 ();
 DECAPx1_ASAP7_75t_R FILLER_51_490 ();
 DECAPx1_ASAP7_75t_R FILLER_51_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_501 ();
 FILLER_ASAP7_75t_R FILLER_51_505 ();
 FILLER_ASAP7_75t_R FILLER_51_513 ();
 DECAPx1_ASAP7_75t_R FILLER_51_523 ();
 FILLER_ASAP7_75t_R FILLER_51_547 ();
 DECAPx6_ASAP7_75t_R FILLER_51_571 ();
 DECAPx2_ASAP7_75t_R FILLER_51_588 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_604 ();
 DECAPx4_ASAP7_75t_R FILLER_51_610 ();
 FILLER_ASAP7_75t_R FILLER_51_626 ();
 FILLER_ASAP7_75t_R FILLER_51_634 ();
 FILLER_ASAP7_75t_R FILLER_51_643 ();
 FILLER_ASAP7_75t_R FILLER_51_648 ();
 DECAPx2_ASAP7_75t_R FILLER_51_660 ();
 DECAPx2_ASAP7_75t_R FILLER_51_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_679 ();
 DECAPx1_ASAP7_75t_R FILLER_51_690 ();
 FILLER_ASAP7_75t_R FILLER_51_701 ();
 DECAPx2_ASAP7_75t_R FILLER_51_723 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_729 ();
 DECAPx2_ASAP7_75t_R FILLER_51_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_744 ();
 FILLER_ASAP7_75t_R FILLER_51_765 ();
 FILLER_ASAP7_75t_R FILLER_51_773 ();
 DECAPx6_ASAP7_75t_R FILLER_51_778 ();
 FILLER_ASAP7_75t_R FILLER_51_792 ();
 FILLER_ASAP7_75t_R FILLER_51_801 ();
 DECAPx2_ASAP7_75t_R FILLER_51_809 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_822 ();
 DECAPx2_ASAP7_75t_R FILLER_51_828 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_834 ();
 DECAPx2_ASAP7_75t_R FILLER_51_843 ();
 FILLER_ASAP7_75t_R FILLER_51_849 ();
 DECAPx6_ASAP7_75t_R FILLER_51_858 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_872 ();
 DECAPx4_ASAP7_75t_R FILLER_51_881 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_891 ();
 DECAPx4_ASAP7_75t_R FILLER_51_902 ();
 DECAPx1_ASAP7_75t_R FILLER_51_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_924 ();
 FILLER_ASAP7_75t_R FILLER_51_927 ();
 FILLER_ASAP7_75t_R FILLER_51_955 ();
 DECAPx6_ASAP7_75t_R FILLER_51_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_974 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1016 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1051 ();
 FILLER_ASAP7_75t_R FILLER_51_1055 ();
 DECAPx4_ASAP7_75t_R FILLER_51_1064 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1107 ();
 FILLER_ASAP7_75t_R FILLER_51_1111 ();
 FILLER_ASAP7_75t_R FILLER_51_1120 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_51_1141 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1163 ();
 FILLER_ASAP7_75t_R FILLER_51_1175 ();
 DECAPx4_ASAP7_75t_R FILLER_51_1184 ();
 FILLER_ASAP7_75t_R FILLER_51_1194 ();
 FILLER_ASAP7_75t_R FILLER_51_1208 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1213 ();
 FILLER_ASAP7_75t_R FILLER_51_1243 ();
 FILLER_ASAP7_75t_R FILLER_51_1253 ();
 DECAPx1_ASAP7_75t_R FILLER_51_1258 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1266 ();
 DECAPx6_ASAP7_75t_R FILLER_51_1298 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_1312 ();
 DECAPx2_ASAP7_75t_R FILLER_51_1323 ();
 FILLER_ASAP7_75t_R FILLER_51_1329 ();
 FILLER_ASAP7_75t_R FILLER_51_1334 ();
 DECAPx4_ASAP7_75t_R FILLER_51_1339 ();
 FILLER_ASAP7_75t_R FILLER_51_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_52_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_8 ();
 FILLER_ASAP7_75t_R FILLER_52_17 ();
 DECAPx4_ASAP7_75t_R FILLER_52_22 ();
 DECAPx4_ASAP7_75t_R FILLER_52_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_48 ();
 DECAPx1_ASAP7_75t_R FILLER_52_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_59 ();
 DECAPx6_ASAP7_75t_R FILLER_52_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_80 ();
 DECAPx2_ASAP7_75t_R FILLER_52_89 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_95 ();
 FILLER_ASAP7_75t_R FILLER_52_136 ();
 FILLER_ASAP7_75t_R FILLER_52_144 ();
 DECAPx1_ASAP7_75t_R FILLER_52_149 ();
 FILLER_ASAP7_75t_R FILLER_52_159 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_169 ();
 FILLER_ASAP7_75t_R FILLER_52_180 ();
 DECAPx6_ASAP7_75t_R FILLER_52_188 ();
 DECAPx2_ASAP7_75t_R FILLER_52_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_208 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_215 ();
 DECAPx4_ASAP7_75t_R FILLER_52_224 ();
 DECAPx1_ASAP7_75t_R FILLER_52_242 ();
 DECAPx10_ASAP7_75t_R FILLER_52_252 ();
 DECAPx10_ASAP7_75t_R FILLER_52_274 ();
 DECAPx6_ASAP7_75t_R FILLER_52_296 ();
 DECAPx1_ASAP7_75t_R FILLER_52_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_314 ();
 DECAPx2_ASAP7_75t_R FILLER_52_341 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_347 ();
 DECAPx1_ASAP7_75t_R FILLER_52_356 ();
 DECAPx2_ASAP7_75t_R FILLER_52_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_372 ();
 FILLER_ASAP7_75t_R FILLER_52_399 ();
 FILLER_ASAP7_75t_R FILLER_52_407 ();
 FILLER_ASAP7_75t_R FILLER_52_415 ();
 DECAPx2_ASAP7_75t_R FILLER_52_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_429 ();
 DECAPx6_ASAP7_75t_R FILLER_52_433 ();
 DECAPx2_ASAP7_75t_R FILLER_52_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_453 ();
 FILLER_ASAP7_75t_R FILLER_52_460 ();
 FILLER_ASAP7_75t_R FILLER_52_464 ();
 FILLER_ASAP7_75t_R FILLER_52_472 ();
 DECAPx2_ASAP7_75t_R FILLER_52_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_506 ();
 FILLER_ASAP7_75t_R FILLER_52_513 ();
 DECAPx2_ASAP7_75t_R FILLER_52_523 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_529 ();
 FILLER_ASAP7_75t_R FILLER_52_550 ();
 FILLER_ASAP7_75t_R FILLER_52_561 ();
 DECAPx4_ASAP7_75t_R FILLER_52_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_579 ();
 FILLER_ASAP7_75t_R FILLER_52_588 ();
 DECAPx1_ASAP7_75t_R FILLER_52_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_601 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_612 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_623 ();
 DECAPx4_ASAP7_75t_R FILLER_52_632 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_642 ();
 FILLER_ASAP7_75t_R FILLER_52_651 ();
 DECAPx1_ASAP7_75t_R FILLER_52_660 ();
 FILLER_ASAP7_75t_R FILLER_52_670 ();
 DECAPx2_ASAP7_75t_R FILLER_52_678 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_684 ();
 FILLER_ASAP7_75t_R FILLER_52_697 ();
 DECAPx2_ASAP7_75t_R FILLER_52_709 ();
 FILLER_ASAP7_75t_R FILLER_52_715 ();
 DECAPx6_ASAP7_75t_R FILLER_52_724 ();
 DECAPx1_ASAP7_75t_R FILLER_52_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_742 ();
 FILLER_ASAP7_75t_R FILLER_52_767 ();
 FILLER_ASAP7_75t_R FILLER_52_773 ();
 FILLER_ASAP7_75t_R FILLER_52_778 ();
 FILLER_ASAP7_75t_R FILLER_52_788 ();
 FILLER_ASAP7_75t_R FILLER_52_798 ();
 FILLER_ASAP7_75t_R FILLER_52_808 ();
 DECAPx2_ASAP7_75t_R FILLER_52_816 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_822 ();
 DECAPx4_ASAP7_75t_R FILLER_52_832 ();
 FILLER_ASAP7_75t_R FILLER_52_849 ();
 FILLER_ASAP7_75t_R FILLER_52_859 ();
 FILLER_ASAP7_75t_R FILLER_52_867 ();
 DECAPx1_ASAP7_75t_R FILLER_52_875 ();
 DECAPx2_ASAP7_75t_R FILLER_52_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_892 ();
 DECAPx4_ASAP7_75t_R FILLER_52_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_909 ();
 DECAPx2_ASAP7_75t_R FILLER_52_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_919 ();
 FILLER_ASAP7_75t_R FILLER_52_926 ();
 DECAPx2_ASAP7_75t_R FILLER_52_934 ();
 FILLER_ASAP7_75t_R FILLER_52_940 ();
 DECAPx4_ASAP7_75t_R FILLER_52_950 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_960 ();
 DECAPx4_ASAP7_75t_R FILLER_52_969 ();
 FILLER_ASAP7_75t_R FILLER_52_979 ();
 FILLER_ASAP7_75t_R FILLER_52_985 ();
 DECAPx1_ASAP7_75t_R FILLER_52_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1042 ();
 DECAPx4_ASAP7_75t_R FILLER_52_1064 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_1084 ();
 FILLER_ASAP7_75t_R FILLER_52_1090 ();
 DECAPx4_ASAP7_75t_R FILLER_52_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1185 ();
 DECAPx6_ASAP7_75t_R FILLER_52_1201 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_1215 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_1228 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_52_1243 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1265 ();
 FILLER_ASAP7_75t_R FILLER_52_1271 ();
 FILLER_ASAP7_75t_R FILLER_52_1279 ();
 FILLER_ASAP7_75t_R FILLER_52_1284 ();
 FILLER_ASAP7_75t_R FILLER_52_1289 ();
 DECAPx1_ASAP7_75t_R FILLER_52_1294 ();
 FILLER_ASAP7_75t_R FILLER_52_1324 ();
 DECAPx1_ASAP7_75t_R FILLER_52_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1333 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1346 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_1352 ();
 DECAPx1_ASAP7_75t_R FILLER_52_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_1365 ();
 DECAPx2_ASAP7_75t_R FILLER_52_1369 ();
 FILLER_ASAP7_75t_R FILLER_52_1375 ();
 DECAPx4_ASAP7_75t_R FILLER_53_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_12 ();
 DECAPx6_ASAP7_75t_R FILLER_53_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_33 ();
 DECAPx1_ASAP7_75t_R FILLER_53_37 ();
 FILLER_ASAP7_75t_R FILLER_53_49 ();
 DECAPx2_ASAP7_75t_R FILLER_53_57 ();
 FILLER_ASAP7_75t_R FILLER_53_63 ();
 DECAPx6_ASAP7_75t_R FILLER_53_71 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_85 ();
 FILLER_ASAP7_75t_R FILLER_53_96 ();
 DECAPx2_ASAP7_75t_R FILLER_53_105 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_111 ();
 DECAPx10_ASAP7_75t_R FILLER_53_120 ();
 DECAPx6_ASAP7_75t_R FILLER_53_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_156 ();
 DECAPx2_ASAP7_75t_R FILLER_53_165 ();
 FILLER_ASAP7_75t_R FILLER_53_171 ();
 DECAPx2_ASAP7_75t_R FILLER_53_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_185 ();
 DECAPx4_ASAP7_75t_R FILLER_53_192 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_202 ();
 DECAPx6_ASAP7_75t_R FILLER_53_231 ();
 DECAPx2_ASAP7_75t_R FILLER_53_253 ();
 FILLER_ASAP7_75t_R FILLER_53_259 ();
 FILLER_ASAP7_75t_R FILLER_53_269 ();
 FILLER_ASAP7_75t_R FILLER_53_280 ();
 DECAPx2_ASAP7_75t_R FILLER_53_285 ();
 DECAPx2_ASAP7_75t_R FILLER_53_297 ();
 DECAPx4_ASAP7_75t_R FILLER_53_309 ();
 DECAPx2_ASAP7_75t_R FILLER_53_325 ();
 FILLER_ASAP7_75t_R FILLER_53_337 ();
 FILLER_ASAP7_75t_R FILLER_53_345 ();
 FILLER_ASAP7_75t_R FILLER_53_355 ();
 DECAPx1_ASAP7_75t_R FILLER_53_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_387 ();
 FILLER_ASAP7_75t_R FILLER_53_414 ();
 DECAPx6_ASAP7_75t_R FILLER_53_442 ();
 FILLER_ASAP7_75t_R FILLER_53_456 ();
 DECAPx4_ASAP7_75t_R FILLER_53_461 ();
 FILLER_ASAP7_75t_R FILLER_53_477 ();
 DECAPx1_ASAP7_75t_R FILLER_53_485 ();
 DECAPx2_ASAP7_75t_R FILLER_53_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_498 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_502 ();
 DECAPx1_ASAP7_75t_R FILLER_53_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_517 ();
 FILLER_ASAP7_75t_R FILLER_53_524 ();
 FILLER_ASAP7_75t_R FILLER_53_533 ();
 FILLER_ASAP7_75t_R FILLER_53_542 ();
 DECAPx4_ASAP7_75t_R FILLER_53_550 ();
 DECAPx4_ASAP7_75t_R FILLER_53_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_578 ();
 DECAPx4_ASAP7_75t_R FILLER_53_589 ();
 FILLER_ASAP7_75t_R FILLER_53_613 ();
 DECAPx6_ASAP7_75t_R FILLER_53_625 ();
 DECAPx2_ASAP7_75t_R FILLER_53_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_645 ();
 DECAPx10_ASAP7_75t_R FILLER_53_652 ();
 FILLER_ASAP7_75t_R FILLER_53_674 ();
 DECAPx1_ASAP7_75t_R FILLER_53_686 ();
 DECAPx10_ASAP7_75t_R FILLER_53_696 ();
 DECAPx2_ASAP7_75t_R FILLER_53_738 ();
 DECAPx2_ASAP7_75t_R FILLER_53_751 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_757 ();
 DECAPx2_ASAP7_75t_R FILLER_53_786 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_792 ();
 DECAPx10_ASAP7_75t_R FILLER_53_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_823 ();
 DECAPx2_ASAP7_75t_R FILLER_53_830 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_836 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_842 ();
 DECAPx6_ASAP7_75t_R FILLER_53_853 ();
 DECAPx2_ASAP7_75t_R FILLER_53_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_873 ();
 FILLER_ASAP7_75t_R FILLER_53_882 ();
 FILLER_ASAP7_75t_R FILLER_53_892 ();
 DECAPx1_ASAP7_75t_R FILLER_53_902 ();
 DECAPx4_ASAP7_75t_R FILLER_53_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_922 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_927 ();
 DECAPx2_ASAP7_75t_R FILLER_53_933 ();
 DECAPx2_ASAP7_75t_R FILLER_53_945 ();
 FILLER_ASAP7_75t_R FILLER_53_961 ();
 FILLER_ASAP7_75t_R FILLER_53_971 ();
 DECAPx10_ASAP7_75t_R FILLER_53_981 ();
 DECAPx1_ASAP7_75t_R FILLER_53_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1010 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_53_1022 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1041 ();
 FILLER_ASAP7_75t_R FILLER_53_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1061 ();
 FILLER_ASAP7_75t_R FILLER_53_1067 ();
 DECAPx4_ASAP7_75t_R FILLER_53_1072 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_53_1095 ();
 DECAPx4_ASAP7_75t_R FILLER_53_1106 ();
 DECAPx6_ASAP7_75t_R FILLER_53_1126 ();
 FILLER_ASAP7_75t_R FILLER_53_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1170 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_1176 ();
 FILLER_ASAP7_75t_R FILLER_53_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1213 ();
 DECAPx4_ASAP7_75t_R FILLER_53_1235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1261 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1283 ();
 FILLER_ASAP7_75t_R FILLER_53_1289 ();
 FILLER_ASAP7_75t_R FILLER_53_1297 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1307 ();
 FILLER_ASAP7_75t_R FILLER_53_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_53_1321 ();
 DECAPx2_ASAP7_75t_R FILLER_53_1343 ();
 FILLER_ASAP7_75t_R FILLER_53_1349 ();
 FILLER_ASAP7_75t_R FILLER_53_1358 ();
 DECAPx4_ASAP7_75t_R FILLER_53_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_1376 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_2 ();
 DECAPx4_ASAP7_75t_R FILLER_54_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_41 ();
 DECAPx6_ASAP7_75t_R FILLER_54_50 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_64 ();
 FILLER_ASAP7_75t_R FILLER_54_73 ();
 DECAPx10_ASAP7_75t_R FILLER_54_81 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_103 ();
 DECAPx1_ASAP7_75t_R FILLER_54_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_136 ();
 DECAPx4_ASAP7_75t_R FILLER_54_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_154 ();
 DECAPx6_ASAP7_75t_R FILLER_54_161 ();
 DECAPx2_ASAP7_75t_R FILLER_54_175 ();
 DECAPx1_ASAP7_75t_R FILLER_54_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_211 ();
 FILLER_ASAP7_75t_R FILLER_54_219 ();
 FILLER_ASAP7_75t_R FILLER_54_228 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_233 ();
 FILLER_ASAP7_75t_R FILLER_54_242 ();
 DECAPx1_ASAP7_75t_R FILLER_54_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_256 ();
 FILLER_ASAP7_75t_R FILLER_54_263 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_291 ();
 FILLER_ASAP7_75t_R FILLER_54_297 ();
 FILLER_ASAP7_75t_R FILLER_54_305 ();
 DECAPx10_ASAP7_75t_R FILLER_54_315 ();
 DECAPx2_ASAP7_75t_R FILLER_54_337 ();
 FILLER_ASAP7_75t_R FILLER_54_346 ();
 DECAPx2_ASAP7_75t_R FILLER_54_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_360 ();
 DECAPx1_ASAP7_75t_R FILLER_54_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_371 ();
 FILLER_ASAP7_75t_R FILLER_54_378 ();
 FILLER_ASAP7_75t_R FILLER_54_386 ();
 DECAPx6_ASAP7_75t_R FILLER_54_391 ();
 DECAPx4_ASAP7_75t_R FILLER_54_408 ();
 DECAPx2_ASAP7_75t_R FILLER_54_424 ();
 FILLER_ASAP7_75t_R FILLER_54_433 ();
 FILLER_ASAP7_75t_R FILLER_54_441 ();
 DECAPx1_ASAP7_75t_R FILLER_54_450 ();
 FILLER_ASAP7_75t_R FILLER_54_460 ();
 DECAPx2_ASAP7_75t_R FILLER_54_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_470 ();
 DECAPx10_ASAP7_75t_R FILLER_54_479 ();
 DECAPx1_ASAP7_75t_R FILLER_54_501 ();
 DECAPx1_ASAP7_75t_R FILLER_54_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_517 ();
 FILLER_ASAP7_75t_R FILLER_54_540 ();
 DECAPx4_ASAP7_75t_R FILLER_54_548 ();
 FILLER_ASAP7_75t_R FILLER_54_566 ();
 DECAPx2_ASAP7_75t_R FILLER_54_574 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_580 ();
 DECAPx4_ASAP7_75t_R FILLER_54_589 ();
 FILLER_ASAP7_75t_R FILLER_54_599 ();
 DECAPx4_ASAP7_75t_R FILLER_54_607 ();
 FILLER_ASAP7_75t_R FILLER_54_617 ();
 FILLER_ASAP7_75t_R FILLER_54_628 ();
 DECAPx2_ASAP7_75t_R FILLER_54_636 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_642 ();
 DECAPx2_ASAP7_75t_R FILLER_54_651 ();
 DECAPx2_ASAP7_75t_R FILLER_54_663 ();
 FILLER_ASAP7_75t_R FILLER_54_669 ();
 DECAPx10_ASAP7_75t_R FILLER_54_677 ();
 DECAPx1_ASAP7_75t_R FILLER_54_699 ();
 DECAPx6_ASAP7_75t_R FILLER_54_709 ();
 DECAPx4_ASAP7_75t_R FILLER_54_729 ();
 FILLER_ASAP7_75t_R FILLER_54_739 ();
 DECAPx10_ASAP7_75t_R FILLER_54_761 ();
 DECAPx10_ASAP7_75t_R FILLER_54_783 ();
 FILLER_ASAP7_75t_R FILLER_54_811 ();
 DECAPx10_ASAP7_75t_R FILLER_54_819 ();
 DECAPx1_ASAP7_75t_R FILLER_54_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_845 ();
 DECAPx4_ASAP7_75t_R FILLER_54_852 ();
 DECAPx1_ASAP7_75t_R FILLER_54_868 ();
 DECAPx10_ASAP7_75t_R FILLER_54_878 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_900 ();
 FILLER_ASAP7_75t_R FILLER_54_911 ();
 DECAPx6_ASAP7_75t_R FILLER_54_921 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_935 ();
 DECAPx6_ASAP7_75t_R FILLER_54_944 ();
 DECAPx2_ASAP7_75t_R FILLER_54_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_964 ();
 DECAPx6_ASAP7_75t_R FILLER_54_971 ();
 DECAPx2_ASAP7_75t_R FILLER_54_985 ();
 DECAPx6_ASAP7_75t_R FILLER_54_999 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1028 ();
 FILLER_ASAP7_75t_R FILLER_54_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_54_1046 ();
 FILLER_ASAP7_75t_R FILLER_54_1052 ();
 FILLER_ASAP7_75t_R FILLER_54_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_54_1092 ();
 DECAPx6_ASAP7_75t_R FILLER_54_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1138 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_1149 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1155 ();
 DECAPx2_ASAP7_75t_R FILLER_54_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1185 ();
 FILLER_ASAP7_75t_R FILLER_54_1192 ();
 FILLER_ASAP7_75t_R FILLER_54_1200 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1209 ();
 DECAPx4_ASAP7_75t_R FILLER_54_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1227 ();
 DECAPx4_ASAP7_75t_R FILLER_54_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_54_1254 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_54_1287 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_1297 ();
 DECAPx1_ASAP7_75t_R FILLER_54_1310 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_1314 ();
 DECAPx2_ASAP7_75t_R FILLER_54_1341 ();
 FILLER_ASAP7_75t_R FILLER_54_1347 ();
 FILLER_ASAP7_75t_R FILLER_54_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_55_2 ();
 FILLER_ASAP7_75t_R FILLER_55_8 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_16 ();
 DECAPx2_ASAP7_75t_R FILLER_55_22 ();
 FILLER_ASAP7_75t_R FILLER_55_34 ();
 DECAPx1_ASAP7_75t_R FILLER_55_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_48 ();
 FILLER_ASAP7_75t_R FILLER_55_55 ();
 DECAPx4_ASAP7_75t_R FILLER_55_63 ();
 DECAPx2_ASAP7_75t_R FILLER_55_81 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_87 ();
 DECAPx4_ASAP7_75t_R FILLER_55_98 ();
 FILLER_ASAP7_75t_R FILLER_55_108 ();
 DECAPx1_ASAP7_75t_R FILLER_55_116 ();
 DECAPx2_ASAP7_75t_R FILLER_55_123 ();
 FILLER_ASAP7_75t_R FILLER_55_129 ();
 FILLER_ASAP7_75t_R FILLER_55_137 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_147 ();
 DECAPx4_ASAP7_75t_R FILLER_55_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_166 ();
 FILLER_ASAP7_75t_R FILLER_55_175 ();
 FILLER_ASAP7_75t_R FILLER_55_183 ();
 DECAPx1_ASAP7_75t_R FILLER_55_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_195 ();
 DECAPx1_ASAP7_75t_R FILLER_55_199 ();
 FILLER_ASAP7_75t_R FILLER_55_210 ();
 FILLER_ASAP7_75t_R FILLER_55_219 ();
 FILLER_ASAP7_75t_R FILLER_55_228 ();
 DECAPx4_ASAP7_75t_R FILLER_55_236 ();
 FILLER_ASAP7_75t_R FILLER_55_246 ();
 FILLER_ASAP7_75t_R FILLER_55_254 ();
 DECAPx1_ASAP7_75t_R FILLER_55_262 ();
 DECAPx2_ASAP7_75t_R FILLER_55_272 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_278 ();
 FILLER_ASAP7_75t_R FILLER_55_307 ();
 DECAPx2_ASAP7_75t_R FILLER_55_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_323 ();
 DECAPx2_ASAP7_75t_R FILLER_55_330 ();
 FILLER_ASAP7_75t_R FILLER_55_336 ();
 DECAPx1_ASAP7_75t_R FILLER_55_344 ();
 FILLER_ASAP7_75t_R FILLER_55_370 ();
 DECAPx10_ASAP7_75t_R FILLER_55_375 ();
 DECAPx10_ASAP7_75t_R FILLER_55_397 ();
 DECAPx1_ASAP7_75t_R FILLER_55_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_423 ();
 DECAPx2_ASAP7_75t_R FILLER_55_430 ();
 DECAPx1_ASAP7_75t_R FILLER_55_444 ();
 FILLER_ASAP7_75t_R FILLER_55_454 ();
 DECAPx1_ASAP7_75t_R FILLER_55_464 ();
 DECAPx2_ASAP7_75t_R FILLER_55_494 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_500 ();
 DECAPx2_ASAP7_75t_R FILLER_55_509 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_515 ();
 FILLER_ASAP7_75t_R FILLER_55_540 ();
 FILLER_ASAP7_75t_R FILLER_55_549 ();
 DECAPx2_ASAP7_75t_R FILLER_55_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_560 ();
 DECAPx4_ASAP7_75t_R FILLER_55_569 ();
 FILLER_ASAP7_75t_R FILLER_55_585 ();
 DECAPx10_ASAP7_75t_R FILLER_55_595 ();
 DECAPx2_ASAP7_75t_R FILLER_55_617 ();
 FILLER_ASAP7_75t_R FILLER_55_623 ();
 DECAPx1_ASAP7_75t_R FILLER_55_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_638 ();
 FILLER_ASAP7_75t_R FILLER_55_645 ();
 DECAPx2_ASAP7_75t_R FILLER_55_655 ();
 FILLER_ASAP7_75t_R FILLER_55_670 ();
 DECAPx2_ASAP7_75t_R FILLER_55_680 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_686 ();
 FILLER_ASAP7_75t_R FILLER_55_709 ();
 DECAPx10_ASAP7_75t_R FILLER_55_718 ();
 DECAPx2_ASAP7_75t_R FILLER_55_740 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_746 ();
 DECAPx6_ASAP7_75t_R FILLER_55_755 ();
 DECAPx1_ASAP7_75t_R FILLER_55_769 ();
 DECAPx2_ASAP7_75t_R FILLER_55_781 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_787 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_796 ();
 FILLER_ASAP7_75t_R FILLER_55_805 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_813 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_822 ();
 FILLER_ASAP7_75t_R FILLER_55_835 ();
 DECAPx10_ASAP7_75t_R FILLER_55_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_870 ();
 DECAPx10_ASAP7_75t_R FILLER_55_877 ();
 DECAPx1_ASAP7_75t_R FILLER_55_899 ();
 DECAPx6_ASAP7_75t_R FILLER_55_909 ();
 FILLER_ASAP7_75t_R FILLER_55_923 ();
 DECAPx2_ASAP7_75t_R FILLER_55_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_933 ();
 DECAPx4_ASAP7_75t_R FILLER_55_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_953 ();
 DECAPx6_ASAP7_75t_R FILLER_55_965 ();
 DECAPx2_ASAP7_75t_R FILLER_55_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_985 ();
 FILLER_ASAP7_75t_R FILLER_55_994 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1006 ();
 FILLER_ASAP7_75t_R FILLER_55_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1049 ();
 FILLER_ASAP7_75t_R FILLER_55_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1067 ();
 DECAPx4_ASAP7_75t_R FILLER_55_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1099 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1106 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_1115 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1153 ();
 DECAPx1_ASAP7_75t_R FILLER_55_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_55_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1204 ();
 FILLER_ASAP7_75t_R FILLER_55_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1238 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_1251 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1257 ();
 FILLER_ASAP7_75t_R FILLER_55_1269 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1297 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_1303 ();
 FILLER_ASAP7_75t_R FILLER_55_1312 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_1321 ();
 FILLER_ASAP7_75t_R FILLER_55_1327 ();
 DECAPx4_ASAP7_75t_R FILLER_55_1341 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1351 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_1365 ();
 DECAPx2_ASAP7_75t_R FILLER_55_1369 ();
 FILLER_ASAP7_75t_R FILLER_55_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_56_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_8 ();
 DECAPx6_ASAP7_75t_R FILLER_56_17 ();
 DECAPx6_ASAP7_75t_R FILLER_56_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_48 ();
 DECAPx1_ASAP7_75t_R FILLER_56_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_61 ();
 FILLER_ASAP7_75t_R FILLER_56_70 ();
 DECAPx1_ASAP7_75t_R FILLER_56_78 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_88 ();
 FILLER_ASAP7_75t_R FILLER_56_97 ();
 DECAPx4_ASAP7_75t_R FILLER_56_102 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_112 ();
 DECAPx2_ASAP7_75t_R FILLER_56_121 ();
 FILLER_ASAP7_75t_R FILLER_56_127 ();
 FILLER_ASAP7_75t_R FILLER_56_132 ();
 DECAPx6_ASAP7_75t_R FILLER_56_140 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_154 ();
 DECAPx1_ASAP7_75t_R FILLER_56_163 ();
 DECAPx2_ASAP7_75t_R FILLER_56_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_195 ();
 DECAPx2_ASAP7_75t_R FILLER_56_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_228 ();
 FILLER_ASAP7_75t_R FILLER_56_237 ();
 DECAPx10_ASAP7_75t_R FILLER_56_245 ();
 DECAPx4_ASAP7_75t_R FILLER_56_267 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_277 ();
 DECAPx2_ASAP7_75t_R FILLER_56_302 ();
 FILLER_ASAP7_75t_R FILLER_56_314 ();
 FILLER_ASAP7_75t_R FILLER_56_342 ();
 DECAPx4_ASAP7_75t_R FILLER_56_354 ();
 FILLER_ASAP7_75t_R FILLER_56_364 ();
 DECAPx2_ASAP7_75t_R FILLER_56_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_378 ();
 DECAPx1_ASAP7_75t_R FILLER_56_385 ();
 DECAPx1_ASAP7_75t_R FILLER_56_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_399 ();
 FILLER_ASAP7_75t_R FILLER_56_426 ();
 DECAPx2_ASAP7_75t_R FILLER_56_434 ();
 DECAPx2_ASAP7_75t_R FILLER_56_446 ();
 FILLER_ASAP7_75t_R FILLER_56_460 ();
 FILLER_ASAP7_75t_R FILLER_56_464 ();
 DECAPx2_ASAP7_75t_R FILLER_56_488 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_500 ();
 DECAPx2_ASAP7_75t_R FILLER_56_509 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_515 ();
 FILLER_ASAP7_75t_R FILLER_56_524 ();
 DECAPx4_ASAP7_75t_R FILLER_56_552 ();
 DECAPx2_ASAP7_75t_R FILLER_56_570 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_576 ();
 DECAPx6_ASAP7_75t_R FILLER_56_587 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_601 ();
 DECAPx4_ASAP7_75t_R FILLER_56_613 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_623 ();
 DECAPx1_ASAP7_75t_R FILLER_56_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_640 ();
 FILLER_ASAP7_75t_R FILLER_56_647 ();
 DECAPx4_ASAP7_75t_R FILLER_56_652 ();
 FILLER_ASAP7_75t_R FILLER_56_662 ();
 DECAPx4_ASAP7_75t_R FILLER_56_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_680 ();
 FILLER_ASAP7_75t_R FILLER_56_693 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_702 ();
 DECAPx1_ASAP7_75t_R FILLER_56_725 ();
 DECAPx1_ASAP7_75t_R FILLER_56_735 ();
 FILLER_ASAP7_75t_R FILLER_56_745 ();
 FILLER_ASAP7_75t_R FILLER_56_754 ();
 FILLER_ASAP7_75t_R FILLER_56_762 ();
 FILLER_ASAP7_75t_R FILLER_56_770 ();
 DECAPx2_ASAP7_75t_R FILLER_56_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_787 ();
 FILLER_ASAP7_75t_R FILLER_56_795 ();
 DECAPx2_ASAP7_75t_R FILLER_56_804 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_810 ();
 FILLER_ASAP7_75t_R FILLER_56_821 ();
 DECAPx1_ASAP7_75t_R FILLER_56_831 ();
 FILLER_ASAP7_75t_R FILLER_56_842 ();
 DECAPx4_ASAP7_75t_R FILLER_56_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_864 ();
 FILLER_ASAP7_75t_R FILLER_56_873 ();
 DECAPx1_ASAP7_75t_R FILLER_56_882 ();
 FILLER_ASAP7_75t_R FILLER_56_894 ();
 DECAPx2_ASAP7_75t_R FILLER_56_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_908 ();
 DECAPx2_ASAP7_75t_R FILLER_56_915 ();
 FILLER_ASAP7_75t_R FILLER_56_927 ();
 FILLER_ASAP7_75t_R FILLER_56_937 ();
 FILLER_ASAP7_75t_R FILLER_56_947 ();
 FILLER_ASAP7_75t_R FILLER_56_952 ();
 DECAPx2_ASAP7_75t_R FILLER_56_960 ();
 FILLER_ASAP7_75t_R FILLER_56_966 ();
 DECAPx1_ASAP7_75t_R FILLER_56_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_978 ();
 DECAPx1_ASAP7_75t_R FILLER_56_982 ();
 FILLER_ASAP7_75t_R FILLER_56_995 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1009 ();
 FILLER_ASAP7_75t_R FILLER_56_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_56_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1036 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1091 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1119 ();
 FILLER_ASAP7_75t_R FILLER_56_1130 ();
 FILLER_ASAP7_75t_R FILLER_56_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1147 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_1153 ();
 DECAPx4_ASAP7_75t_R FILLER_56_1159 ();
 FILLER_ASAP7_75t_R FILLER_56_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_56_1177 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_1187 ();
 FILLER_ASAP7_75t_R FILLER_56_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1211 ();
 DECAPx6_ASAP7_75t_R FILLER_56_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1238 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_1266 ();
 FILLER_ASAP7_75t_R FILLER_56_1277 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_1282 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_56_1303 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1325 ();
 FILLER_ASAP7_75t_R FILLER_56_1331 ();
 DECAPx2_ASAP7_75t_R FILLER_56_1341 ();
 FILLER_ASAP7_75t_R FILLER_56_1347 ();
 FILLER_ASAP7_75t_R FILLER_56_1375 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_2 ();
 FILLER_ASAP7_75t_R FILLER_57_31 ();
 DECAPx6_ASAP7_75t_R FILLER_57_36 ();
 DECAPx4_ASAP7_75t_R FILLER_57_56 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_66 ();
 DECAPx10_ASAP7_75t_R FILLER_57_72 ();
 DECAPx4_ASAP7_75t_R FILLER_57_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_104 ();
 DECAPx6_ASAP7_75t_R FILLER_57_131 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_145 ();
 DECAPx2_ASAP7_75t_R FILLER_57_156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_162 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_171 ();
 DECAPx6_ASAP7_75t_R FILLER_57_186 ();
 FILLER_ASAP7_75t_R FILLER_57_200 ();
 FILLER_ASAP7_75t_R FILLER_57_208 ();
 FILLER_ASAP7_75t_R FILLER_57_216 ();
 FILLER_ASAP7_75t_R FILLER_57_221 ();
 DECAPx1_ASAP7_75t_R FILLER_57_226 ();
 DECAPx2_ASAP7_75t_R FILLER_57_238 ();
 FILLER_ASAP7_75t_R FILLER_57_250 ();
 FILLER_ASAP7_75t_R FILLER_57_258 ();
 DECAPx6_ASAP7_75t_R FILLER_57_263 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_283 ();
 DECAPx10_ASAP7_75t_R FILLER_57_292 ();
 DECAPx2_ASAP7_75t_R FILLER_57_314 ();
 DECAPx1_ASAP7_75t_R FILLER_57_326 ();
 DECAPx1_ASAP7_75t_R FILLER_57_333 ();
 DECAPx6_ASAP7_75t_R FILLER_57_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_358 ();
 FILLER_ASAP7_75t_R FILLER_57_385 ();
 FILLER_ASAP7_75t_R FILLER_57_390 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_400 ();
 FILLER_ASAP7_75t_R FILLER_57_409 ();
 FILLER_ASAP7_75t_R FILLER_57_417 ();
 DECAPx10_ASAP7_75t_R FILLER_57_422 ();
 DECAPx4_ASAP7_75t_R FILLER_57_444 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_454 ();
 DECAPx6_ASAP7_75t_R FILLER_57_463 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_477 ();
 FILLER_ASAP7_75t_R FILLER_57_483 ();
 DECAPx2_ASAP7_75t_R FILLER_57_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_517 ();
 FILLER_ASAP7_75t_R FILLER_57_524 ();
 FILLER_ASAP7_75t_R FILLER_57_533 ();
 FILLER_ASAP7_75t_R FILLER_57_542 ();
 DECAPx2_ASAP7_75t_R FILLER_57_551 ();
 DECAPx2_ASAP7_75t_R FILLER_57_565 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_571 ();
 DECAPx2_ASAP7_75t_R FILLER_57_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_586 ();
 DECAPx2_ASAP7_75t_R FILLER_57_593 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_599 ();
 FILLER_ASAP7_75t_R FILLER_57_612 ();
 DECAPx1_ASAP7_75t_R FILLER_57_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_624 ();
 DECAPx10_ASAP7_75t_R FILLER_57_631 ();
 DECAPx4_ASAP7_75t_R FILLER_57_653 ();
 FILLER_ASAP7_75t_R FILLER_57_663 ();
 DECAPx2_ASAP7_75t_R FILLER_57_672 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_678 ();
 DECAPx10_ASAP7_75t_R FILLER_57_687 ();
 DECAPx4_ASAP7_75t_R FILLER_57_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_719 ();
 FILLER_ASAP7_75t_R FILLER_57_740 ();
 FILLER_ASAP7_75t_R FILLER_57_764 ();
 DECAPx10_ASAP7_75t_R FILLER_57_774 ();
 DECAPx2_ASAP7_75t_R FILLER_57_796 ();
 FILLER_ASAP7_75t_R FILLER_57_802 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_810 ();
 DECAPx10_ASAP7_75t_R FILLER_57_819 ();
 FILLER_ASAP7_75t_R FILLER_57_850 ();
 FILLER_ASAP7_75t_R FILLER_57_861 ();
 DECAPx4_ASAP7_75t_R FILLER_57_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_881 ();
 FILLER_ASAP7_75t_R FILLER_57_888 ();
 DECAPx2_ASAP7_75t_R FILLER_57_896 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_902 ();
 FILLER_ASAP7_75t_R FILLER_57_914 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_922 ();
 FILLER_ASAP7_75t_R FILLER_57_927 ();
 FILLER_ASAP7_75t_R FILLER_57_939 ();
 DECAPx6_ASAP7_75t_R FILLER_57_947 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_961 ();
 FILLER_ASAP7_75t_R FILLER_57_973 ();
 DECAPx2_ASAP7_75t_R FILLER_57_981 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_987 ();
 FILLER_ASAP7_75t_R FILLER_57_996 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1008 ();
 DECAPx6_ASAP7_75t_R FILLER_57_1012 ();
 FILLER_ASAP7_75t_R FILLER_57_1034 ();
 FILLER_ASAP7_75t_R FILLER_57_1042 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1079 ();
 DECAPx6_ASAP7_75t_R FILLER_57_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1154 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1167 ();
 FILLER_ASAP7_75t_R FILLER_57_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1178 ();
 FILLER_ASAP7_75t_R FILLER_57_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_57_1234 ();
 DECAPx4_ASAP7_75t_R FILLER_57_1256 ();
 DECAPx6_ASAP7_75t_R FILLER_57_1272 ();
 DECAPx1_ASAP7_75t_R FILLER_57_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_1290 ();
 DECAPx6_ASAP7_75t_R FILLER_57_1297 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_1311 ();
 FILLER_ASAP7_75t_R FILLER_57_1321 ();
 FILLER_ASAP7_75t_R FILLER_57_1329 ();
 DECAPx6_ASAP7_75t_R FILLER_57_1334 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1348 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1360 ();
 DECAPx2_ASAP7_75t_R FILLER_57_1369 ();
 FILLER_ASAP7_75t_R FILLER_57_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_58_2 ();
 DECAPx1_ASAP7_75t_R FILLER_58_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_18 ();
 DECAPx10_ASAP7_75t_R FILLER_58_22 ();
 DECAPx1_ASAP7_75t_R FILLER_58_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_74 ();
 DECAPx2_ASAP7_75t_R FILLER_58_81 ();
 DECAPx2_ASAP7_75t_R FILLER_58_90 ();
 FILLER_ASAP7_75t_R FILLER_58_96 ();
 FILLER_ASAP7_75t_R FILLER_58_110 ();
 FILLER_ASAP7_75t_R FILLER_58_118 ();
 DECAPx6_ASAP7_75t_R FILLER_58_123 ();
 DECAPx2_ASAP7_75t_R FILLER_58_137 ();
 FILLER_ASAP7_75t_R FILLER_58_149 ();
 DECAPx10_ASAP7_75t_R FILLER_58_159 ();
 DECAPx2_ASAP7_75t_R FILLER_58_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_187 ();
 FILLER_ASAP7_75t_R FILLER_58_194 ();
 DECAPx10_ASAP7_75t_R FILLER_58_199 ();
 DECAPx6_ASAP7_75t_R FILLER_58_221 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_235 ();
 FILLER_ASAP7_75t_R FILLER_58_264 ();
 DECAPx2_ASAP7_75t_R FILLER_58_292 ();
 FILLER_ASAP7_75t_R FILLER_58_298 ();
 FILLER_ASAP7_75t_R FILLER_58_306 ();
 DECAPx10_ASAP7_75t_R FILLER_58_311 ();
 DECAPx6_ASAP7_75t_R FILLER_58_333 ();
 DECAPx1_ASAP7_75t_R FILLER_58_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_351 ();
 FILLER_ASAP7_75t_R FILLER_58_360 ();
 DECAPx1_ASAP7_75t_R FILLER_58_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_372 ();
 FILLER_ASAP7_75t_R FILLER_58_376 ();
 DECAPx4_ASAP7_75t_R FILLER_58_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_396 ();
 DECAPx10_ASAP7_75t_R FILLER_58_403 ();
 DECAPx1_ASAP7_75t_R FILLER_58_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_429 ();
 DECAPx4_ASAP7_75t_R FILLER_58_436 ();
 FILLER_ASAP7_75t_R FILLER_58_446 ();
 DECAPx2_ASAP7_75t_R FILLER_58_456 ();
 DECAPx10_ASAP7_75t_R FILLER_58_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_486 ();
 DECAPx2_ASAP7_75t_R FILLER_58_493 ();
 DECAPx6_ASAP7_75t_R FILLER_58_502 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_516 ();
 DECAPx2_ASAP7_75t_R FILLER_58_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_531 ();
 FILLER_ASAP7_75t_R FILLER_58_539 ();
 FILLER_ASAP7_75t_R FILLER_58_547 ();
 FILLER_ASAP7_75t_R FILLER_58_555 ();
 DECAPx2_ASAP7_75t_R FILLER_58_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_570 ();
 DECAPx2_ASAP7_75t_R FILLER_58_577 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_583 ();
 DECAPx1_ASAP7_75t_R FILLER_58_593 ();
 DECAPx2_ASAP7_75t_R FILLER_58_603 ();
 DECAPx2_ASAP7_75t_R FILLER_58_615 ();
 FILLER_ASAP7_75t_R FILLER_58_627 ();
 DECAPx1_ASAP7_75t_R FILLER_58_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_639 ();
 FILLER_ASAP7_75t_R FILLER_58_650 ();
 DECAPx2_ASAP7_75t_R FILLER_58_658 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_664 ();
 DECAPx2_ASAP7_75t_R FILLER_58_677 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_683 ();
 DECAPx1_ASAP7_75t_R FILLER_58_690 ();
 FILLER_ASAP7_75t_R FILLER_58_701 ();
 DECAPx4_ASAP7_75t_R FILLER_58_709 ();
 DECAPx1_ASAP7_75t_R FILLER_58_726 ();
 DECAPx6_ASAP7_75t_R FILLER_58_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_747 ();
 DECAPx1_ASAP7_75t_R FILLER_58_754 ();
 DECAPx4_ASAP7_75t_R FILLER_58_766 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_776 ();
 FILLER_ASAP7_75t_R FILLER_58_786 ();
 DECAPx10_ASAP7_75t_R FILLER_58_798 ();
 DECAPx2_ASAP7_75t_R FILLER_58_820 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_826 ();
 FILLER_ASAP7_75t_R FILLER_58_836 ();
 DECAPx6_ASAP7_75t_R FILLER_58_844 ();
 FILLER_ASAP7_75t_R FILLER_58_858 ();
 FILLER_ASAP7_75t_R FILLER_58_866 ();
 DECAPx10_ASAP7_75t_R FILLER_58_874 ();
 DECAPx4_ASAP7_75t_R FILLER_58_896 ();
 DECAPx10_ASAP7_75t_R FILLER_58_909 ();
 DECAPx6_ASAP7_75t_R FILLER_58_931 ();
 DECAPx1_ASAP7_75t_R FILLER_58_945 ();
 FILLER_ASAP7_75t_R FILLER_58_955 ();
 FILLER_ASAP7_75t_R FILLER_58_963 ();
 DECAPx10_ASAP7_75t_R FILLER_58_968 ();
 DECAPx6_ASAP7_75t_R FILLER_58_990 ();
 FILLER_ASAP7_75t_R FILLER_58_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_58_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1056 ();
 FILLER_ASAP7_75t_R FILLER_58_1067 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1078 ();
 FILLER_ASAP7_75t_R FILLER_58_1084 ();
 FILLER_ASAP7_75t_R FILLER_58_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_58_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_58_1167 ();
 FILLER_ASAP7_75t_R FILLER_58_1197 ();
 DECAPx1_ASAP7_75t_R FILLER_58_1211 ();
 FILLER_ASAP7_75t_R FILLER_58_1241 ();
 FILLER_ASAP7_75t_R FILLER_58_1252 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_1298 ();
 DECAPx2_ASAP7_75t_R FILLER_58_1309 ();
 DECAPx6_ASAP7_75t_R FILLER_58_1341 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_1355 ();
 DECAPx4_ASAP7_75t_R FILLER_58_1365 ();
 FILLER_ASAP7_75t_R FILLER_58_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_59_2 ();
 FILLER_ASAP7_75t_R FILLER_59_30 ();
 DECAPx2_ASAP7_75t_R FILLER_59_38 ();
 FILLER_ASAP7_75t_R FILLER_59_44 ();
 DECAPx2_ASAP7_75t_R FILLER_59_52 ();
 DECAPx4_ASAP7_75t_R FILLER_59_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_71 ();
 FILLER_ASAP7_75t_R FILLER_59_98 ();
 DECAPx4_ASAP7_75t_R FILLER_59_112 ();
 FILLER_ASAP7_75t_R FILLER_59_128 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_136 ();
 FILLER_ASAP7_75t_R FILLER_59_142 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_147 ();
 DECAPx2_ASAP7_75t_R FILLER_59_156 ();
 DECAPx2_ASAP7_75t_R FILLER_59_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_174 ();
 DECAPx2_ASAP7_75t_R FILLER_59_201 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_207 ();
 DECAPx10_ASAP7_75t_R FILLER_59_216 ();
 DECAPx4_ASAP7_75t_R FILLER_59_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_248 ();
 FILLER_ASAP7_75t_R FILLER_59_255 ();
 DECAPx2_ASAP7_75t_R FILLER_59_263 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_269 ();
 FILLER_ASAP7_75t_R FILLER_59_278 ();
 DECAPx1_ASAP7_75t_R FILLER_59_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_287 ();
 DECAPx2_ASAP7_75t_R FILLER_59_314 ();
 FILLER_ASAP7_75t_R FILLER_59_320 ();
 DECAPx2_ASAP7_75t_R FILLER_59_328 ();
 DECAPx6_ASAP7_75t_R FILLER_59_340 ();
 DECAPx6_ASAP7_75t_R FILLER_59_361 ();
 DECAPx1_ASAP7_75t_R FILLER_59_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_379 ();
 DECAPx10_ASAP7_75t_R FILLER_59_386 ();
 DECAPx2_ASAP7_75t_R FILLER_59_408 ();
 FILLER_ASAP7_75t_R FILLER_59_420 ();
 DECAPx2_ASAP7_75t_R FILLER_59_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_431 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_443 ();
 FILLER_ASAP7_75t_R FILLER_59_454 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_464 ();
 DECAPx4_ASAP7_75t_R FILLER_59_493 ();
 FILLER_ASAP7_75t_R FILLER_59_503 ();
 FILLER_ASAP7_75t_R FILLER_59_511 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_539 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_545 ();
 FILLER_ASAP7_75t_R FILLER_59_554 ();
 FILLER_ASAP7_75t_R FILLER_59_562 ();
 DECAPx6_ASAP7_75t_R FILLER_59_570 ();
 DECAPx2_ASAP7_75t_R FILLER_59_584 ();
 DECAPx4_ASAP7_75t_R FILLER_59_599 ();
 DECAPx2_ASAP7_75t_R FILLER_59_617 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_623 ();
 DECAPx2_ASAP7_75t_R FILLER_59_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_641 ();
 FILLER_ASAP7_75t_R FILLER_59_648 ();
 DECAPx2_ASAP7_75t_R FILLER_59_662 ();
 FILLER_ASAP7_75t_R FILLER_59_668 ();
 DECAPx6_ASAP7_75t_R FILLER_59_678 ();
 DECAPx1_ASAP7_75t_R FILLER_59_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_716 ();
 DECAPx6_ASAP7_75t_R FILLER_59_723 ();
 DECAPx2_ASAP7_75t_R FILLER_59_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_743 ();
 DECAPx2_ASAP7_75t_R FILLER_59_750 ();
 FILLER_ASAP7_75t_R FILLER_59_764 ();
 DECAPx10_ASAP7_75t_R FILLER_59_774 ();
 DECAPx4_ASAP7_75t_R FILLER_59_799 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_815 ();
 DECAPx2_ASAP7_75t_R FILLER_59_821 ();
 FILLER_ASAP7_75t_R FILLER_59_827 ();
 DECAPx4_ASAP7_75t_R FILLER_59_849 ();
 DECAPx10_ASAP7_75t_R FILLER_59_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_887 ();
 DECAPx2_ASAP7_75t_R FILLER_59_896 ();
 FILLER_ASAP7_75t_R FILLER_59_902 ();
 DECAPx6_ASAP7_75t_R FILLER_59_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_924 ();
 DECAPx10_ASAP7_75t_R FILLER_59_927 ();
 DECAPx6_ASAP7_75t_R FILLER_59_949 ();
 FILLER_ASAP7_75t_R FILLER_59_963 ();
 FILLER_ASAP7_75t_R FILLER_59_971 ();
 DECAPx2_ASAP7_75t_R FILLER_59_981 ();
 FILLER_ASAP7_75t_R FILLER_59_987 ();
 DECAPx2_ASAP7_75t_R FILLER_59_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1012 ();
 DECAPx6_ASAP7_75t_R FILLER_59_1021 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_1035 ();
 FILLER_ASAP7_75t_R FILLER_59_1045 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1053 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_1059 ();
 FILLER_ASAP7_75t_R FILLER_59_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1096 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_1102 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_59_1130 ();
 FILLER_ASAP7_75t_R FILLER_59_1144 ();
 FILLER_ASAP7_75t_R FILLER_59_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1177 ();
 FILLER_ASAP7_75t_R FILLER_59_1183 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1188 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_1198 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1204 ();
 FILLER_ASAP7_75t_R FILLER_59_1220 ();
 FILLER_ASAP7_75t_R FILLER_59_1230 ();
 DECAPx1_ASAP7_75t_R FILLER_59_1235 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1246 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_1252 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1281 ();
 FILLER_ASAP7_75t_R FILLER_59_1313 ();
 DECAPx4_ASAP7_75t_R FILLER_59_1321 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1331 ();
 DECAPx2_ASAP7_75t_R FILLER_59_1342 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_1348 ();
 FILLER_ASAP7_75t_R FILLER_59_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_60_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_8 ();
 DECAPx1_ASAP7_75t_R FILLER_60_15 ();
 DECAPx10_ASAP7_75t_R FILLER_60_45 ();
 DECAPx2_ASAP7_75t_R FILLER_60_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_73 ();
 DECAPx2_ASAP7_75t_R FILLER_60_80 ();
 FILLER_ASAP7_75t_R FILLER_60_86 ();
 DECAPx1_ASAP7_75t_R FILLER_60_94 ();
 DECAPx1_ASAP7_75t_R FILLER_60_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_105 ();
 FILLER_ASAP7_75t_R FILLER_60_112 ();
 DECAPx1_ASAP7_75t_R FILLER_60_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_124 ();
 DECAPx2_ASAP7_75t_R FILLER_60_151 ();
 FILLER_ASAP7_75t_R FILLER_60_183 ();
 DECAPx2_ASAP7_75t_R FILLER_60_191 ();
 FILLER_ASAP7_75t_R FILLER_60_223 ();
 FILLER_ASAP7_75t_R FILLER_60_228 ();
 FILLER_ASAP7_75t_R FILLER_60_238 ();
 DECAPx10_ASAP7_75t_R FILLER_60_246 ();
 DECAPx4_ASAP7_75t_R FILLER_60_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_278 ();
 DECAPx4_ASAP7_75t_R FILLER_60_285 ();
 FILLER_ASAP7_75t_R FILLER_60_301 ();
 DECAPx2_ASAP7_75t_R FILLER_60_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_312 ();
 FILLER_ASAP7_75t_R FILLER_60_339 ();
 FILLER_ASAP7_75t_R FILLER_60_349 ();
 DECAPx10_ASAP7_75t_R FILLER_60_357 ();
 DECAPx2_ASAP7_75t_R FILLER_60_379 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_385 ();
 DECAPx4_ASAP7_75t_R FILLER_60_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_406 ();
 DECAPx1_ASAP7_75t_R FILLER_60_433 ();
 DECAPx2_ASAP7_75t_R FILLER_60_445 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_451 ();
 FILLER_ASAP7_75t_R FILLER_60_460 ();
 DECAPx1_ASAP7_75t_R FILLER_60_464 ();
 FILLER_ASAP7_75t_R FILLER_60_471 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_479 ();
 DECAPx2_ASAP7_75t_R FILLER_60_485 ();
 DECAPx2_ASAP7_75t_R FILLER_60_517 ();
 FILLER_ASAP7_75t_R FILLER_60_523 ();
 FILLER_ASAP7_75t_R FILLER_60_531 ();
 FILLER_ASAP7_75t_R FILLER_60_541 ();
 DECAPx2_ASAP7_75t_R FILLER_60_549 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_555 ();
 DECAPx6_ASAP7_75t_R FILLER_60_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_578 ();
 FILLER_ASAP7_75t_R FILLER_60_585 ();
 DECAPx6_ASAP7_75t_R FILLER_60_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_607 ();
 DECAPx4_ASAP7_75t_R FILLER_60_618 ();
 DECAPx4_ASAP7_75t_R FILLER_60_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_648 ();
 DECAPx2_ASAP7_75t_R FILLER_60_656 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_662 ();
 FILLER_ASAP7_75t_R FILLER_60_671 ();
 DECAPx10_ASAP7_75t_R FILLER_60_679 ();
 DECAPx2_ASAP7_75t_R FILLER_60_701 ();
 FILLER_ASAP7_75t_R FILLER_60_707 ();
 FILLER_ASAP7_75t_R FILLER_60_729 ();
 DECAPx10_ASAP7_75t_R FILLER_60_738 ();
 FILLER_ASAP7_75t_R FILLER_60_760 ();
 DECAPx2_ASAP7_75t_R FILLER_60_770 ();
 FILLER_ASAP7_75t_R FILLER_60_782 ();
 FILLER_ASAP7_75t_R FILLER_60_791 ();
 DECAPx1_ASAP7_75t_R FILLER_60_800 ();
 DECAPx1_ASAP7_75t_R FILLER_60_807 ();
 DECAPx2_ASAP7_75t_R FILLER_60_814 ();
 FILLER_ASAP7_75t_R FILLER_60_820 ();
 DECAPx6_ASAP7_75t_R FILLER_60_832 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_846 ();
 DECAPx2_ASAP7_75t_R FILLER_60_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_858 ();
 DECAPx1_ASAP7_75t_R FILLER_60_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_872 ();
 FILLER_ASAP7_75t_R FILLER_60_876 ();
 FILLER_ASAP7_75t_R FILLER_60_887 ();
 FILLER_ASAP7_75t_R FILLER_60_897 ();
 FILLER_ASAP7_75t_R FILLER_60_905 ();
 DECAPx6_ASAP7_75t_R FILLER_60_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_928 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_936 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_947 ();
 DECAPx4_ASAP7_75t_R FILLER_60_976 ();
 FILLER_ASAP7_75t_R FILLER_60_986 ();
 FILLER_ASAP7_75t_R FILLER_60_996 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1028 ();
 FILLER_ASAP7_75t_R FILLER_60_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1062 ();
 DECAPx4_ASAP7_75t_R FILLER_60_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1080 ();
 DECAPx6_ASAP7_75t_R FILLER_60_1102 ();
 FILLER_ASAP7_75t_R FILLER_60_1116 ();
 FILLER_ASAP7_75t_R FILLER_60_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1172 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1194 ();
 DECAPx6_ASAP7_75t_R FILLER_60_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1219 ();
 DECAPx4_ASAP7_75t_R FILLER_60_1228 ();
 FILLER_ASAP7_75t_R FILLER_60_1250 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1263 ();
 FILLER_ASAP7_75t_R FILLER_60_1274 ();
 FILLER_ASAP7_75t_R FILLER_60_1279 ();
 DECAPx2_ASAP7_75t_R FILLER_60_1284 ();
 FILLER_ASAP7_75t_R FILLER_60_1290 ();
 FILLER_ASAP7_75t_R FILLER_60_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_60_1305 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_1327 ();
 FILLER_ASAP7_75t_R FILLER_60_1336 ();
 FILLER_ASAP7_75t_R FILLER_60_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_60_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_1376 ();
 FILLER_ASAP7_75t_R FILLER_61_2 ();
 FILLER_ASAP7_75t_R FILLER_61_30 ();
 DECAPx1_ASAP7_75t_R FILLER_61_39 ();
 FILLER_ASAP7_75t_R FILLER_61_51 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_56 ();
 DECAPx4_ASAP7_75t_R FILLER_61_67 ();
 FILLER_ASAP7_75t_R FILLER_61_77 ();
 FILLER_ASAP7_75t_R FILLER_61_105 ();
 DECAPx10_ASAP7_75t_R FILLER_61_133 ();
 DECAPx4_ASAP7_75t_R FILLER_61_155 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_165 ();
 FILLER_ASAP7_75t_R FILLER_61_174 ();
 DECAPx10_ASAP7_75t_R FILLER_61_179 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_201 ();
 FILLER_ASAP7_75t_R FILLER_61_210 ();
 DECAPx2_ASAP7_75t_R FILLER_61_215 ();
 FILLER_ASAP7_75t_R FILLER_61_221 ();
 FILLER_ASAP7_75t_R FILLER_61_229 ();
 FILLER_ASAP7_75t_R FILLER_61_239 ();
 DECAPx2_ASAP7_75t_R FILLER_61_247 ();
 FILLER_ASAP7_75t_R FILLER_61_253 ();
 DECAPx4_ASAP7_75t_R FILLER_61_261 ();
 FILLER_ASAP7_75t_R FILLER_61_277 ();
 FILLER_ASAP7_75t_R FILLER_61_301 ();
 DECAPx2_ASAP7_75t_R FILLER_61_309 ();
 FILLER_ASAP7_75t_R FILLER_61_315 ();
 DECAPx1_ASAP7_75t_R FILLER_61_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_327 ();
 DECAPx2_ASAP7_75t_R FILLER_61_331 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_337 ();
 DECAPx6_ASAP7_75t_R FILLER_61_343 ();
 DECAPx1_ASAP7_75t_R FILLER_61_383 ();
 FILLER_ASAP7_75t_R FILLER_61_393 ();
 DECAPx1_ASAP7_75t_R FILLER_61_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_409 ();
 DECAPx4_ASAP7_75t_R FILLER_61_416 ();
 FILLER_ASAP7_75t_R FILLER_61_440 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_448 ();
 DECAPx6_ASAP7_75t_R FILLER_61_457 ();
 DECAPx6_ASAP7_75t_R FILLER_61_477 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_491 ();
 DECAPx2_ASAP7_75t_R FILLER_61_500 ();
 FILLER_ASAP7_75t_R FILLER_61_512 ();
 DECAPx4_ASAP7_75t_R FILLER_61_517 ();
 FILLER_ASAP7_75t_R FILLER_61_530 ();
 DECAPx6_ASAP7_75t_R FILLER_61_540 ();
 DECAPx1_ASAP7_75t_R FILLER_61_554 ();
 DECAPx1_ASAP7_75t_R FILLER_61_564 ();
 FILLER_ASAP7_75t_R FILLER_61_574 ();
 FILLER_ASAP7_75t_R FILLER_61_582 ();
 DECAPx2_ASAP7_75t_R FILLER_61_590 ();
 FILLER_ASAP7_75t_R FILLER_61_596 ();
 FILLER_ASAP7_75t_R FILLER_61_604 ();
 DECAPx10_ASAP7_75t_R FILLER_61_618 ();
 DECAPx2_ASAP7_75t_R FILLER_61_640 ();
 FILLER_ASAP7_75t_R FILLER_61_646 ();
 FILLER_ASAP7_75t_R FILLER_61_654 ();
 DECAPx2_ASAP7_75t_R FILLER_61_662 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_668 ();
 DECAPx2_ASAP7_75t_R FILLER_61_677 ();
 FILLER_ASAP7_75t_R FILLER_61_690 ();
 DECAPx4_ASAP7_75t_R FILLER_61_698 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_708 ();
 DECAPx4_ASAP7_75t_R FILLER_61_718 ();
 FILLER_ASAP7_75t_R FILLER_61_728 ();
 DECAPx2_ASAP7_75t_R FILLER_61_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_756 ();
 DECAPx6_ASAP7_75t_R FILLER_61_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_777 ();
 FILLER_ASAP7_75t_R FILLER_61_784 ();
 DECAPx2_ASAP7_75t_R FILLER_61_792 ();
 FILLER_ASAP7_75t_R FILLER_61_798 ();
 DECAPx10_ASAP7_75t_R FILLER_61_803 ();
 FILLER_ASAP7_75t_R FILLER_61_825 ();
 DECAPx2_ASAP7_75t_R FILLER_61_835 ();
 FILLER_ASAP7_75t_R FILLER_61_841 ();
 DECAPx2_ASAP7_75t_R FILLER_61_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_859 ();
 DECAPx6_ASAP7_75t_R FILLER_61_866 ();
 FILLER_ASAP7_75t_R FILLER_61_880 ();
 FILLER_ASAP7_75t_R FILLER_61_888 ();
 DECAPx2_ASAP7_75t_R FILLER_61_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_902 ();
 FILLER_ASAP7_75t_R FILLER_61_923 ();
 DECAPx2_ASAP7_75t_R FILLER_61_927 ();
 FILLER_ASAP7_75t_R FILLER_61_941 ();
 DECAPx2_ASAP7_75t_R FILLER_61_949 ();
 FILLER_ASAP7_75t_R FILLER_61_962 ();
 DECAPx10_ASAP7_75t_R FILLER_61_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_989 ();
 DECAPx4_ASAP7_75t_R FILLER_61_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1006 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1015 ();
 FILLER_ASAP7_75t_R FILLER_61_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1094 ();
 FILLER_ASAP7_75t_R FILLER_61_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1132 ();
 FILLER_ASAP7_75t_R FILLER_61_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1144 ();
 FILLER_ASAP7_75t_R FILLER_61_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_61_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1167 ();
 FILLER_ASAP7_75t_R FILLER_61_1173 ();
 FILLER_ASAP7_75t_R FILLER_61_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1195 ();
 DECAPx4_ASAP7_75t_R FILLER_61_1209 ();
 FILLER_ASAP7_75t_R FILLER_61_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1231 ();
 FILLER_ASAP7_75t_R FILLER_61_1237 ();
 DECAPx4_ASAP7_75t_R FILLER_61_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_61_1277 ();
 DECAPx6_ASAP7_75t_R FILLER_61_1299 ();
 FILLER_ASAP7_75t_R FILLER_61_1313 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1327 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_1333 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1343 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_1349 ();
 DECAPx4_ASAP7_75t_R FILLER_61_1355 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_1365 ();
 DECAPx2_ASAP7_75t_R FILLER_61_1369 ();
 FILLER_ASAP7_75t_R FILLER_61_1375 ();
 DECAPx1_ASAP7_75t_R FILLER_62_2 ();
 DECAPx2_ASAP7_75t_R FILLER_62_12 ();
 FILLER_ASAP7_75t_R FILLER_62_25 ();
 FILLER_ASAP7_75t_R FILLER_62_34 ();
 DECAPx1_ASAP7_75t_R FILLER_62_39 ();
 DECAPx1_ASAP7_75t_R FILLER_62_51 ();
 FILLER_ASAP7_75t_R FILLER_62_61 ();
 FILLER_ASAP7_75t_R FILLER_62_71 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_79 ();
 FILLER_ASAP7_75t_R FILLER_62_88 ();
 DECAPx10_ASAP7_75t_R FILLER_62_96 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_118 ();
 DECAPx6_ASAP7_75t_R FILLER_62_124 ();
 DECAPx2_ASAP7_75t_R FILLER_62_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_144 ();
 FILLER_ASAP7_75t_R FILLER_62_151 ();
 DECAPx10_ASAP7_75t_R FILLER_62_156 ();
 DECAPx1_ASAP7_75t_R FILLER_62_178 ();
 FILLER_ASAP7_75t_R FILLER_62_188 ();
 DECAPx4_ASAP7_75t_R FILLER_62_193 ();
 FILLER_ASAP7_75t_R FILLER_62_203 ();
 FILLER_ASAP7_75t_R FILLER_62_211 ();
 DECAPx1_ASAP7_75t_R FILLER_62_219 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_226 ();
 DECAPx4_ASAP7_75t_R FILLER_62_235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_245 ();
 FILLER_ASAP7_75t_R FILLER_62_256 ();
 FILLER_ASAP7_75t_R FILLER_62_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_274 ();
 DECAPx2_ASAP7_75t_R FILLER_62_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_291 ();
 FILLER_ASAP7_75t_R FILLER_62_318 ();
 DECAPx6_ASAP7_75t_R FILLER_62_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_337 ();
 DECAPx4_ASAP7_75t_R FILLER_62_346 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_356 ();
 FILLER_ASAP7_75t_R FILLER_62_365 ();
 FILLER_ASAP7_75t_R FILLER_62_373 ();
 DECAPx6_ASAP7_75t_R FILLER_62_401 ();
 DECAPx2_ASAP7_75t_R FILLER_62_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_421 ();
 DECAPx10_ASAP7_75t_R FILLER_62_428 ();
 DECAPx1_ASAP7_75t_R FILLER_62_450 ();
 FILLER_ASAP7_75t_R FILLER_62_460 ();
 DECAPx10_ASAP7_75t_R FILLER_62_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_486 ();
 DECAPx10_ASAP7_75t_R FILLER_62_490 ();
 DECAPx6_ASAP7_75t_R FILLER_62_512 ();
 DECAPx1_ASAP7_75t_R FILLER_62_526 ();
 DECAPx1_ASAP7_75t_R FILLER_62_536 ();
 DECAPx6_ASAP7_75t_R FILLER_62_546 ();
 DECAPx6_ASAP7_75t_R FILLER_62_566 ();
 DECAPx1_ASAP7_75t_R FILLER_62_580 ();
 FILLER_ASAP7_75t_R FILLER_62_594 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_602 ();
 DECAPx10_ASAP7_75t_R FILLER_62_611 ();
 FILLER_ASAP7_75t_R FILLER_62_633 ();
 DECAPx6_ASAP7_75t_R FILLER_62_641 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_655 ();
 DECAPx6_ASAP7_75t_R FILLER_62_664 ();
 DECAPx1_ASAP7_75t_R FILLER_62_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_682 ();
 DECAPx10_ASAP7_75t_R FILLER_62_703 ();
 DECAPx4_ASAP7_75t_R FILLER_62_725 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_735 ();
 DECAPx6_ASAP7_75t_R FILLER_62_744 ();
 DECAPx4_ASAP7_75t_R FILLER_62_761 ();
 DECAPx2_ASAP7_75t_R FILLER_62_777 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_783 ();
 DECAPx6_ASAP7_75t_R FILLER_62_812 ();
 FILLER_ASAP7_75t_R FILLER_62_826 ();
 DECAPx6_ASAP7_75t_R FILLER_62_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_845 ();
 DECAPx2_ASAP7_75t_R FILLER_62_858 ();
 DECAPx10_ASAP7_75t_R FILLER_62_867 ();
 DECAPx6_ASAP7_75t_R FILLER_62_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_903 ();
 FILLER_ASAP7_75t_R FILLER_62_909 ();
 DECAPx2_ASAP7_75t_R FILLER_62_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_923 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_930 ();
 DECAPx10_ASAP7_75t_R FILLER_62_939 ();
 DECAPx10_ASAP7_75t_R FILLER_62_961 ();
 DECAPx1_ASAP7_75t_R FILLER_62_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_987 ();
 DECAPx4_ASAP7_75t_R FILLER_62_995 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_1005 ();
 FILLER_ASAP7_75t_R FILLER_62_1034 ();
 FILLER_ASAP7_75t_R FILLER_62_1042 ();
 DECAPx6_ASAP7_75t_R FILLER_62_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1068 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_62_1122 ();
 DECAPx4_ASAP7_75t_R FILLER_62_1138 ();
 FILLER_ASAP7_75t_R FILLER_62_1174 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_1182 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_1211 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_1240 ();
 DECAPx1_ASAP7_75t_R FILLER_62_1252 ();
 DECAPx4_ASAP7_75t_R FILLER_62_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1269 ();
 FILLER_ASAP7_75t_R FILLER_62_1278 ();
 DECAPx4_ASAP7_75t_R FILLER_62_1286 ();
 FILLER_ASAP7_75t_R FILLER_62_1296 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1306 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1321 ();
 DECAPx1_ASAP7_75t_R FILLER_62_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_1329 ();
 DECAPx6_ASAP7_75t_R FILLER_62_1337 ();
 DECAPx1_ASAP7_75t_R FILLER_62_1351 ();
 DECAPx1_ASAP7_75t_R FILLER_62_1362 ();
 DECAPx2_ASAP7_75t_R FILLER_62_1369 ();
 FILLER_ASAP7_75t_R FILLER_62_1375 ();
 DECAPx4_ASAP7_75t_R FILLER_63_2 ();
 FILLER_ASAP7_75t_R FILLER_63_12 ();
 FILLER_ASAP7_75t_R FILLER_63_17 ();
 FILLER_ASAP7_75t_R FILLER_63_25 ();
 FILLER_ASAP7_75t_R FILLER_63_34 ();
 FILLER_ASAP7_75t_R FILLER_63_43 ();
 DECAPx6_ASAP7_75t_R FILLER_63_51 ();
 DECAPx4_ASAP7_75t_R FILLER_63_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_81 ();
 DECAPx4_ASAP7_75t_R FILLER_63_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_118 ();
 DECAPx2_ASAP7_75t_R FILLER_63_125 ();
 FILLER_ASAP7_75t_R FILLER_63_131 ();
 DECAPx1_ASAP7_75t_R FILLER_63_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_163 ();
 DECAPx4_ASAP7_75t_R FILLER_63_172 ();
 FILLER_ASAP7_75t_R FILLER_63_182 ();
 FILLER_ASAP7_75t_R FILLER_63_190 ();
 FILLER_ASAP7_75t_R FILLER_63_198 ();
 DECAPx1_ASAP7_75t_R FILLER_63_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_207 ();
 DECAPx6_ASAP7_75t_R FILLER_63_234 ();
 DECAPx1_ASAP7_75t_R FILLER_63_248 ();
 DECAPx2_ASAP7_75t_R FILLER_63_258 ();
 FILLER_ASAP7_75t_R FILLER_63_264 ();
 DECAPx1_ASAP7_75t_R FILLER_63_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_276 ();
 DECAPx6_ASAP7_75t_R FILLER_63_285 ();
 FILLER_ASAP7_75t_R FILLER_63_305 ();
 DECAPx2_ASAP7_75t_R FILLER_63_310 ();
 DECAPx2_ASAP7_75t_R FILLER_63_322 ();
 FILLER_ASAP7_75t_R FILLER_63_334 ();
 FILLER_ASAP7_75t_R FILLER_63_342 ();
 FILLER_ASAP7_75t_R FILLER_63_352 ();
 DECAPx4_ASAP7_75t_R FILLER_63_361 ();
 DECAPx1_ASAP7_75t_R FILLER_63_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_378 ();
 DECAPx1_ASAP7_75t_R FILLER_63_385 ();
 FILLER_ASAP7_75t_R FILLER_63_395 ();
 DECAPx6_ASAP7_75t_R FILLER_63_400 ();
 DECAPx2_ASAP7_75t_R FILLER_63_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_446 ();
 DECAPx1_ASAP7_75t_R FILLER_63_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_477 ();
 DECAPx1_ASAP7_75t_R FILLER_63_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_488 ();
 FILLER_ASAP7_75t_R FILLER_63_515 ();
 DECAPx1_ASAP7_75t_R FILLER_63_523 ();
 DECAPx4_ASAP7_75t_R FILLER_63_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_563 ();
 DECAPx10_ASAP7_75t_R FILLER_63_574 ();
 DECAPx10_ASAP7_75t_R FILLER_63_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_618 ();
 FILLER_ASAP7_75t_R FILLER_63_625 ();
 FILLER_ASAP7_75t_R FILLER_63_633 ();
 DECAPx2_ASAP7_75t_R FILLER_63_642 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_648 ();
 DECAPx2_ASAP7_75t_R FILLER_63_657 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_663 ();
 DECAPx1_ASAP7_75t_R FILLER_63_672 ();
 DECAPx6_ASAP7_75t_R FILLER_63_683 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_697 ();
 DECAPx2_ASAP7_75t_R FILLER_63_706 ();
 FILLER_ASAP7_75t_R FILLER_63_712 ();
 FILLER_ASAP7_75t_R FILLER_63_721 ();
 DECAPx2_ASAP7_75t_R FILLER_63_729 ();
 FILLER_ASAP7_75t_R FILLER_63_735 ();
 FILLER_ASAP7_75t_R FILLER_63_763 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_772 ();
 FILLER_ASAP7_75t_R FILLER_63_782 ();
 DECAPx6_ASAP7_75t_R FILLER_63_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_804 ();
 FILLER_ASAP7_75t_R FILLER_63_825 ();
 FILLER_ASAP7_75t_R FILLER_63_834 ();
 DECAPx2_ASAP7_75t_R FILLER_63_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_848 ();
 DECAPx1_ASAP7_75t_R FILLER_63_856 ();
 FILLER_ASAP7_75t_R FILLER_63_866 ();
 DECAPx6_ASAP7_75t_R FILLER_63_877 ();
 FILLER_ASAP7_75t_R FILLER_63_891 ();
 FILLER_ASAP7_75t_R FILLER_63_899 ();
 FILLER_ASAP7_75t_R FILLER_63_907 ();
 DECAPx4_ASAP7_75t_R FILLER_63_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_922 ();
 DECAPx6_ASAP7_75t_R FILLER_63_927 ();
 DECAPx2_ASAP7_75t_R FILLER_63_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_947 ();
 FILLER_ASAP7_75t_R FILLER_63_954 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_962 ();
 DECAPx2_ASAP7_75t_R FILLER_63_975 ();
 FILLER_ASAP7_75t_R FILLER_63_993 ();
 DECAPx2_ASAP7_75t_R FILLER_63_1003 ();
 FILLER_ASAP7_75t_R FILLER_63_1015 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_63_1026 ();
 FILLER_ASAP7_75t_R FILLER_63_1039 ();
 FILLER_ASAP7_75t_R FILLER_63_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_63_1054 ();
 FILLER_ASAP7_75t_R FILLER_63_1060 ();
 FILLER_ASAP7_75t_R FILLER_63_1074 ();
 FILLER_ASAP7_75t_R FILLER_63_1083 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1099 ();
 DECAPx2_ASAP7_75t_R FILLER_63_1121 ();
 FILLER_ASAP7_75t_R FILLER_63_1127 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_63_1144 ();
 DECAPx6_ASAP7_75t_R FILLER_63_1166 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1180 ();
 DECAPx2_ASAP7_75t_R FILLER_63_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1207 ();
 FILLER_ASAP7_75t_R FILLER_63_1218 ();
 FILLER_ASAP7_75t_R FILLER_63_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1233 ();
 FILLER_ASAP7_75t_R FILLER_63_1240 ();
 DECAPx2_ASAP7_75t_R FILLER_63_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1285 ();
 FILLER_ASAP7_75t_R FILLER_63_1295 ();
 DECAPx4_ASAP7_75t_R FILLER_63_1323 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1333 ();
 DECAPx1_ASAP7_75t_R FILLER_63_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_1348 ();
 FILLER_ASAP7_75t_R FILLER_63_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_64_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_8 ();
 FILLER_ASAP7_75t_R FILLER_64_35 ();
 DECAPx6_ASAP7_75t_R FILLER_64_43 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_60 ();
 DECAPx4_ASAP7_75t_R FILLER_64_69 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_79 ();
 DECAPx2_ASAP7_75t_R FILLER_64_88 ();
 FILLER_ASAP7_75t_R FILLER_64_94 ();
 DECAPx2_ASAP7_75t_R FILLER_64_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_105 ();
 DECAPx2_ASAP7_75t_R FILLER_64_132 ();
 FILLER_ASAP7_75t_R FILLER_64_144 ();
 DECAPx1_ASAP7_75t_R FILLER_64_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_156 ();
 FILLER_ASAP7_75t_R FILLER_64_163 ();
 FILLER_ASAP7_75t_R FILLER_64_173 ();
 DECAPx1_ASAP7_75t_R FILLER_64_181 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_193 ();
 DECAPx10_ASAP7_75t_R FILLER_64_204 ();
 DECAPx10_ASAP7_75t_R FILLER_64_226 ();
 FILLER_ASAP7_75t_R FILLER_64_254 ();
 DECAPx6_ASAP7_75t_R FILLER_64_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_273 ();
 FILLER_ASAP7_75t_R FILLER_64_280 ();
 DECAPx10_ASAP7_75t_R FILLER_64_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_307 ();
 DECAPx1_ASAP7_75t_R FILLER_64_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_338 ();
 DECAPx10_ASAP7_75t_R FILLER_64_347 ();
 DECAPx10_ASAP7_75t_R FILLER_64_369 ();
 DECAPx2_ASAP7_75t_R FILLER_64_391 ();
 DECAPx2_ASAP7_75t_R FILLER_64_403 ();
 FILLER_ASAP7_75t_R FILLER_64_409 ();
 FILLER_ASAP7_75t_R FILLER_64_417 ();
 DECAPx1_ASAP7_75t_R FILLER_64_425 ();
 DECAPx6_ASAP7_75t_R FILLER_64_432 ();
 DECAPx1_ASAP7_75t_R FILLER_64_446 ();
 DECAPx2_ASAP7_75t_R FILLER_64_456 ();
 FILLER_ASAP7_75t_R FILLER_64_464 ();
 DECAPx1_ASAP7_75t_R FILLER_64_469 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_499 ();
 FILLER_ASAP7_75t_R FILLER_64_505 ();
 FILLER_ASAP7_75t_R FILLER_64_513 ();
 DECAPx10_ASAP7_75t_R FILLER_64_523 ();
 FILLER_ASAP7_75t_R FILLER_64_548 ();
 DECAPx4_ASAP7_75t_R FILLER_64_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_563 ();
 FILLER_ASAP7_75t_R FILLER_64_570 ();
 FILLER_ASAP7_75t_R FILLER_64_578 ();
 DECAPx2_ASAP7_75t_R FILLER_64_586 ();
 FILLER_ASAP7_75t_R FILLER_64_592 ();
 DECAPx2_ASAP7_75t_R FILLER_64_600 ();
 FILLER_ASAP7_75t_R FILLER_64_606 ();
 DECAPx6_ASAP7_75t_R FILLER_64_614 ();
 FILLER_ASAP7_75t_R FILLER_64_635 ();
 DECAPx10_ASAP7_75t_R FILLER_64_647 ();
 DECAPx2_ASAP7_75t_R FILLER_64_669 ();
 FILLER_ASAP7_75t_R FILLER_64_675 ();
 DECAPx2_ASAP7_75t_R FILLER_64_697 ();
 FILLER_ASAP7_75t_R FILLER_64_709 ();
 DECAPx6_ASAP7_75t_R FILLER_64_731 ();
 DECAPx2_ASAP7_75t_R FILLER_64_745 ();
 DECAPx2_ASAP7_75t_R FILLER_64_754 ();
 FILLER_ASAP7_75t_R FILLER_64_760 ();
 DECAPx2_ASAP7_75t_R FILLER_64_768 ();
 FILLER_ASAP7_75t_R FILLER_64_774 ();
 FILLER_ASAP7_75t_R FILLER_64_802 ();
 DECAPx2_ASAP7_75t_R FILLER_64_807 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_813 ();
 DECAPx2_ASAP7_75t_R FILLER_64_842 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_848 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_871 ();
 FILLER_ASAP7_75t_R FILLER_64_880 ();
 FILLER_ASAP7_75t_R FILLER_64_888 ();
 FILLER_ASAP7_75t_R FILLER_64_898 ();
 FILLER_ASAP7_75t_R FILLER_64_909 ();
 DECAPx6_ASAP7_75t_R FILLER_64_917 ();
 FILLER_ASAP7_75t_R FILLER_64_940 ();
 DECAPx1_ASAP7_75t_R FILLER_64_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_949 ();
 DECAPx2_ASAP7_75t_R FILLER_64_976 ();
 FILLER_ASAP7_75t_R FILLER_64_982 ();
 FILLER_ASAP7_75t_R FILLER_64_990 ();
 DECAPx10_ASAP7_75t_R FILLER_64_995 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1017 ();
 DECAPx4_ASAP7_75t_R FILLER_64_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_64_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_64_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1087 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_1093 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1122 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_1128 ();
 FILLER_ASAP7_75t_R FILLER_64_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1148 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_1154 ();
 FILLER_ASAP7_75t_R FILLER_64_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_64_1216 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1238 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_1244 ();
 DECAPx4_ASAP7_75t_R FILLER_64_1253 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_1263 ();
 FILLER_ASAP7_75t_R FILLER_64_1274 ();
 DECAPx6_ASAP7_75t_R FILLER_64_1302 ();
 FILLER_ASAP7_75t_R FILLER_64_1316 ();
 FILLER_ASAP7_75t_R FILLER_64_1344 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1349 ();
 FILLER_ASAP7_75t_R FILLER_64_1355 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_1363 ();
 DECAPx2_ASAP7_75t_R FILLER_64_1369 ();
 FILLER_ASAP7_75t_R FILLER_64_1375 ();
 DECAPx4_ASAP7_75t_R FILLER_65_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_12 ();
 FILLER_ASAP7_75t_R FILLER_65_21 ();
 DECAPx4_ASAP7_75t_R FILLER_65_26 ();
 FILLER_ASAP7_75t_R FILLER_65_36 ();
 DECAPx2_ASAP7_75t_R FILLER_65_44 ();
 DECAPx2_ASAP7_75t_R FILLER_65_56 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_62 ();
 DECAPx6_ASAP7_75t_R FILLER_65_71 ();
 DECAPx2_ASAP7_75t_R FILLER_65_85 ();
 DECAPx6_ASAP7_75t_R FILLER_65_97 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_117 ();
 DECAPx4_ASAP7_75t_R FILLER_65_123 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_159 ();
 DECAPx4_ASAP7_75t_R FILLER_65_168 ();
 FILLER_ASAP7_75t_R FILLER_65_178 ();
 FILLER_ASAP7_75t_R FILLER_65_187 ();
 DECAPx4_ASAP7_75t_R FILLER_65_197 ();
 FILLER_ASAP7_75t_R FILLER_65_207 ();
 DECAPx4_ASAP7_75t_R FILLER_65_217 ();
 FILLER_ASAP7_75t_R FILLER_65_233 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_261 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_290 ();
 FILLER_ASAP7_75t_R FILLER_65_299 ();
 DECAPx1_ASAP7_75t_R FILLER_65_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_311 ();
 DECAPx1_ASAP7_75t_R FILLER_65_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_322 ();
 DECAPx2_ASAP7_75t_R FILLER_65_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_332 ();
 FILLER_ASAP7_75t_R FILLER_65_336 ();
 DECAPx2_ASAP7_75t_R FILLER_65_344 ();
 DECAPx1_ASAP7_75t_R FILLER_65_376 ();
 DECAPx2_ASAP7_75t_R FILLER_65_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_392 ();
 DECAPx4_ASAP7_75t_R FILLER_65_419 ();
 FILLER_ASAP7_75t_R FILLER_65_429 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_438 ();
 DECAPx10_ASAP7_75t_R FILLER_65_447 ();
 DECAPx2_ASAP7_75t_R FILLER_65_469 ();
 DECAPx2_ASAP7_75t_R FILLER_65_481 ();
 FILLER_ASAP7_75t_R FILLER_65_493 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_501 ();
 DECAPx2_ASAP7_75t_R FILLER_65_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_513 ();
 DECAPx10_ASAP7_75t_R FILLER_65_522 ();
 DECAPx1_ASAP7_75t_R FILLER_65_544 ();
 DECAPx4_ASAP7_75t_R FILLER_65_554 ();
 DECAPx1_ASAP7_75t_R FILLER_65_570 ();
 DECAPx4_ASAP7_75t_R FILLER_65_580 ();
 FILLER_ASAP7_75t_R FILLER_65_597 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_605 ();
 FILLER_ASAP7_75t_R FILLER_65_618 ();
 DECAPx4_ASAP7_75t_R FILLER_65_628 ();
 FILLER_ASAP7_75t_R FILLER_65_638 ();
 FILLER_ASAP7_75t_R FILLER_65_648 ();
 FILLER_ASAP7_75t_R FILLER_65_658 ();
 DECAPx4_ASAP7_75t_R FILLER_65_668 ();
 FILLER_ASAP7_75t_R FILLER_65_678 ();
 DECAPx10_ASAP7_75t_R FILLER_65_686 ();
 DECAPx4_ASAP7_75t_R FILLER_65_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_718 ();
 FILLER_ASAP7_75t_R FILLER_65_725 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_733 ();
 DECAPx10_ASAP7_75t_R FILLER_65_743 ();
 DECAPx4_ASAP7_75t_R FILLER_65_765 ();
 FILLER_ASAP7_75t_R FILLER_65_775 ();
 DECAPx2_ASAP7_75t_R FILLER_65_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_789 ();
 DECAPx6_ASAP7_75t_R FILLER_65_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_807 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_822 ();
 FILLER_ASAP7_75t_R FILLER_65_831 ();
 DECAPx4_ASAP7_75t_R FILLER_65_836 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_846 ();
 DECAPx4_ASAP7_75t_R FILLER_65_855 ();
 DECAPx10_ASAP7_75t_R FILLER_65_869 ();
 FILLER_ASAP7_75t_R FILLER_65_891 ();
 DECAPx4_ASAP7_75t_R FILLER_65_901 ();
 DECAPx2_ASAP7_75t_R FILLER_65_919 ();
 FILLER_ASAP7_75t_R FILLER_65_927 ();
 FILLER_ASAP7_75t_R FILLER_65_935 ();
 DECAPx2_ASAP7_75t_R FILLER_65_943 ();
 FILLER_ASAP7_75t_R FILLER_65_949 ();
 DECAPx2_ASAP7_75t_R FILLER_65_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_960 ();
 FILLER_ASAP7_75t_R FILLER_65_969 ();
 DECAPx6_ASAP7_75t_R FILLER_65_974 ();
 FILLER_ASAP7_75t_R FILLER_65_988 ();
 DECAPx1_ASAP7_75t_R FILLER_65_999 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_1006 ();
 FILLER_ASAP7_75t_R FILLER_65_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1024 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_1030 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1040 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_1046 ();
 DECAPx1_ASAP7_75t_R FILLER_65_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1079 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1094 ();
 FILLER_ASAP7_75t_R FILLER_65_1103 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_1137 ();
 DECAPx1_ASAP7_75t_R FILLER_65_1142 ();
 FILLER_ASAP7_75t_R FILLER_65_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1180 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_1186 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_1199 ();
 FILLER_ASAP7_75t_R FILLER_65_1205 ();
 DECAPx6_ASAP7_75t_R FILLER_65_1217 ();
 DECAPx1_ASAP7_75t_R FILLER_65_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_65_1242 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1264 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_1270 ();
 DECAPx2_ASAP7_75t_R FILLER_65_1283 ();
 FILLER_ASAP7_75t_R FILLER_65_1289 ();
 DECAPx1_ASAP7_75t_R FILLER_65_1294 ();
 DECAPx4_ASAP7_75t_R FILLER_65_1301 ();
 FILLER_ASAP7_75t_R FILLER_65_1311 ();
 DECAPx4_ASAP7_75t_R FILLER_65_1323 ();
 DECAPx4_ASAP7_75t_R FILLER_65_1336 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_1346 ();
 FILLER_ASAP7_75t_R FILLER_65_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_66_2 ();
 DECAPx2_ASAP7_75t_R FILLER_66_24 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_30 ();
 DECAPx2_ASAP7_75t_R FILLER_66_59 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_65 ();
 FILLER_ASAP7_75t_R FILLER_66_74 ();
 DECAPx2_ASAP7_75t_R FILLER_66_79 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_85 ();
 DECAPx2_ASAP7_75t_R FILLER_66_114 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_120 ();
 DECAPx6_ASAP7_75t_R FILLER_66_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_143 ();
 FILLER_ASAP7_75t_R FILLER_66_150 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_155 ();
 DECAPx10_ASAP7_75t_R FILLER_66_161 ();
 DECAPx6_ASAP7_75t_R FILLER_66_183 ();
 FILLER_ASAP7_75t_R FILLER_66_203 ();
 FILLER_ASAP7_75t_R FILLER_66_211 ();
 FILLER_ASAP7_75t_R FILLER_66_239 ();
 FILLER_ASAP7_75t_R FILLER_66_247 ();
 DECAPx6_ASAP7_75t_R FILLER_66_252 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_266 ();
 DECAPx1_ASAP7_75t_R FILLER_66_275 ();
 DECAPx2_ASAP7_75t_R FILLER_66_282 ();
 DECAPx4_ASAP7_75t_R FILLER_66_314 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_324 ();
 DECAPx6_ASAP7_75t_R FILLER_66_333 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_347 ();
 FILLER_ASAP7_75t_R FILLER_66_356 ();
 FILLER_ASAP7_75t_R FILLER_66_364 ();
 DECAPx6_ASAP7_75t_R FILLER_66_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_406 ();
 DECAPx1_ASAP7_75t_R FILLER_66_410 ();
 DECAPx4_ASAP7_75t_R FILLER_66_417 ();
 FILLER_ASAP7_75t_R FILLER_66_427 ();
 FILLER_ASAP7_75t_R FILLER_66_455 ();
 FILLER_ASAP7_75t_R FILLER_66_460 ();
 DECAPx2_ASAP7_75t_R FILLER_66_464 ();
 DECAPx10_ASAP7_75t_R FILLER_66_476 ();
 DECAPx4_ASAP7_75t_R FILLER_66_498 ();
 FILLER_ASAP7_75t_R FILLER_66_508 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_516 ();
 FILLER_ASAP7_75t_R FILLER_66_525 ();
 FILLER_ASAP7_75t_R FILLER_66_533 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_541 ();
 FILLER_ASAP7_75t_R FILLER_66_552 ();
 DECAPx6_ASAP7_75t_R FILLER_66_562 ();
 DECAPx1_ASAP7_75t_R FILLER_66_576 ();
 DECAPx2_ASAP7_75t_R FILLER_66_586 ();
 FILLER_ASAP7_75t_R FILLER_66_592 ();
 FILLER_ASAP7_75t_R FILLER_66_604 ();
 FILLER_ASAP7_75t_R FILLER_66_612 ();
 FILLER_ASAP7_75t_R FILLER_66_620 ();
 DECAPx10_ASAP7_75t_R FILLER_66_628 ();
 DECAPx2_ASAP7_75t_R FILLER_66_650 ();
 FILLER_ASAP7_75t_R FILLER_66_656 ();
 DECAPx10_ASAP7_75t_R FILLER_66_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_700 ();
 DECAPx10_ASAP7_75t_R FILLER_66_708 ();
 DECAPx2_ASAP7_75t_R FILLER_66_730 ();
 FILLER_ASAP7_75t_R FILLER_66_756 ();
 DECAPx4_ASAP7_75t_R FILLER_66_764 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_774 ();
 DECAPx4_ASAP7_75t_R FILLER_66_797 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_807 ();
 DECAPx6_ASAP7_75t_R FILLER_66_817 ();
 DECAPx1_ASAP7_75t_R FILLER_66_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_835 ();
 DECAPx2_ASAP7_75t_R FILLER_66_839 ();
 FILLER_ASAP7_75t_R FILLER_66_845 ();
 DECAPx6_ASAP7_75t_R FILLER_66_854 ();
 DECAPx1_ASAP7_75t_R FILLER_66_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_872 ();
 DECAPx2_ASAP7_75t_R FILLER_66_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_885 ();
 DECAPx6_ASAP7_75t_R FILLER_66_896 ();
 DECAPx1_ASAP7_75t_R FILLER_66_910 ();
 DECAPx4_ASAP7_75t_R FILLER_66_920 ();
 FILLER_ASAP7_75t_R FILLER_66_930 ();
 DECAPx10_ASAP7_75t_R FILLER_66_940 ();
 DECAPx2_ASAP7_75t_R FILLER_66_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_968 ();
 DECAPx6_ASAP7_75t_R FILLER_66_975 ();
 FILLER_ASAP7_75t_R FILLER_66_989 ();
 FILLER_ASAP7_75t_R FILLER_66_997 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1005 ();
 FILLER_ASAP7_75t_R FILLER_66_1029 ();
 FILLER_ASAP7_75t_R FILLER_66_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_66_1055 ();
 FILLER_ASAP7_75t_R FILLER_66_1061 ();
 DECAPx4_ASAP7_75t_R FILLER_66_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_66_1083 ();
 FILLER_ASAP7_75t_R FILLER_66_1105 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1119 ();
 DECAPx6_ASAP7_75t_R FILLER_66_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1137 ();
 DECAPx4_ASAP7_75t_R FILLER_66_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1154 ();
 DECAPx2_ASAP7_75t_R FILLER_66_1161 ();
 FILLER_ASAP7_75t_R FILLER_66_1167 ();
 FILLER_ASAP7_75t_R FILLER_66_1189 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1221 ();
 FILLER_ASAP7_75t_R FILLER_66_1226 ();
 DECAPx2_ASAP7_75t_R FILLER_66_1237 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_1243 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1255 ();
 DECAPx4_ASAP7_75t_R FILLER_66_1269 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_1279 ();
 DECAPx1_ASAP7_75t_R FILLER_66_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1312 ();
 DECAPx4_ASAP7_75t_R FILLER_66_1323 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_1333 ();
 DECAPx4_ASAP7_75t_R FILLER_66_1344 ();
 FILLER_ASAP7_75t_R FILLER_66_1354 ();
 FILLER_ASAP7_75t_R FILLER_66_1363 ();
 DECAPx2_ASAP7_75t_R FILLER_66_1371 ();
 DECAPx10_ASAP7_75t_R FILLER_67_2 ();
 DECAPx10_ASAP7_75t_R FILLER_67_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_46 ();
 DECAPx4_ASAP7_75t_R FILLER_67_50 ();
 FILLER_ASAP7_75t_R FILLER_67_60 ();
 DECAPx2_ASAP7_75t_R FILLER_67_88 ();
 FILLER_ASAP7_75t_R FILLER_67_94 ();
 FILLER_ASAP7_75t_R FILLER_67_102 ();
 DECAPx2_ASAP7_75t_R FILLER_67_107 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_67_113 ();
 DECAPx1_ASAP7_75t_R FILLER_67_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_123 ();
 FILLER_ASAP7_75t_R FILLER_67_132 ();
 DECAPx6_ASAP7_75t_R FILLER_67_140 ();
 DECAPx2_ASAP7_75t_R FILLER_67_160 ();
 FILLER_ASAP7_75t_R FILLER_67_166 ();
 FILLER_ASAP7_75t_R FILLER_67_174 ();
 DECAPx2_ASAP7_75t_R FILLER_67_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_190 ();
 DECAPx4_ASAP7_75t_R FILLER_67_197 ();
 DECAPx4_ASAP7_75t_R FILLER_67_210 ();
 FILLER_ASAP7_75t_R FILLER_67_226 ();
 FILLER_ASAP7_75t_R FILLER_67_231 ();
 DECAPx10_ASAP7_75t_R FILLER_67_236 ();
 DECAPx10_ASAP7_75t_R FILLER_67_258 ();
 DECAPx10_ASAP7_75t_R FILLER_67_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_302 ();
 DECAPx4_ASAP7_75t_R FILLER_67_306 ();
 FILLER_ASAP7_75t_R FILLER_67_316 ();
 DECAPx6_ASAP7_75t_R FILLER_67_344 ();
 DECAPx2_ASAP7_75t_R FILLER_67_358 ();
 DECAPx2_ASAP7_75t_R FILLER_67_367 ();
 DECAPx2_ASAP7_75t_R FILLER_67_379 ();
 FILLER_ASAP7_75t_R FILLER_67_388 ();
 DECAPx1_ASAP7_75t_R FILLER_67_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_397 ();
 DECAPx4_ASAP7_75t_R FILLER_67_424 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_67_440 ();
 DECAPx4_ASAP7_75t_R FILLER_67_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_456 ();
 DECAPx1_ASAP7_75t_R FILLER_67_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_487 ();
 DECAPx2_ASAP7_75t_R FILLER_67_498 ();
 FILLER_ASAP7_75t_R FILLER_67_507 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_67_515 ();
 FILLER_ASAP7_75t_R FILLER_67_536 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_67_544 ();
 DECAPx4_ASAP7_75t_R FILLER_67_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_563 ();
 DECAPx10_ASAP7_75t_R FILLER_67_571 ();
 DECAPx10_ASAP7_75t_R FILLER_67_593 ();
 DECAPx4_ASAP7_75t_R FILLER_67_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_625 ();
 DECAPx4_ASAP7_75t_R FILLER_67_633 ();
 DECAPx10_ASAP7_75t_R FILLER_67_650 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_67_672 ();
 DECAPx6_ASAP7_75t_R FILLER_67_682 ();
 FILLER_ASAP7_75t_R FILLER_67_702 ();
 DECAPx6_ASAP7_75t_R FILLER_67_724 ();
 DECAPx1_ASAP7_75t_R FILLER_67_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_742 ();
 FILLER_ASAP7_75t_R FILLER_67_749 ();
 DECAPx2_ASAP7_75t_R FILLER_67_757 ();
 DECAPx4_ASAP7_75t_R FILLER_67_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_780 ();
 DECAPx6_ASAP7_75t_R FILLER_67_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_798 ();
 FILLER_ASAP7_75t_R FILLER_67_802 ();
 DECAPx2_ASAP7_75t_R FILLER_67_816 ();
 FILLER_ASAP7_75t_R FILLER_67_834 ();
 DECAPx1_ASAP7_75t_R FILLER_67_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_846 ();
 DECAPx2_ASAP7_75t_R FILLER_67_867 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_67_873 ();
 FILLER_ASAP7_75t_R FILLER_67_883 ();
 DECAPx6_ASAP7_75t_R FILLER_67_897 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_67_911 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_67_922 ();
 DECAPx6_ASAP7_75t_R FILLER_67_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_941 ();
 FILLER_ASAP7_75t_R FILLER_67_954 ();
 DECAPx1_ASAP7_75t_R FILLER_67_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_966 ();
 DECAPx1_ASAP7_75t_R FILLER_67_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_981 ();
 DECAPx10_ASAP7_75t_R FILLER_67_985 ();
 DECAPx6_ASAP7_75t_R FILLER_67_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_67_1034 ();
 DECAPx4_ASAP7_75t_R FILLER_67_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1082 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_67_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1101 ();
 FILLER_ASAP7_75t_R FILLER_67_1119 ();
 DECAPx1_ASAP7_75t_R FILLER_67_1131 ();
 DECAPx6_ASAP7_75t_R FILLER_67_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1158 ();
 DECAPx1_ASAP7_75t_R FILLER_67_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1173 ();
 FILLER_ASAP7_75t_R FILLER_67_1182 ();
 DECAPx1_ASAP7_75t_R FILLER_67_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_67_1198 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_67_1204 ();
 DECAPx6_ASAP7_75t_R FILLER_67_1214 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_1228 ();
 FILLER_ASAP7_75t_R FILLER_67_1241 ();
 DECAPx1_ASAP7_75t_R FILLER_67_1249 ();
 FILLER_ASAP7_75t_R FILLER_67_1279 ();
 DECAPx4_ASAP7_75t_R FILLER_67_1284 ();
 FILLER_ASAP7_75t_R FILLER_67_1294 ();
 DECAPx1_ASAP7_75t_R FILLER_67_1299 ();
 FILLER_ASAP7_75t_R FILLER_67_1315 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_67_1343 ();
 FILLER_ASAP7_75t_R FILLER_67_1351 ();
 FILLER_ASAP7_75t_R FILLER_67_1360 ();
 FILLER_ASAP7_75t_R FILLER_67_1368 ();
 FILLER_ASAP7_75t_R FILLER_67_1375 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_2 ();
 FILLER_ASAP7_75t_R FILLER_68_31 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_36 ();
 DECAPx1_ASAP7_75t_R FILLER_68_42 ();
 DECAPx10_ASAP7_75t_R FILLER_68_52 ();
 DECAPx10_ASAP7_75t_R FILLER_68_74 ();
 DECAPx2_ASAP7_75t_R FILLER_68_96 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_102 ();
 DECAPx6_ASAP7_75t_R FILLER_68_111 ();
 FILLER_ASAP7_75t_R FILLER_68_125 ();
 DECAPx2_ASAP7_75t_R FILLER_68_135 ();
 FILLER_ASAP7_75t_R FILLER_68_141 ();
 FILLER_ASAP7_75t_R FILLER_68_169 ();
 FILLER_ASAP7_75t_R FILLER_68_193 ();
 DECAPx10_ASAP7_75t_R FILLER_68_201 ();
 DECAPx10_ASAP7_75t_R FILLER_68_223 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_245 ();
 FILLER_ASAP7_75t_R FILLER_68_254 ();
 DECAPx10_ASAP7_75t_R FILLER_68_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_287 ();
 DECAPx1_ASAP7_75t_R FILLER_68_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_298 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_302 ();
 DECAPx4_ASAP7_75t_R FILLER_68_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_321 ();
 FILLER_ASAP7_75t_R FILLER_68_328 ();
 FILLER_ASAP7_75t_R FILLER_68_333 ();
 DECAPx10_ASAP7_75t_R FILLER_68_341 ();
 DECAPx6_ASAP7_75t_R FILLER_68_363 ();
 DECAPx1_ASAP7_75t_R FILLER_68_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_381 ();
 DECAPx2_ASAP7_75t_R FILLER_68_404 ();
 FILLER_ASAP7_75t_R FILLER_68_410 ();
 FILLER_ASAP7_75t_R FILLER_68_418 ();
 DECAPx10_ASAP7_75t_R FILLER_68_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_445 ();
 DECAPx4_ASAP7_75t_R FILLER_68_452 ();
 FILLER_ASAP7_75t_R FILLER_68_464 ();
 FILLER_ASAP7_75t_R FILLER_68_472 ();
 DECAPx2_ASAP7_75t_R FILLER_68_477 ();
 FILLER_ASAP7_75t_R FILLER_68_509 ();
 DECAPx6_ASAP7_75t_R FILLER_68_533 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_547 ();
 DECAPx2_ASAP7_75t_R FILLER_68_556 ();
 FILLER_ASAP7_75t_R FILLER_68_562 ();
 DECAPx6_ASAP7_75t_R FILLER_68_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_598 ();
 DECAPx6_ASAP7_75t_R FILLER_68_606 ();
 FILLER_ASAP7_75t_R FILLER_68_620 ();
 FILLER_ASAP7_75t_R FILLER_68_642 ();
 DECAPx4_ASAP7_75t_R FILLER_68_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_674 ();
 DECAPx4_ASAP7_75t_R FILLER_68_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_705 ();
 FILLER_ASAP7_75t_R FILLER_68_712 ();
 DECAPx4_ASAP7_75t_R FILLER_68_721 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_731 ();
 DECAPx6_ASAP7_75t_R FILLER_68_740 ();
 DECAPx1_ASAP7_75t_R FILLER_68_754 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_784 ();
 DECAPx1_ASAP7_75t_R FILLER_68_813 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_831 ();
 DECAPx2_ASAP7_75t_R FILLER_68_840 ();
 FILLER_ASAP7_75t_R FILLER_68_846 ();
 DECAPx2_ASAP7_75t_R FILLER_68_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_860 ();
 DECAPx10_ASAP7_75t_R FILLER_68_868 ();
 DECAPx2_ASAP7_75t_R FILLER_68_890 ();
 FILLER_ASAP7_75t_R FILLER_68_896 ();
 DECAPx4_ASAP7_75t_R FILLER_68_906 ();
 DECAPx1_ASAP7_75t_R FILLER_68_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_928 ();
 DECAPx4_ASAP7_75t_R FILLER_68_932 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_942 ();
 DECAPx2_ASAP7_75t_R FILLER_68_948 ();
 FILLER_ASAP7_75t_R FILLER_68_954 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_964 ();
 DECAPx4_ASAP7_75t_R FILLER_68_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1003 ();
 DECAPx4_ASAP7_75t_R FILLER_68_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1040 ();
 DECAPx1_ASAP7_75t_R FILLER_68_1044 ();
 DECAPx4_ASAP7_75t_R FILLER_68_1058 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_1068 ();
 FILLER_ASAP7_75t_R FILLER_68_1081 ();
 DECAPx4_ASAP7_75t_R FILLER_68_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1119 ();
 FILLER_ASAP7_75t_R FILLER_68_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_68_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1230 ();
 FILLER_ASAP7_75t_R FILLER_68_1258 ();
 DECAPx1_ASAP7_75t_R FILLER_68_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1267 ();
 DECAPx6_ASAP7_75t_R FILLER_68_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1285 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1293 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_68_1305 ();
 DECAPx1_ASAP7_75t_R FILLER_68_1327 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_1331 ();
 FILLER_ASAP7_75t_R FILLER_68_1335 ();
 DECAPx2_ASAP7_75t_R FILLER_68_1340 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_1346 ();
 FILLER_ASAP7_75t_R FILLER_68_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_69_2 ();
 FILLER_ASAP7_75t_R FILLER_69_14 ();
 FILLER_ASAP7_75t_R FILLER_69_22 ();
 FILLER_ASAP7_75t_R FILLER_69_50 ();
 DECAPx2_ASAP7_75t_R FILLER_69_60 ();
 FILLER_ASAP7_75t_R FILLER_69_66 ();
 FILLER_ASAP7_75t_R FILLER_69_76 ();
 DECAPx4_ASAP7_75t_R FILLER_69_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_91 ();
 DECAPx10_ASAP7_75t_R FILLER_69_118 ();
 DECAPx2_ASAP7_75t_R FILLER_69_140 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_146 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_155 ();
 DECAPx1_ASAP7_75t_R FILLER_69_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_165 ();
 FILLER_ASAP7_75t_R FILLER_69_169 ();
 FILLER_ASAP7_75t_R FILLER_69_179 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_187 ();
 DECAPx6_ASAP7_75t_R FILLER_69_216 ();
 DECAPx1_ASAP7_75t_R FILLER_69_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_234 ();
 FILLER_ASAP7_75t_R FILLER_69_243 ();
 FILLER_ASAP7_75t_R FILLER_69_251 ();
 DECAPx6_ASAP7_75t_R FILLER_69_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_273 ();
 DECAPx1_ASAP7_75t_R FILLER_69_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_304 ();
 FILLER_ASAP7_75t_R FILLER_69_313 ();
 DECAPx2_ASAP7_75t_R FILLER_69_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_327 ();
 DECAPx2_ASAP7_75t_R FILLER_69_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_360 ();
 DECAPx4_ASAP7_75t_R FILLER_69_369 ();
 FILLER_ASAP7_75t_R FILLER_69_385 ();
 FILLER_ASAP7_75t_R FILLER_69_393 ();
 FILLER_ASAP7_75t_R FILLER_69_401 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_409 ();
 FILLER_ASAP7_75t_R FILLER_69_420 ();
 DECAPx2_ASAP7_75t_R FILLER_69_428 ();
 FILLER_ASAP7_75t_R FILLER_69_440 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_445 ();
 DECAPx6_ASAP7_75t_R FILLER_69_456 ();
 FILLER_ASAP7_75t_R FILLER_69_470 ();
 DECAPx2_ASAP7_75t_R FILLER_69_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_484 ();
 FILLER_ASAP7_75t_R FILLER_69_491 ();
 DECAPx1_ASAP7_75t_R FILLER_69_499 ();
 FILLER_ASAP7_75t_R FILLER_69_509 ();
 FILLER_ASAP7_75t_R FILLER_69_519 ();
 DECAPx2_ASAP7_75t_R FILLER_69_529 ();
 FILLER_ASAP7_75t_R FILLER_69_535 ();
 FILLER_ASAP7_75t_R FILLER_69_543 ();
 DECAPx2_ASAP7_75t_R FILLER_69_571 ();
 FILLER_ASAP7_75t_R FILLER_69_581 ();
 FILLER_ASAP7_75t_R FILLER_69_590 ();
 FILLER_ASAP7_75t_R FILLER_69_598 ();
 DECAPx10_ASAP7_75t_R FILLER_69_620 ();
 DECAPx4_ASAP7_75t_R FILLER_69_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_652 ();
 FILLER_ASAP7_75t_R FILLER_69_681 ();
 DECAPx2_ASAP7_75t_R FILLER_69_689 ();
 FILLER_ASAP7_75t_R FILLER_69_701 ();
 DECAPx1_ASAP7_75t_R FILLER_69_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_713 ();
 FILLER_ASAP7_75t_R FILLER_69_734 ();
 DECAPx6_ASAP7_75t_R FILLER_69_742 ();
 DECAPx2_ASAP7_75t_R FILLER_69_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_762 ();
 DECAPx1_ASAP7_75t_R FILLER_69_769 ();
 DECAPx1_ASAP7_75t_R FILLER_69_776 ();
 DECAPx4_ASAP7_75t_R FILLER_69_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_793 ();
 FILLER_ASAP7_75t_R FILLER_69_801 ();
 DECAPx1_ASAP7_75t_R FILLER_69_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_813 ();
 DECAPx2_ASAP7_75t_R FILLER_69_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_825 ();
 DECAPx1_ASAP7_75t_R FILLER_69_838 ();
 DECAPx4_ASAP7_75t_R FILLER_69_849 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_859 ();
 FILLER_ASAP7_75t_R FILLER_69_882 ();
 DECAPx6_ASAP7_75t_R FILLER_69_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_904 ();
 DECAPx4_ASAP7_75t_R FILLER_69_915 ();
 FILLER_ASAP7_75t_R FILLER_69_927 ();
 DECAPx1_ASAP7_75t_R FILLER_69_937 ();
 FILLER_ASAP7_75t_R FILLER_69_950 ();
 DECAPx1_ASAP7_75t_R FILLER_69_958 ();
 DECAPx2_ASAP7_75t_R FILLER_69_968 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_974 ();
 DECAPx2_ASAP7_75t_R FILLER_69_983 ();
 DECAPx1_ASAP7_75t_R FILLER_69_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_69_1022 ();
 FILLER_ASAP7_75t_R FILLER_69_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1068 ();
 DECAPx6_ASAP7_75t_R FILLER_69_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_69_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1100 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_1106 ();
 FILLER_ASAP7_75t_R FILLER_69_1119 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1129 ();
 FILLER_ASAP7_75t_R FILLER_69_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1175 ();
 FILLER_ASAP7_75t_R FILLER_69_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1201 ();
 FILLER_ASAP7_75t_R FILLER_69_1207 ();
 DECAPx6_ASAP7_75t_R FILLER_69_1215 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1238 ();
 DECAPx4_ASAP7_75t_R FILLER_69_1260 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_1270 ();
 DECAPx4_ASAP7_75t_R FILLER_69_1276 ();
 FILLER_ASAP7_75t_R FILLER_69_1286 ();
 FILLER_ASAP7_75t_R FILLER_69_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_69_1319 ();
 DECAPx2_ASAP7_75t_R FILLER_69_1341 ();
 FILLER_ASAP7_75t_R FILLER_69_1347 ();
 FILLER_ASAP7_75t_R FILLER_69_1356 ();
 FILLER_ASAP7_75t_R FILLER_69_1361 ();
 FILLER_ASAP7_75t_R FILLER_69_1368 ();
 FILLER_ASAP7_75t_R FILLER_69_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_70_2 ();
 DECAPx2_ASAP7_75t_R FILLER_70_14 ();
 DECAPx1_ASAP7_75t_R FILLER_70_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_27 ();
 DECAPx4_ASAP7_75t_R FILLER_70_34 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_44 ();
 DECAPx2_ASAP7_75t_R FILLER_70_55 ();
 FILLER_ASAP7_75t_R FILLER_70_67 ();
 DECAPx2_ASAP7_75t_R FILLER_70_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_81 ();
 FILLER_ASAP7_75t_R FILLER_70_88 ();
 FILLER_ASAP7_75t_R FILLER_70_96 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_104 ();
 DECAPx2_ASAP7_75t_R FILLER_70_110 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_116 ();
 DECAPx2_ASAP7_75t_R FILLER_70_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_128 ();
 DECAPx10_ASAP7_75t_R FILLER_70_135 ();
 DECAPx6_ASAP7_75t_R FILLER_70_157 ();
 DECAPx1_ASAP7_75t_R FILLER_70_171 ();
 DECAPx4_ASAP7_75t_R FILLER_70_181 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_191 ();
 DECAPx1_ASAP7_75t_R FILLER_70_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_204 ();
 DECAPx2_ASAP7_75t_R FILLER_70_208 ();
 FILLER_ASAP7_75t_R FILLER_70_214 ();
 DECAPx1_ASAP7_75t_R FILLER_70_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_226 ();
 FILLER_ASAP7_75t_R FILLER_70_233 ();
 DECAPx1_ASAP7_75t_R FILLER_70_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_247 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_254 ();
 FILLER_ASAP7_75t_R FILLER_70_265 ();
 FILLER_ASAP7_75t_R FILLER_70_281 ();
 FILLER_ASAP7_75t_R FILLER_70_289 ();
 DECAPx4_ASAP7_75t_R FILLER_70_294 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_304 ();
 DECAPx10_ASAP7_75t_R FILLER_70_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_337 ();
 FILLER_ASAP7_75t_R FILLER_70_341 ();
 DECAPx1_ASAP7_75t_R FILLER_70_349 ();
 FILLER_ASAP7_75t_R FILLER_70_359 ();
 FILLER_ASAP7_75t_R FILLER_70_369 ();
 FILLER_ASAP7_75t_R FILLER_70_386 ();
 DECAPx2_ASAP7_75t_R FILLER_70_403 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_409 ();
 DECAPx2_ASAP7_75t_R FILLER_70_420 ();
 FILLER_ASAP7_75t_R FILLER_70_452 ();
 FILLER_ASAP7_75t_R FILLER_70_460 ();
 DECAPx2_ASAP7_75t_R FILLER_70_464 ();
 FILLER_ASAP7_75t_R FILLER_70_478 ();
 DECAPx4_ASAP7_75t_R FILLER_70_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_496 ();
 DECAPx6_ASAP7_75t_R FILLER_70_500 ();
 FILLER_ASAP7_75t_R FILLER_70_520 ();
 FILLER_ASAP7_75t_R FILLER_70_528 ();
 DECAPx1_ASAP7_75t_R FILLER_70_544 ();
 FILLER_ASAP7_75t_R FILLER_70_560 ();
 FILLER_ASAP7_75t_R FILLER_70_565 ();
 DECAPx2_ASAP7_75t_R FILLER_70_574 ();
 FILLER_ASAP7_75t_R FILLER_70_580 ();
 DECAPx4_ASAP7_75t_R FILLER_70_602 ();
 FILLER_ASAP7_75t_R FILLER_70_612 ();
 DECAPx6_ASAP7_75t_R FILLER_70_622 ();
 DECAPx10_ASAP7_75t_R FILLER_70_643 ();
 FILLER_ASAP7_75t_R FILLER_70_665 ();
 DECAPx1_ASAP7_75t_R FILLER_70_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_691 ();
 DECAPx2_ASAP7_75t_R FILLER_70_698 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_704 ();
 DECAPx2_ASAP7_75t_R FILLER_70_714 ();
 FILLER_ASAP7_75t_R FILLER_70_720 ();
 DECAPx4_ASAP7_75t_R FILLER_70_728 ();
 FILLER_ASAP7_75t_R FILLER_70_738 ();
 DECAPx2_ASAP7_75t_R FILLER_70_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_752 ();
 FILLER_ASAP7_75t_R FILLER_70_759 ();
 DECAPx10_ASAP7_75t_R FILLER_70_767 ();
 DECAPx4_ASAP7_75t_R FILLER_70_789 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_799 ();
 DECAPx10_ASAP7_75t_R FILLER_70_805 ();
 DECAPx6_ASAP7_75t_R FILLER_70_827 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_841 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_852 ();
 FILLER_ASAP7_75t_R FILLER_70_858 ();
 DECAPx4_ASAP7_75t_R FILLER_70_866 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_876 ();
 FILLER_ASAP7_75t_R FILLER_70_883 ();
 DECAPx4_ASAP7_75t_R FILLER_70_892 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_902 ();
 DECAPx10_ASAP7_75t_R FILLER_70_911 ();
 DECAPx4_ASAP7_75t_R FILLER_70_933 ();
 DECAPx4_ASAP7_75t_R FILLER_70_949 ();
 FILLER_ASAP7_75t_R FILLER_70_973 ();
 FILLER_ASAP7_75t_R FILLER_70_989 ();
 DECAPx2_ASAP7_75t_R FILLER_70_994 ();
 FILLER_ASAP7_75t_R FILLER_70_1003 ();
 DECAPx4_ASAP7_75t_R FILLER_70_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_70_1035 ();
 FILLER_ASAP7_75t_R FILLER_70_1045 ();
 FILLER_ASAP7_75t_R FILLER_70_1054 ();
 FILLER_ASAP7_75t_R FILLER_70_1062 ();
 FILLER_ASAP7_75t_R FILLER_70_1070 ();
 DECAPx6_ASAP7_75t_R FILLER_70_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1097 ();
 FILLER_ASAP7_75t_R FILLER_70_1103 ();
 DECAPx6_ASAP7_75t_R FILLER_70_1115 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_1129 ();
 FILLER_ASAP7_75t_R FILLER_70_1158 ();
 FILLER_ASAP7_75t_R FILLER_70_1186 ();
 FILLER_ASAP7_75t_R FILLER_70_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1206 ();
 DECAPx4_ASAP7_75t_R FILLER_70_1218 ();
 DECAPx2_ASAP7_75t_R FILLER_70_1234 ();
 FILLER_ASAP7_75t_R FILLER_70_1248 ();
 FILLER_ASAP7_75t_R FILLER_70_1253 ();
 DECAPx1_ASAP7_75t_R FILLER_70_1281 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1285 ();
 DECAPx1_ASAP7_75t_R FILLER_70_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_1296 ();
 DECAPx1_ASAP7_75t_R FILLER_70_1323 ();
 FILLER_ASAP7_75t_R FILLER_70_1337 ();
 FILLER_ASAP7_75t_R FILLER_70_1347 ();
 FILLER_ASAP7_75t_R FILLER_70_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_71_2 ();
 DECAPx6_ASAP7_75t_R FILLER_71_24 ();
 DECAPx2_ASAP7_75t_R FILLER_71_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_44 ();
 DECAPx6_ASAP7_75t_R FILLER_71_51 ();
 DECAPx1_ASAP7_75t_R FILLER_71_65 ();
 DECAPx10_ASAP7_75t_R FILLER_71_75 ();
 DECAPx2_ASAP7_75t_R FILLER_71_97 ();
 FILLER_ASAP7_75t_R FILLER_71_103 ();
 DECAPx2_ASAP7_75t_R FILLER_71_111 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_117 ();
 FILLER_ASAP7_75t_R FILLER_71_128 ();
 FILLER_ASAP7_75t_R FILLER_71_138 ();
 DECAPx2_ASAP7_75t_R FILLER_71_146 ();
 FILLER_ASAP7_75t_R FILLER_71_152 ();
 FILLER_ASAP7_75t_R FILLER_71_160 ();
 DECAPx1_ASAP7_75t_R FILLER_71_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_169 ();
 DECAPx4_ASAP7_75t_R FILLER_71_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_206 ();
 FILLER_ASAP7_75t_R FILLER_71_233 ();
 DECAPx10_ASAP7_75t_R FILLER_71_241 ();
 DECAPx1_ASAP7_75t_R FILLER_71_263 ();
 DECAPx10_ASAP7_75t_R FILLER_71_277 ();
 DECAPx6_ASAP7_75t_R FILLER_71_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_313 ();
 DECAPx4_ASAP7_75t_R FILLER_71_321 ();
 DECAPx6_ASAP7_75t_R FILLER_71_337 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_351 ();
 DECAPx1_ASAP7_75t_R FILLER_71_357 ();
 DECAPx6_ASAP7_75t_R FILLER_71_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_381 ();
 DECAPx10_ASAP7_75t_R FILLER_71_390 ();
 DECAPx6_ASAP7_75t_R FILLER_71_412 ();
 DECAPx1_ASAP7_75t_R FILLER_71_426 ();
 DECAPx1_ASAP7_75t_R FILLER_71_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_440 ();
 FILLER_ASAP7_75t_R FILLER_71_447 ();
 FILLER_ASAP7_75t_R FILLER_71_457 ();
 DECAPx1_ASAP7_75t_R FILLER_71_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_469 ();
 DECAPx6_ASAP7_75t_R FILLER_71_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_492 ();
 FILLER_ASAP7_75t_R FILLER_71_499 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_504 ();
 DECAPx1_ASAP7_75t_R FILLER_71_513 ();
 FILLER_ASAP7_75t_R FILLER_71_539 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_551 ();
 DECAPx2_ASAP7_75t_R FILLER_71_566 ();
 FILLER_ASAP7_75t_R FILLER_71_586 ();
 FILLER_ASAP7_75t_R FILLER_71_594 ();
 DECAPx4_ASAP7_75t_R FILLER_71_600 ();
 FILLER_ASAP7_75t_R FILLER_71_610 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_632 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_655 ();
 FILLER_ASAP7_75t_R FILLER_71_664 ();
 DECAPx10_ASAP7_75t_R FILLER_71_673 ();
 DECAPx2_ASAP7_75t_R FILLER_71_695 ();
 DECAPx10_ASAP7_75t_R FILLER_71_707 ();
 DECAPx1_ASAP7_75t_R FILLER_71_735 ();
 DECAPx1_ASAP7_75t_R FILLER_71_745 ();
 DECAPx4_ASAP7_75t_R FILLER_71_764 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_774 ();
 DECAPx6_ASAP7_75t_R FILLER_71_783 ();
 DECAPx2_ASAP7_75t_R FILLER_71_800 ();
 FILLER_ASAP7_75t_R FILLER_71_806 ();
 DECAPx4_ASAP7_75t_R FILLER_71_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_844 ();
 DECAPx10_ASAP7_75t_R FILLER_71_855 ();
 DECAPx4_ASAP7_75t_R FILLER_71_877 ();
 FILLER_ASAP7_75t_R FILLER_71_893 ();
 DECAPx1_ASAP7_75t_R FILLER_71_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_905 ();
 DECAPx4_ASAP7_75t_R FILLER_71_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_922 ();
 DECAPx2_ASAP7_75t_R FILLER_71_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_933 ();
 DECAPx1_ASAP7_75t_R FILLER_71_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_941 ();
 DECAPx2_ASAP7_75t_R FILLER_71_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_954 ();
 FILLER_ASAP7_75t_R FILLER_71_958 ();
 DECAPx2_ASAP7_75t_R FILLER_71_986 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1000 ();
 DECAPx6_ASAP7_75t_R FILLER_71_1022 ();
 FILLER_ASAP7_75t_R FILLER_71_1036 ();
 DECAPx2_ASAP7_75t_R FILLER_71_1050 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_1056 ();
 FILLER_ASAP7_75t_R FILLER_71_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_71_1113 ();
 FILLER_ASAP7_75t_R FILLER_71_1135 ();
 FILLER_ASAP7_75t_R FILLER_71_1145 ();
 FILLER_ASAP7_75t_R FILLER_71_1150 ();
 FILLER_ASAP7_75t_R FILLER_71_1162 ();
 FILLER_ASAP7_75t_R FILLER_71_1172 ();
 DECAPx4_ASAP7_75t_R FILLER_71_1177 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_1187 ();
 FILLER_ASAP7_75t_R FILLER_71_1193 ();
 FILLER_ASAP7_75t_R FILLER_71_1198 ();
 FILLER_ASAP7_75t_R FILLER_71_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_71_1237 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_1243 ();
 FILLER_ASAP7_75t_R FILLER_71_1255 ();
 DECAPx2_ASAP7_75t_R FILLER_71_1263 ();
 DECAPx6_ASAP7_75t_R FILLER_71_1272 ();
 DECAPx1_ASAP7_75t_R FILLER_71_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1290 ();
 DECAPx1_ASAP7_75t_R FILLER_71_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1305 ();
 FILLER_ASAP7_75t_R FILLER_71_1316 ();
 DECAPx1_ASAP7_75t_R FILLER_71_1321 ();
 DECAPx6_ASAP7_75t_R FILLER_71_1328 ();
 DECAPx2_ASAP7_75t_R FILLER_71_1342 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_1348 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_1355 ();
 FILLER_ASAP7_75t_R FILLER_71_1361 ();
 FILLER_ASAP7_75t_R FILLER_71_1368 ();
 FILLER_ASAP7_75t_R FILLER_71_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_72_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_8 ();
 DECAPx1_ASAP7_75t_R FILLER_72_15 ();
 DECAPx4_ASAP7_75t_R FILLER_72_22 ();
 FILLER_ASAP7_75t_R FILLER_72_32 ();
 DECAPx10_ASAP7_75t_R FILLER_72_37 ();
 FILLER_ASAP7_75t_R FILLER_72_59 ();
 DECAPx4_ASAP7_75t_R FILLER_72_87 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_123 ();
 FILLER_ASAP7_75t_R FILLER_72_132 ();
 FILLER_ASAP7_75t_R FILLER_72_141 ();
 DECAPx1_ASAP7_75t_R FILLER_72_169 ();
 DECAPx1_ASAP7_75t_R FILLER_72_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_183 ();
 DECAPx4_ASAP7_75t_R FILLER_72_187 ();
 DECAPx2_ASAP7_75t_R FILLER_72_203 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_209 ();
 DECAPx1_ASAP7_75t_R FILLER_72_218 ();
 DECAPx6_ASAP7_75t_R FILLER_72_225 ();
 DECAPx2_ASAP7_75t_R FILLER_72_239 ();
 DECAPx10_ASAP7_75t_R FILLER_72_253 ();
 FILLER_ASAP7_75t_R FILLER_72_281 ();
 DECAPx2_ASAP7_75t_R FILLER_72_286 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_295 ();
 DECAPx10_ASAP7_75t_R FILLER_72_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_328 ();
 DECAPx6_ASAP7_75t_R FILLER_72_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_369 ();
 DECAPx10_ASAP7_75t_R FILLER_72_376 ();
 DECAPx2_ASAP7_75t_R FILLER_72_404 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_410 ();
 FILLER_ASAP7_75t_R FILLER_72_419 ();
 DECAPx10_ASAP7_75t_R FILLER_72_427 ();
 DECAPx4_ASAP7_75t_R FILLER_72_449 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_459 ();
 DECAPx2_ASAP7_75t_R FILLER_72_464 ();
 FILLER_ASAP7_75t_R FILLER_72_470 ();
 FILLER_ASAP7_75t_R FILLER_72_478 ();
 DECAPx1_ASAP7_75t_R FILLER_72_483 ();
 FILLER_ASAP7_75t_R FILLER_72_513 ();
 DECAPx2_ASAP7_75t_R FILLER_72_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_529 ();
 DECAPx2_ASAP7_75t_R FILLER_72_536 ();
 FILLER_ASAP7_75t_R FILLER_72_542 ();
 FILLER_ASAP7_75t_R FILLER_72_556 ();
 DECAPx1_ASAP7_75t_R FILLER_72_570 ();
 FILLER_ASAP7_75t_R FILLER_72_588 ();
 DECAPx4_ASAP7_75t_R FILLER_72_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_606 ();
 FILLER_ASAP7_75t_R FILLER_72_617 ();
 DECAPx4_ASAP7_75t_R FILLER_72_623 ();
 FILLER_ASAP7_75t_R FILLER_72_633 ();
 DECAPx6_ASAP7_75t_R FILLER_72_641 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_675 ();
 FILLER_ASAP7_75t_R FILLER_72_685 ();
 DECAPx2_ASAP7_75t_R FILLER_72_693 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_705 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_715 ();
 DECAPx1_ASAP7_75t_R FILLER_72_740 ();
 FILLER_ASAP7_75t_R FILLER_72_754 ();
 DECAPx4_ASAP7_75t_R FILLER_72_762 ();
 FILLER_ASAP7_75t_R FILLER_72_780 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_808 ();
 FILLER_ASAP7_75t_R FILLER_72_818 ();
 FILLER_ASAP7_75t_R FILLER_72_826 ();
 DECAPx10_ASAP7_75t_R FILLER_72_831 ();
 DECAPx6_ASAP7_75t_R FILLER_72_853 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_867 ();
 FILLER_ASAP7_75t_R FILLER_72_877 ();
 DECAPx4_ASAP7_75t_R FILLER_72_885 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_895 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_910 ();
 FILLER_ASAP7_75t_R FILLER_72_921 ();
 FILLER_ASAP7_75t_R FILLER_72_931 ();
 FILLER_ASAP7_75t_R FILLER_72_941 ();
 DECAPx2_ASAP7_75t_R FILLER_72_951 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_957 ();
 FILLER_ASAP7_75t_R FILLER_72_963 ();
 DECAPx2_ASAP7_75t_R FILLER_72_972 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_988 ();
 FILLER_ASAP7_75t_R FILLER_72_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_72_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_72_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_72_1076 ();
 FILLER_ASAP7_75t_R FILLER_72_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_72_1090 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_1096 ();
 FILLER_ASAP7_75t_R FILLER_72_1102 ();
 DECAPx4_ASAP7_75t_R FILLER_72_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1120 ();
 FILLER_ASAP7_75t_R FILLER_72_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1137 ();
 DECAPx6_ASAP7_75t_R FILLER_72_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1210 ();
 DECAPx4_ASAP7_75t_R FILLER_72_1214 ();
 FILLER_ASAP7_75t_R FILLER_72_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1251 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_1255 ();
 DECAPx2_ASAP7_75t_R FILLER_72_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_72_1278 ();
 DECAPx4_ASAP7_75t_R FILLER_72_1300 ();
 FILLER_ASAP7_75t_R FILLER_72_1336 ();
 DECAPx6_ASAP7_75t_R FILLER_72_1341 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1355 ();
 DECAPx2_ASAP7_75t_R FILLER_72_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_1369 ();
 FILLER_ASAP7_75t_R FILLER_72_1375 ();
 FILLER_ASAP7_75t_R FILLER_73_2 ();
 DECAPx2_ASAP7_75t_R FILLER_73_30 ();
 FILLER_ASAP7_75t_R FILLER_73_42 ();
 FILLER_ASAP7_75t_R FILLER_73_52 ();
 DECAPx1_ASAP7_75t_R FILLER_73_60 ();
 DECAPx2_ASAP7_75t_R FILLER_73_70 ();
 DECAPx4_ASAP7_75t_R FILLER_73_79 ();
 FILLER_ASAP7_75t_R FILLER_73_99 ();
 DECAPx1_ASAP7_75t_R FILLER_73_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_111 ();
 DECAPx10_ASAP7_75t_R FILLER_73_115 ();
 DECAPx4_ASAP7_75t_R FILLER_73_137 ();
 FILLER_ASAP7_75t_R FILLER_73_147 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_155 ();
 DECAPx10_ASAP7_75t_R FILLER_73_161 ();
 DECAPx1_ASAP7_75t_R FILLER_73_183 ();
 DECAPx1_ASAP7_75t_R FILLER_73_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_217 ();
 DECAPx4_ASAP7_75t_R FILLER_73_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_234 ();
 DECAPx2_ASAP7_75t_R FILLER_73_238 ();
 FILLER_ASAP7_75t_R FILLER_73_244 ();
 DECAPx4_ASAP7_75t_R FILLER_73_254 ();
 FILLER_ASAP7_75t_R FILLER_73_264 ();
 DECAPx2_ASAP7_75t_R FILLER_73_292 ();
 DECAPx1_ASAP7_75t_R FILLER_73_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_310 ();
 DECAPx1_ASAP7_75t_R FILLER_73_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_322 ();
 FILLER_ASAP7_75t_R FILLER_73_329 ();
 DECAPx1_ASAP7_75t_R FILLER_73_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_341 ();
 FILLER_ASAP7_75t_R FILLER_73_364 ();
 DECAPx2_ASAP7_75t_R FILLER_73_392 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_398 ();
 DECAPx4_ASAP7_75t_R FILLER_73_409 ();
 FILLER_ASAP7_75t_R FILLER_73_419 ();
 DECAPx2_ASAP7_75t_R FILLER_73_429 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_435 ();
 DECAPx6_ASAP7_75t_R FILLER_73_444 ();
 DECAPx1_ASAP7_75t_R FILLER_73_458 ();
 FILLER_ASAP7_75t_R FILLER_73_488 ();
 DECAPx2_ASAP7_75t_R FILLER_73_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_502 ();
 FILLER_ASAP7_75t_R FILLER_73_509 ();
 FILLER_ASAP7_75t_R FILLER_73_517 ();
 DECAPx1_ASAP7_75t_R FILLER_73_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_529 ();
 FILLER_ASAP7_75t_R FILLER_73_542 ();
 FILLER_ASAP7_75t_R FILLER_73_556 ();
 FILLER_ASAP7_75t_R FILLER_73_572 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_588 ();
 FILLER_ASAP7_75t_R FILLER_73_605 ();
 DECAPx2_ASAP7_75t_R FILLER_73_619 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_625 ();
 DECAPx6_ASAP7_75t_R FILLER_73_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_646 ();
 FILLER_ASAP7_75t_R FILLER_73_653 ();
 DECAPx2_ASAP7_75t_R FILLER_73_662 ();
 DECAPx1_ASAP7_75t_R FILLER_73_674 ();
 DECAPx2_ASAP7_75t_R FILLER_73_698 ();
 FILLER_ASAP7_75t_R FILLER_73_704 ();
 DECAPx1_ASAP7_75t_R FILLER_73_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_730 ();
 DECAPx10_ASAP7_75t_R FILLER_73_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_759 ();
 DECAPx2_ASAP7_75t_R FILLER_73_766 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_772 ();
 FILLER_ASAP7_75t_R FILLER_73_781 ();
 DECAPx4_ASAP7_75t_R FILLER_73_789 ();
 FILLER_ASAP7_75t_R FILLER_73_799 ();
 DECAPx6_ASAP7_75t_R FILLER_73_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_821 ();
 DECAPx1_ASAP7_75t_R FILLER_73_825 ();
 DECAPx1_ASAP7_75t_R FILLER_73_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_841 ();
 DECAPx2_ASAP7_75t_R FILLER_73_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_854 ();
 DECAPx1_ASAP7_75t_R FILLER_73_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_865 ();
 FILLER_ASAP7_75t_R FILLER_73_869 ();
 DECAPx1_ASAP7_75t_R FILLER_73_891 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_907 ();
 DECAPx4_ASAP7_75t_R FILLER_73_913 ();
 FILLER_ASAP7_75t_R FILLER_73_923 ();
 DECAPx4_ASAP7_75t_R FILLER_73_927 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_937 ();
 DECAPx10_ASAP7_75t_R FILLER_73_946 ();
 DECAPx4_ASAP7_75t_R FILLER_73_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_978 ();
 DECAPx10_ASAP7_75t_R FILLER_73_987 ();
 DECAPx1_ASAP7_75t_R FILLER_73_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1013 ();
 FILLER_ASAP7_75t_R FILLER_73_1022 ();
 DECAPx6_ASAP7_75t_R FILLER_73_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1041 ();
 FILLER_ASAP7_75t_R FILLER_73_1068 ();
 DECAPx4_ASAP7_75t_R FILLER_73_1073 ();
 DECAPx1_ASAP7_75t_R FILLER_73_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1099 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1108 ();
 FILLER_ASAP7_75t_R FILLER_73_1114 ();
 FILLER_ASAP7_75t_R FILLER_73_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1150 ();
 DECAPx4_ASAP7_75t_R FILLER_73_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1182 ();
 FILLER_ASAP7_75t_R FILLER_73_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1238 ();
 DECAPx1_ASAP7_75t_R FILLER_73_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_73_1294 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1316 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_1322 ();
 FILLER_ASAP7_75t_R FILLER_73_1332 ();
 DECAPx2_ASAP7_75t_R FILLER_73_1341 ();
 FILLER_ASAP7_75t_R FILLER_73_1347 ();
 FILLER_ASAP7_75t_R FILLER_73_1375 ();
 FILLER_ASAP7_75t_R FILLER_74_2 ();
 FILLER_ASAP7_75t_R FILLER_74_10 ();
 DECAPx1_ASAP7_75t_R FILLER_74_38 ();
 DECAPx4_ASAP7_75t_R FILLER_74_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_60 ();
 DECAPx1_ASAP7_75t_R FILLER_74_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_71 ();
 DECAPx2_ASAP7_75t_R FILLER_74_78 ();
 FILLER_ASAP7_75t_R FILLER_74_90 ();
 DECAPx10_ASAP7_75t_R FILLER_74_95 ();
 DECAPx6_ASAP7_75t_R FILLER_74_117 ();
 DECAPx10_ASAP7_75t_R FILLER_74_137 ();
 FILLER_ASAP7_75t_R FILLER_74_159 ();
 DECAPx2_ASAP7_75t_R FILLER_74_167 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_74_173 ();
 DECAPx4_ASAP7_75t_R FILLER_74_182 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_74_198 ();
 DECAPx1_ASAP7_75t_R FILLER_74_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_208 ();
 DECAPx1_ASAP7_75t_R FILLER_74_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_239 ();
 FILLER_ASAP7_75t_R FILLER_74_246 ();
 FILLER_ASAP7_75t_R FILLER_74_254 ();
 DECAPx2_ASAP7_75t_R FILLER_74_262 ();
 FILLER_ASAP7_75t_R FILLER_74_268 ();
 FILLER_ASAP7_75t_R FILLER_74_276 ();
 DECAPx4_ASAP7_75t_R FILLER_74_284 ();
 FILLER_ASAP7_75t_R FILLER_74_300 ();
 DECAPx4_ASAP7_75t_R FILLER_74_308 ();
 FILLER_ASAP7_75t_R FILLER_74_318 ();
 FILLER_ASAP7_75t_R FILLER_74_326 ();
 DECAPx2_ASAP7_75t_R FILLER_74_334 ();
 FILLER_ASAP7_75t_R FILLER_74_340 ();
 FILLER_ASAP7_75t_R FILLER_74_345 ();
 DECAPx4_ASAP7_75t_R FILLER_74_357 ();
 DECAPx2_ASAP7_75t_R FILLER_74_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_379 ();
 DECAPx6_ASAP7_75t_R FILLER_74_383 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_74_397 ();
 DECAPx2_ASAP7_75t_R FILLER_74_408 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_74_414 ();
 DECAPx2_ASAP7_75t_R FILLER_74_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_434 ();
 DECAPx2_ASAP7_75t_R FILLER_74_443 ();
 FILLER_ASAP7_75t_R FILLER_74_449 ();
 DECAPx1_ASAP7_75t_R FILLER_74_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_461 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_74_464 ();
 DECAPx1_ASAP7_75t_R FILLER_74_473 ();
 DECAPx10_ASAP7_75t_R FILLER_74_480 ();
 DECAPx2_ASAP7_75t_R FILLER_74_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_508 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_74_517 ();
 FILLER_ASAP7_75t_R FILLER_74_526 ();
 FILLER_ASAP7_75t_R FILLER_74_550 ();
 DECAPx2_ASAP7_75t_R FILLER_74_564 ();
 FILLER_ASAP7_75t_R FILLER_74_570 ();
 DECAPx2_ASAP7_75t_R FILLER_74_586 ();
 FILLER_ASAP7_75t_R FILLER_74_606 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_74_618 ();
 FILLER_ASAP7_75t_R FILLER_74_633 ();
 DECAPx6_ASAP7_75t_R FILLER_74_642 ();
 DECAPx10_ASAP7_75t_R FILLER_74_663 ();
 DECAPx10_ASAP7_75t_R FILLER_74_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_714 ();
 DECAPx2_ASAP7_75t_R FILLER_74_721 ();
 DECAPx10_ASAP7_75t_R FILLER_74_734 ();
 DECAPx1_ASAP7_75t_R FILLER_74_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_760 ();
 DECAPx2_ASAP7_75t_R FILLER_74_781 ();
 FILLER_ASAP7_75t_R FILLER_74_787 ();
 FILLER_ASAP7_75t_R FILLER_74_792 ();
 DECAPx6_ASAP7_75t_R FILLER_74_805 ();
 DECAPx1_ASAP7_75t_R FILLER_74_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_823 ();
 DECAPx2_ASAP7_75t_R FILLER_74_830 ();
 FILLER_ASAP7_75t_R FILLER_74_844 ();
 FILLER_ASAP7_75t_R FILLER_74_852 ();
 DECAPx2_ASAP7_75t_R FILLER_74_860 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_74_866 ();
 DECAPx10_ASAP7_75t_R FILLER_74_878 ();
 DECAPx2_ASAP7_75t_R FILLER_74_900 ();
 DECAPx6_ASAP7_75t_R FILLER_74_909 ();
 DECAPx2_ASAP7_75t_R FILLER_74_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_929 ();
 FILLER_ASAP7_75t_R FILLER_74_933 ();
 DECAPx1_ASAP7_75t_R FILLER_74_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_965 ();
 DECAPx2_ASAP7_75t_R FILLER_74_972 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_74_988 ();
 DECAPx4_ASAP7_75t_R FILLER_74_994 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_74_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1015 ();
 FILLER_ASAP7_75t_R FILLER_74_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1033 ();
 FILLER_ASAP7_75t_R FILLER_74_1049 ();
 FILLER_ASAP7_75t_R FILLER_74_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1080 ();
 FILLER_ASAP7_75t_R FILLER_74_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1122 ();
 DECAPx4_ASAP7_75t_R FILLER_74_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1149 ();
 FILLER_ASAP7_75t_R FILLER_74_1156 ();
 FILLER_ASAP7_75t_R FILLER_74_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1174 ();
 FILLER_ASAP7_75t_R FILLER_74_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1214 ();
 FILLER_ASAP7_75t_R FILLER_74_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1259 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_74_1266 ();
 FILLER_ASAP7_75t_R FILLER_74_1275 ();
 DECAPx4_ASAP7_75t_R FILLER_74_1303 ();
 FILLER_ASAP7_75t_R FILLER_74_1313 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1322 ();
 FILLER_ASAP7_75t_R FILLER_74_1328 ();
 DECAPx1_ASAP7_75t_R FILLER_74_1333 ();
 DECAPx4_ASAP7_75t_R FILLER_74_1347 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_1357 ();
 FILLER_ASAP7_75t_R FILLER_74_1364 ();
 DECAPx2_ASAP7_75t_R FILLER_74_1369 ();
 FILLER_ASAP7_75t_R FILLER_74_1375 ();
 DECAPx4_ASAP7_75t_R FILLER_75_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_12 ();
 FILLER_ASAP7_75t_R FILLER_75_21 ();
 FILLER_ASAP7_75t_R FILLER_75_29 ();
 DECAPx1_ASAP7_75t_R FILLER_75_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_38 ();
 DECAPx10_ASAP7_75t_R FILLER_75_45 ();
 DECAPx4_ASAP7_75t_R FILLER_75_67 ();
 DECAPx1_ASAP7_75t_R FILLER_75_103 ();
 DECAPx1_ASAP7_75t_R FILLER_75_113 ();
 DECAPx6_ASAP7_75t_R FILLER_75_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_137 ();
 FILLER_ASAP7_75t_R FILLER_75_144 ();
 DECAPx2_ASAP7_75t_R FILLER_75_152 ();
 DECAPx2_ASAP7_75t_R FILLER_75_166 ();
 DECAPx6_ASAP7_75t_R FILLER_75_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_212 ();
 DECAPx1_ASAP7_75t_R FILLER_75_219 ();
 DECAPx2_ASAP7_75t_R FILLER_75_226 ();
 DECAPx2_ASAP7_75t_R FILLER_75_258 ();
 FILLER_ASAP7_75t_R FILLER_75_264 ();
 DECAPx10_ASAP7_75t_R FILLER_75_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_314 ();
 DECAPx2_ASAP7_75t_R FILLER_75_323 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_329 ();
 FILLER_ASAP7_75t_R FILLER_75_338 ();
 FILLER_ASAP7_75t_R FILLER_75_346 ();
 DECAPx6_ASAP7_75t_R FILLER_75_356 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_370 ();
 FILLER_ASAP7_75t_R FILLER_75_379 ();
 DECAPx2_ASAP7_75t_R FILLER_75_384 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_390 ();
 FILLER_ASAP7_75t_R FILLER_75_396 ();
 DECAPx2_ASAP7_75t_R FILLER_75_404 ();
 DECAPx2_ASAP7_75t_R FILLER_75_417 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_423 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_432 ();
 DECAPx1_ASAP7_75t_R FILLER_75_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_447 ();
 DECAPx4_ASAP7_75t_R FILLER_75_474 ();
 FILLER_ASAP7_75t_R FILLER_75_484 ();
 DECAPx2_ASAP7_75t_R FILLER_75_489 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_495 ();
 DECAPx4_ASAP7_75t_R FILLER_75_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_511 ();
 DECAPx2_ASAP7_75t_R FILLER_75_520 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_526 ();
 FILLER_ASAP7_75t_R FILLER_75_551 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_565 ();
 DECAPx2_ASAP7_75t_R FILLER_75_582 ();
 FILLER_ASAP7_75t_R FILLER_75_602 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_611 ();
 DECAPx2_ASAP7_75t_R FILLER_75_621 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_627 ();
 FILLER_ASAP7_75t_R FILLER_75_650 ();
 DECAPx6_ASAP7_75t_R FILLER_75_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_686 ();
 DECAPx4_ASAP7_75t_R FILLER_75_707 ();
 FILLER_ASAP7_75t_R FILLER_75_717 ();
 DECAPx1_ASAP7_75t_R FILLER_75_725 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_749 ();
 DECAPx1_ASAP7_75t_R FILLER_75_758 ();
 DECAPx6_ASAP7_75t_R FILLER_75_768 ();
 DECAPx2_ASAP7_75t_R FILLER_75_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_788 ();
 DECAPx6_ASAP7_75t_R FILLER_75_793 ();
 FILLER_ASAP7_75t_R FILLER_75_814 ();
 DECAPx2_ASAP7_75t_R FILLER_75_822 ();
 FILLER_ASAP7_75t_R FILLER_75_828 ();
 FILLER_ASAP7_75t_R FILLER_75_840 ();
 FILLER_ASAP7_75t_R FILLER_75_850 ();
 DECAPx2_ASAP7_75t_R FILLER_75_858 ();
 DECAPx10_ASAP7_75t_R FILLER_75_867 ();
 DECAPx4_ASAP7_75t_R FILLER_75_889 ();
 FILLER_ASAP7_75t_R FILLER_75_899 ();
 DECAPx6_ASAP7_75t_R FILLER_75_909 ();
 FILLER_ASAP7_75t_R FILLER_75_923 ();
 FILLER_ASAP7_75t_R FILLER_75_927 ();
 DECAPx2_ASAP7_75t_R FILLER_75_941 ();
 FILLER_ASAP7_75t_R FILLER_75_947 ();
 FILLER_ASAP7_75t_R FILLER_75_952 ();
 DECAPx2_ASAP7_75t_R FILLER_75_966 ();
 DECAPx4_ASAP7_75t_R FILLER_75_979 ();
 FILLER_ASAP7_75t_R FILLER_75_989 ();
 DECAPx1_ASAP7_75t_R FILLER_75_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_75_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1054 ();
 FILLER_ASAP7_75t_R FILLER_75_1060 ();
 FILLER_ASAP7_75t_R FILLER_75_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_75_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_75_1097 ();
 DECAPx1_ASAP7_75t_R FILLER_75_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_75_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1144 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_1151 ();
 FILLER_ASAP7_75t_R FILLER_75_1164 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_1192 ();
 FILLER_ASAP7_75t_R FILLER_75_1198 ();
 FILLER_ASAP7_75t_R FILLER_75_1226 ();
 FILLER_ASAP7_75t_R FILLER_75_1235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_1249 ();
 DECAPx6_ASAP7_75t_R FILLER_75_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1276 ();
 DECAPx4_ASAP7_75t_R FILLER_75_1284 ();
 DECAPx2_ASAP7_75t_R FILLER_75_1301 ();
 DECAPx1_ASAP7_75t_R FILLER_75_1310 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_1314 ();
 FILLER_ASAP7_75t_R FILLER_75_1341 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_1350 ();
 FILLER_ASAP7_75t_R FILLER_75_1360 ();
 FILLER_ASAP7_75t_R FILLER_75_1368 ();
 FILLER_ASAP7_75t_R FILLER_75_1375 ();
 FILLER_ASAP7_75t_R FILLER_76_2 ();
 DECAPx2_ASAP7_75t_R FILLER_76_30 ();
 FILLER_ASAP7_75t_R FILLER_76_36 ();
 DECAPx2_ASAP7_75t_R FILLER_76_44 ();
 FILLER_ASAP7_75t_R FILLER_76_50 ();
 FILLER_ASAP7_75t_R FILLER_76_55 ();
 DECAPx6_ASAP7_75t_R FILLER_76_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_79 ();
 DECAPx6_ASAP7_75t_R FILLER_76_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_100 ();
 DECAPx2_ASAP7_75t_R FILLER_76_127 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_136 ();
 DECAPx4_ASAP7_75t_R FILLER_76_147 ();
 FILLER_ASAP7_75t_R FILLER_76_157 ();
 DECAPx2_ASAP7_75t_R FILLER_76_167 ();
 FILLER_ASAP7_75t_R FILLER_76_173 ();
 DECAPx1_ASAP7_75t_R FILLER_76_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_185 ();
 DECAPx10_ASAP7_75t_R FILLER_76_189 ();
 DECAPx10_ASAP7_75t_R FILLER_76_211 ();
 FILLER_ASAP7_75t_R FILLER_76_233 ();
 DECAPx1_ASAP7_75t_R FILLER_76_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_245 ();
 DECAPx6_ASAP7_75t_R FILLER_76_249 ();
 DECAPx1_ASAP7_75t_R FILLER_76_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_267 ();
 DECAPx2_ASAP7_75t_R FILLER_76_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_280 ();
 DECAPx1_ASAP7_75t_R FILLER_76_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_288 ();
 DECAPx2_ASAP7_75t_R FILLER_76_295 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_301 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_307 ();
 DECAPx4_ASAP7_75t_R FILLER_76_317 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_327 ();
 DECAPx4_ASAP7_75t_R FILLER_76_356 ();
 FILLER_ASAP7_75t_R FILLER_76_392 ();
 DECAPx1_ASAP7_75t_R FILLER_76_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_409 ();
 DECAPx1_ASAP7_75t_R FILLER_76_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_422 ();
 DECAPx4_ASAP7_75t_R FILLER_76_429 ();
 DECAPx2_ASAP7_75t_R FILLER_76_445 ();
 DECAPx1_ASAP7_75t_R FILLER_76_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_461 ();
 FILLER_ASAP7_75t_R FILLER_76_464 ();
 FILLER_ASAP7_75t_R FILLER_76_469 ();
 FILLER_ASAP7_75t_R FILLER_76_497 ();
 FILLER_ASAP7_75t_R FILLER_76_505 ();
 FILLER_ASAP7_75t_R FILLER_76_513 ();
 FILLER_ASAP7_75t_R FILLER_76_533 ();
 DECAPx1_ASAP7_75t_R FILLER_76_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_547 ();
 DECAPx2_ASAP7_75t_R FILLER_76_560 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_566 ();
 DECAPx2_ASAP7_75t_R FILLER_76_583 ();
 FILLER_ASAP7_75t_R FILLER_76_597 ();
 DECAPx2_ASAP7_75t_R FILLER_76_607 ();
 DECAPx1_ASAP7_75t_R FILLER_76_627 ();
 FILLER_ASAP7_75t_R FILLER_76_657 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_666 ();
 DECAPx1_ASAP7_75t_R FILLER_76_689 ();
 FILLER_ASAP7_75t_R FILLER_76_700 ();
 DECAPx2_ASAP7_75t_R FILLER_76_709 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_715 ();
 FILLER_ASAP7_75t_R FILLER_76_724 ();
 DECAPx6_ASAP7_75t_R FILLER_76_732 ();
 DECAPx1_ASAP7_75t_R FILLER_76_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_750 ();
 FILLER_ASAP7_75t_R FILLER_76_759 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_768 ();
 DECAPx10_ASAP7_75t_R FILLER_76_776 ();
 DECAPx1_ASAP7_75t_R FILLER_76_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_802 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_806 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_815 ();
 DECAPx6_ASAP7_75t_R FILLER_76_828 ();
 DECAPx2_ASAP7_75t_R FILLER_76_842 ();
 DECAPx1_ASAP7_75t_R FILLER_76_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_860 ();
 DECAPx1_ASAP7_75t_R FILLER_76_870 ();
 FILLER_ASAP7_75t_R FILLER_76_880 ();
 FILLER_ASAP7_75t_R FILLER_76_888 ();
 DECAPx1_ASAP7_75t_R FILLER_76_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_900 ();
 DECAPx2_ASAP7_75t_R FILLER_76_910 ();
 DECAPx2_ASAP7_75t_R FILLER_76_928 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_934 ();
 FILLER_ASAP7_75t_R FILLER_76_963 ();
 FILLER_ASAP7_75t_R FILLER_76_968 ();
 DECAPx6_ASAP7_75t_R FILLER_76_973 ();
 DECAPx2_ASAP7_75t_R FILLER_76_987 ();
 FILLER_ASAP7_75t_R FILLER_76_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1009 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_1015 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1021 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_1035 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1044 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1065 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1091 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1102 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_1111 ();
 FILLER_ASAP7_75t_R FILLER_76_1117 ();
 FILLER_ASAP7_75t_R FILLER_76_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1155 ();
 DECAPx4_ASAP7_75t_R FILLER_76_1168 ();
 FILLER_ASAP7_75t_R FILLER_76_1178 ();
 DECAPx6_ASAP7_75t_R FILLER_76_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1203 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_1212 ();
 DECAPx4_ASAP7_75t_R FILLER_76_1218 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_1228 ();
 FILLER_ASAP7_75t_R FILLER_76_1237 ();
 DECAPx4_ASAP7_75t_R FILLER_76_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1252 ();
 DECAPx1_ASAP7_75t_R FILLER_76_1261 ();
 DECAPx2_ASAP7_75t_R FILLER_76_1271 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_1277 ();
 FILLER_ASAP7_75t_R FILLER_76_1290 ();
 FILLER_ASAP7_75t_R FILLER_76_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_76_1326 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_1348 ();
 FILLER_ASAP7_75t_R FILLER_76_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_77_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_8 ();
 DECAPx4_ASAP7_75t_R FILLER_77_17 ();
 FILLER_ASAP7_75t_R FILLER_77_27 ();
 DECAPx1_ASAP7_75t_R FILLER_77_55 ();
 FILLER_ASAP7_75t_R FILLER_77_65 ();
 DECAPx1_ASAP7_75t_R FILLER_77_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_77 ();
 FILLER_ASAP7_75t_R FILLER_77_88 ();
 DECAPx2_ASAP7_75t_R FILLER_77_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_102 ();
 DECAPx2_ASAP7_75t_R FILLER_77_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_115 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_119 ();
 FILLER_ASAP7_75t_R FILLER_77_128 ();
 DECAPx2_ASAP7_75t_R FILLER_77_133 ();
 FILLER_ASAP7_75t_R FILLER_77_145 ();
 DECAPx2_ASAP7_75t_R FILLER_77_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_161 ();
 DECAPx10_ASAP7_75t_R FILLER_77_168 ();
 DECAPx6_ASAP7_75t_R FILLER_77_190 ();
 FILLER_ASAP7_75t_R FILLER_77_210 ();
 DECAPx6_ASAP7_75t_R FILLER_77_215 ();
 FILLER_ASAP7_75t_R FILLER_77_229 ();
 DECAPx10_ASAP7_75t_R FILLER_77_237 ();
 DECAPx6_ASAP7_75t_R FILLER_77_259 ();
 DECAPx1_ASAP7_75t_R FILLER_77_273 ();
 DECAPx2_ASAP7_75t_R FILLER_77_303 ();
 DECAPx2_ASAP7_75t_R FILLER_77_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_321 ();
 FILLER_ASAP7_75t_R FILLER_77_330 ();
 DECAPx2_ASAP7_75t_R FILLER_77_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_344 ();
 DECAPx6_ASAP7_75t_R FILLER_77_348 ();
 FILLER_ASAP7_75t_R FILLER_77_368 ();
 DECAPx10_ASAP7_75t_R FILLER_77_376 ();
 DECAPx1_ASAP7_75t_R FILLER_77_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_402 ();
 FILLER_ASAP7_75t_R FILLER_77_425 ();
 DECAPx10_ASAP7_75t_R FILLER_77_435 ();
 DECAPx4_ASAP7_75t_R FILLER_77_457 ();
 FILLER_ASAP7_75t_R FILLER_77_467 ();
 FILLER_ASAP7_75t_R FILLER_77_475 ();
 FILLER_ASAP7_75t_R FILLER_77_483 ();
 FILLER_ASAP7_75t_R FILLER_77_511 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_521 ();
 FILLER_ASAP7_75t_R FILLER_77_530 ();
 FILLER_ASAP7_75t_R FILLER_77_550 ();
 DECAPx1_ASAP7_75t_R FILLER_77_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_568 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_587 ();
 FILLER_ASAP7_75t_R FILLER_77_598 ();
 FILLER_ASAP7_75t_R FILLER_77_608 ();
 FILLER_ASAP7_75t_R FILLER_77_622 ();
 DECAPx1_ASAP7_75t_R FILLER_77_629 ();
 DECAPx2_ASAP7_75t_R FILLER_77_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_644 ();
 DECAPx10_ASAP7_75t_R FILLER_77_648 ();
 FILLER_ASAP7_75t_R FILLER_77_677 ();
 DECAPx6_ASAP7_75t_R FILLER_77_683 ();
 DECAPx1_ASAP7_75t_R FILLER_77_697 ();
 FILLER_ASAP7_75t_R FILLER_77_721 ();
 DECAPx1_ASAP7_75t_R FILLER_77_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_733 ();
 FILLER_ASAP7_75t_R FILLER_77_742 ();
 DECAPx6_ASAP7_75t_R FILLER_77_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_766 ();
 FILLER_ASAP7_75t_R FILLER_77_770 ();
 FILLER_ASAP7_75t_R FILLER_77_778 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_788 ();
 DECAPx10_ASAP7_75t_R FILLER_77_811 ();
 DECAPx10_ASAP7_75t_R FILLER_77_833 ();
 DECAPx1_ASAP7_75t_R FILLER_77_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_859 ();
 FILLER_ASAP7_75t_R FILLER_77_866 ();
 FILLER_ASAP7_75t_R FILLER_77_876 ();
 FILLER_ASAP7_75t_R FILLER_77_884 ();
 FILLER_ASAP7_75t_R FILLER_77_892 ();
 FILLER_ASAP7_75t_R FILLER_77_897 ();
 FILLER_ASAP7_75t_R FILLER_77_905 ();
 DECAPx4_ASAP7_75t_R FILLER_77_913 ();
 FILLER_ASAP7_75t_R FILLER_77_923 ();
 FILLER_ASAP7_75t_R FILLER_77_927 ();
 DECAPx4_ASAP7_75t_R FILLER_77_941 ();
 DECAPx10_ASAP7_75t_R FILLER_77_954 ();
 DECAPx1_ASAP7_75t_R FILLER_77_976 ();
 DECAPx4_ASAP7_75t_R FILLER_77_989 ();
 FILLER_ASAP7_75t_R FILLER_77_999 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1008 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_1030 ();
 FILLER_ASAP7_75t_R FILLER_77_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1087 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1119 ();
 FILLER_ASAP7_75t_R FILLER_77_1125 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1133 ();
 FILLER_ASAP7_75t_R FILLER_77_1139 ();
 FILLER_ASAP7_75t_R FILLER_77_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1174 ();
 FILLER_ASAP7_75t_R FILLER_77_1180 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1202 ();
 DECAPx4_ASAP7_75t_R FILLER_77_1224 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_1234 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1249 ();
 DECAPx4_ASAP7_75t_R FILLER_77_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_1273 ();
 DECAPx6_ASAP7_75t_R FILLER_77_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_77_1302 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1324 ();
 FILLER_ASAP7_75t_R FILLER_77_1330 ();
 DECAPx4_ASAP7_75t_R FILLER_77_1340 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_1350 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1360 ();
 DECAPx2_ASAP7_75t_R FILLER_77_1369 ();
 FILLER_ASAP7_75t_R FILLER_77_1375 ();
 DECAPx1_ASAP7_75t_R FILLER_78_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_6 ();
 DECAPx1_ASAP7_75t_R FILLER_78_13 ();
 DECAPx4_ASAP7_75t_R FILLER_78_20 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_78_30 ();
 DECAPx1_ASAP7_75t_R FILLER_78_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_43 ();
 DECAPx2_ASAP7_75t_R FILLER_78_47 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_78_53 ();
 DECAPx10_ASAP7_75t_R FILLER_78_62 ();
 DECAPx2_ASAP7_75t_R FILLER_78_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_78_96 ();
 DECAPx4_ASAP7_75t_R FILLER_78_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_115 ();
 DECAPx6_ASAP7_75t_R FILLER_78_142 ();
 FILLER_ASAP7_75t_R FILLER_78_156 ();
 DECAPx6_ASAP7_75t_R FILLER_78_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_179 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_78_186 ();
 DECAPx1_ASAP7_75t_R FILLER_78_192 ();
 DECAPx2_ASAP7_75t_R FILLER_78_222 ();
 FILLER_ASAP7_75t_R FILLER_78_234 ();
 DECAPx2_ASAP7_75t_R FILLER_78_254 ();
 DECAPx1_ASAP7_75t_R FILLER_78_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_274 ();
 FILLER_ASAP7_75t_R FILLER_78_282 ();
 FILLER_ASAP7_75t_R FILLER_78_291 ();
 FILLER_ASAP7_75t_R FILLER_78_299 ();
 DECAPx2_ASAP7_75t_R FILLER_78_304 ();
 DECAPx1_ASAP7_75t_R FILLER_78_316 ();
 DECAPx4_ASAP7_75t_R FILLER_78_326 ();
 DECAPx1_ASAP7_75t_R FILLER_78_342 ();
 DECAPx1_ASAP7_75t_R FILLER_78_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_356 ();
 DECAPx6_ASAP7_75t_R FILLER_78_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_397 ();
 DECAPx2_ASAP7_75t_R FILLER_78_404 ();
 FILLER_ASAP7_75t_R FILLER_78_413 ();
 DECAPx6_ASAP7_75t_R FILLER_78_421 ();
 DECAPx1_ASAP7_75t_R FILLER_78_435 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_78_442 ();
 DECAPx4_ASAP7_75t_R FILLER_78_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_461 ();
 FILLER_ASAP7_75t_R FILLER_78_464 ();
 FILLER_ASAP7_75t_R FILLER_78_488 ();
 FILLER_ASAP7_75t_R FILLER_78_496 ();
 DECAPx2_ASAP7_75t_R FILLER_78_520 ();
 FILLER_ASAP7_75t_R FILLER_78_526 ();
 DECAPx2_ASAP7_75t_R FILLER_78_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_540 ();
 DECAPx2_ASAP7_75t_R FILLER_78_563 ();
 FILLER_ASAP7_75t_R FILLER_78_591 ();
 FILLER_ASAP7_75t_R FILLER_78_607 ();
 DECAPx4_ASAP7_75t_R FILLER_78_617 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_78_627 ();
 DECAPx6_ASAP7_75t_R FILLER_78_636 ();
 FILLER_ASAP7_75t_R FILLER_78_650 ();
 DECAPx10_ASAP7_75t_R FILLER_78_659 ();
 DECAPx6_ASAP7_75t_R FILLER_78_681 ();
 FILLER_ASAP7_75t_R FILLER_78_695 ();
 DECAPx10_ASAP7_75t_R FILLER_78_703 ();
 DECAPx10_ASAP7_75t_R FILLER_78_725 ();
 DECAPx2_ASAP7_75t_R FILLER_78_747 ();
 DECAPx2_ASAP7_75t_R FILLER_78_769 ();
 FILLER_ASAP7_75t_R FILLER_78_775 ();
 FILLER_ASAP7_75t_R FILLER_78_787 ();
 DECAPx2_ASAP7_75t_R FILLER_78_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_803 ();
 DECAPx6_ASAP7_75t_R FILLER_78_810 ();
 FILLER_ASAP7_75t_R FILLER_78_824 ();
 FILLER_ASAP7_75t_R FILLER_78_829 ();
 FILLER_ASAP7_75t_R FILLER_78_843 ();
 DECAPx4_ASAP7_75t_R FILLER_78_848 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_78_858 ();
 DECAPx10_ASAP7_75t_R FILLER_78_867 ();
 DECAPx4_ASAP7_75t_R FILLER_78_889 ();
 FILLER_ASAP7_75t_R FILLER_78_899 ();
 DECAPx4_ASAP7_75t_R FILLER_78_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_917 ();
 DECAPx6_ASAP7_75t_R FILLER_78_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_944 ();
 DECAPx4_ASAP7_75t_R FILLER_78_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_963 ();
 DECAPx1_ASAP7_75t_R FILLER_78_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_975 ();
 DECAPx2_ASAP7_75t_R FILLER_78_982 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_78_988 ();
 DECAPx6_ASAP7_75t_R FILLER_78_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1008 ();
 FILLER_ASAP7_75t_R FILLER_78_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_78_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1078 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_78_1084 ();
 FILLER_ASAP7_75t_R FILLER_78_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_78_1105 ();
 FILLER_ASAP7_75t_R FILLER_78_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_78_1124 ();
 FILLER_ASAP7_75t_R FILLER_78_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1167 ();
 DECAPx1_ASAP7_75t_R FILLER_78_1183 ();
 FILLER_ASAP7_75t_R FILLER_78_1199 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1217 ();
 DECAPx6_ASAP7_75t_R FILLER_78_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1258 ();
 FILLER_ASAP7_75t_R FILLER_78_1269 ();
 DECAPx6_ASAP7_75t_R FILLER_78_1297 ();
 FILLER_ASAP7_75t_R FILLER_78_1311 ();
 DECAPx2_ASAP7_75t_R FILLER_78_1320 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_1326 ();
 FILLER_ASAP7_75t_R FILLER_78_1333 ();
 DECAPx1_ASAP7_75t_R FILLER_78_1345 ();
 FILLER_ASAP7_75t_R FILLER_78_1375 ();
 DECAPx4_ASAP7_75t_R FILLER_79_2 ();
 FILLER_ASAP7_75t_R FILLER_79_12 ();
 FILLER_ASAP7_75t_R FILLER_79_20 ();
 DECAPx10_ASAP7_75t_R FILLER_79_28 ();
 DECAPx6_ASAP7_75t_R FILLER_79_50 ();
 DECAPx1_ASAP7_75t_R FILLER_79_64 ();
 FILLER_ASAP7_75t_R FILLER_79_74 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_79 ();
 FILLER_ASAP7_75t_R FILLER_79_92 ();
 FILLER_ASAP7_75t_R FILLER_79_97 ();
 DECAPx4_ASAP7_75t_R FILLER_79_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_117 ();
 DECAPx10_ASAP7_75t_R FILLER_79_124 ();
 DECAPx4_ASAP7_75t_R FILLER_79_146 ();
 FILLER_ASAP7_75t_R FILLER_79_156 ();
 DECAPx2_ASAP7_75t_R FILLER_79_165 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_171 ();
 FILLER_ASAP7_75t_R FILLER_79_200 ();
 FILLER_ASAP7_75t_R FILLER_79_208 ();
 FILLER_ASAP7_75t_R FILLER_79_236 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_244 ();
 FILLER_ASAP7_75t_R FILLER_79_273 ();
 FILLER_ASAP7_75t_R FILLER_79_282 ();
 FILLER_ASAP7_75t_R FILLER_79_291 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_296 ();
 DECAPx1_ASAP7_75t_R FILLER_79_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_329 ();
 DECAPx4_ASAP7_75t_R FILLER_79_356 ();
 FILLER_ASAP7_75t_R FILLER_79_366 ();
 FILLER_ASAP7_75t_R FILLER_79_374 ();
 DECAPx2_ASAP7_75t_R FILLER_79_379 ();
 FILLER_ASAP7_75t_R FILLER_79_385 ();
 DECAPx2_ASAP7_75t_R FILLER_79_413 ();
 FILLER_ASAP7_75t_R FILLER_79_425 ();
 DECAPx2_ASAP7_75t_R FILLER_79_430 ();
 FILLER_ASAP7_75t_R FILLER_79_442 ();
 FILLER_ASAP7_75t_R FILLER_79_470 ();
 FILLER_ASAP7_75t_R FILLER_79_478 ();
 DECAPx6_ASAP7_75t_R FILLER_79_483 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_497 ();
 DECAPx2_ASAP7_75t_R FILLER_79_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_509 ();
 DECAPx1_ASAP7_75t_R FILLER_79_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_520 ();
 FILLER_ASAP7_75t_R FILLER_79_547 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_561 ();
 FILLER_ASAP7_75t_R FILLER_79_578 ();
 FILLER_ASAP7_75t_R FILLER_79_602 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_610 ();
 DECAPx4_ASAP7_75t_R FILLER_79_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_631 ();
 FILLER_ASAP7_75t_R FILLER_79_658 ();
 DECAPx6_ASAP7_75t_R FILLER_79_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_694 ();
 FILLER_ASAP7_75t_R FILLER_79_701 ();
 DECAPx2_ASAP7_75t_R FILLER_79_709 ();
 FILLER_ASAP7_75t_R FILLER_79_715 ();
 DECAPx6_ASAP7_75t_R FILLER_79_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_737 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_745 ();
 FILLER_ASAP7_75t_R FILLER_79_754 ();
 DECAPx10_ASAP7_75t_R FILLER_79_762 ();
 DECAPx1_ASAP7_75t_R FILLER_79_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_788 ();
 DECAPx2_ASAP7_75t_R FILLER_79_795 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_801 ();
 FILLER_ASAP7_75t_R FILLER_79_810 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_824 ();
 DECAPx1_ASAP7_75t_R FILLER_79_839 ();
 DECAPx1_ASAP7_75t_R FILLER_79_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_857 ();
 DECAPx2_ASAP7_75t_R FILLER_79_861 ();
 DECAPx4_ASAP7_75t_R FILLER_79_875 ();
 DECAPx2_ASAP7_75t_R FILLER_79_893 ();
 FILLER_ASAP7_75t_R FILLER_79_899 ();
 FILLER_ASAP7_75t_R FILLER_79_909 ();
 DECAPx2_ASAP7_75t_R FILLER_79_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_924 ();
 DECAPx4_ASAP7_75t_R FILLER_79_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_937 ();
 FILLER_ASAP7_75t_R FILLER_79_941 ();
 DECAPx2_ASAP7_75t_R FILLER_79_955 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_961 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_974 ();
 DECAPx1_ASAP7_75t_R FILLER_79_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_79_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_79_1049 ();
 DECAPx1_ASAP7_75t_R FILLER_79_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_79_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_79_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_79_1136 ();
 FILLER_ASAP7_75t_R FILLER_79_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_79_1158 ();
 DECAPx4_ASAP7_75t_R FILLER_79_1188 ();
 FILLER_ASAP7_75t_R FILLER_79_1198 ();
 FILLER_ASAP7_75t_R FILLER_79_1226 ();
 FILLER_ASAP7_75t_R FILLER_79_1234 ();
 DECAPx2_ASAP7_75t_R FILLER_79_1246 ();
 FILLER_ASAP7_75t_R FILLER_79_1278 ();
 FILLER_ASAP7_75t_R FILLER_79_1286 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_79_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1305 ();
 FILLER_ASAP7_75t_R FILLER_79_1312 ();
 DECAPx6_ASAP7_75t_R FILLER_79_1340 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_1354 ();
 DECAPx1_ASAP7_75t_R FILLER_79_1361 ();
 FILLER_ASAP7_75t_R FILLER_79_1368 ();
 FILLER_ASAP7_75t_R FILLER_79_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_80_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_8 ();
 DECAPx2_ASAP7_75t_R FILLER_80_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_43 ();
 DECAPx4_ASAP7_75t_R FILLER_80_52 ();
 FILLER_ASAP7_75t_R FILLER_80_88 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_100 ();
 DECAPx6_ASAP7_75t_R FILLER_80_109 ();
 FILLER_ASAP7_75t_R FILLER_80_129 ();
 DECAPx2_ASAP7_75t_R FILLER_80_137 ();
 FILLER_ASAP7_75t_R FILLER_80_153 ();
 FILLER_ASAP7_75t_R FILLER_80_163 ();
 FILLER_ASAP7_75t_R FILLER_80_172 ();
 FILLER_ASAP7_75t_R FILLER_80_180 ();
 DECAPx10_ASAP7_75t_R FILLER_80_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_210 ();
 FILLER_ASAP7_75t_R FILLER_80_217 ();
 FILLER_ASAP7_75t_R FILLER_80_225 ();
 DECAPx2_ASAP7_75t_R FILLER_80_230 ();
 DECAPx1_ASAP7_75t_R FILLER_80_242 ();
 FILLER_ASAP7_75t_R FILLER_80_252 ();
 DECAPx1_ASAP7_75t_R FILLER_80_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_268 ();
 FILLER_ASAP7_75t_R FILLER_80_276 ();
 FILLER_ASAP7_75t_R FILLER_80_304 ();
 FILLER_ASAP7_75t_R FILLER_80_312 ();
 DECAPx10_ASAP7_75t_R FILLER_80_317 ();
 DECAPx2_ASAP7_75t_R FILLER_80_339 ();
 DECAPx1_ASAP7_75t_R FILLER_80_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_352 ();
 DECAPx6_ASAP7_75t_R FILLER_80_356 ();
 FILLER_ASAP7_75t_R FILLER_80_376 ();
 DECAPx2_ASAP7_75t_R FILLER_80_384 ();
 FILLER_ASAP7_75t_R FILLER_80_390 ();
 DECAPx1_ASAP7_75t_R FILLER_80_398 ();
 DECAPx2_ASAP7_75t_R FILLER_80_405 ();
 DECAPx2_ASAP7_75t_R FILLER_80_437 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_443 ();
 FILLER_ASAP7_75t_R FILLER_80_460 ();
 DECAPx2_ASAP7_75t_R FILLER_80_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_470 ();
 FILLER_ASAP7_75t_R FILLER_80_478 ();
 DECAPx2_ASAP7_75t_R FILLER_80_486 ();
 FILLER_ASAP7_75t_R FILLER_80_492 ();
 DECAPx1_ASAP7_75t_R FILLER_80_500 ();
 FILLER_ASAP7_75t_R FILLER_80_510 ();
 FILLER_ASAP7_75t_R FILLER_80_515 ();
 DECAPx1_ASAP7_75t_R FILLER_80_520 ();
 DECAPx1_ASAP7_75t_R FILLER_80_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_534 ();
 DECAPx2_ASAP7_75t_R FILLER_80_538 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_544 ();
 FILLER_ASAP7_75t_R FILLER_80_559 ();
 DECAPx2_ASAP7_75t_R FILLER_80_583 ();
 DECAPx4_ASAP7_75t_R FILLER_80_597 ();
 FILLER_ASAP7_75t_R FILLER_80_611 ();
 DECAPx2_ASAP7_75t_R FILLER_80_621 ();
 FILLER_ASAP7_75t_R FILLER_80_627 ();
 FILLER_ASAP7_75t_R FILLER_80_639 ();
 DECAPx2_ASAP7_75t_R FILLER_80_647 ();
 DECAPx2_ASAP7_75t_R FILLER_80_660 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_666 ();
 FILLER_ASAP7_75t_R FILLER_80_676 ();
 FILLER_ASAP7_75t_R FILLER_80_698 ();
 DECAPx1_ASAP7_75t_R FILLER_80_706 ();
 FILLER_ASAP7_75t_R FILLER_80_717 ();
 DECAPx6_ASAP7_75t_R FILLER_80_726 ();
 FILLER_ASAP7_75t_R FILLER_80_749 ();
 FILLER_ASAP7_75t_R FILLER_80_757 ();
 DECAPx2_ASAP7_75t_R FILLER_80_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_771 ();
 FILLER_ASAP7_75t_R FILLER_80_779 ();
 FILLER_ASAP7_75t_R FILLER_80_787 ();
 DECAPx2_ASAP7_75t_R FILLER_80_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_801 ();
 DECAPx2_ASAP7_75t_R FILLER_80_814 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_820 ();
 DECAPx2_ASAP7_75t_R FILLER_80_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_841 ();
 FILLER_ASAP7_75t_R FILLER_80_854 ();
 DECAPx2_ASAP7_75t_R FILLER_80_859 ();
 DECAPx4_ASAP7_75t_R FILLER_80_873 ();
 FILLER_ASAP7_75t_R FILLER_80_895 ();
 FILLER_ASAP7_75t_R FILLER_80_903 ();
 DECAPx2_ASAP7_75t_R FILLER_80_913 ();
 FILLER_ASAP7_75t_R FILLER_80_919 ();
 DECAPx2_ASAP7_75t_R FILLER_80_933 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_939 ();
 FILLER_ASAP7_75t_R FILLER_80_950 ();
 DECAPx2_ASAP7_75t_R FILLER_80_960 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_966 ();
 FILLER_ASAP7_75t_R FILLER_80_975 ();
 DECAPx2_ASAP7_75t_R FILLER_80_984 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_990 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1015 ();
 FILLER_ASAP7_75t_R FILLER_80_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1028 ();
 FILLER_ASAP7_75t_R FILLER_80_1034 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_80_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1104 ();
 FILLER_ASAP7_75t_R FILLER_80_1110 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1115 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_80_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1168 ();
 FILLER_ASAP7_75t_R FILLER_80_1177 ();
 FILLER_ASAP7_75t_R FILLER_80_1182 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1208 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1217 ();
 FILLER_ASAP7_75t_R FILLER_80_1231 ();
 FILLER_ASAP7_75t_R FILLER_80_1236 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1241 ();
 DECAPx1_ASAP7_75t_R FILLER_80_1263 ();
 DECAPx6_ASAP7_75t_R FILLER_80_1270 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1321 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1327 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1331 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_1337 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1346 ();
 DECAPx2_ASAP7_75t_R FILLER_80_1359 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_1365 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_1374 ();
 DECAPx4_ASAP7_75t_R FILLER_81_2 ();
 FILLER_ASAP7_75t_R FILLER_81_12 ();
 DECAPx1_ASAP7_75t_R FILLER_81_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_24 ();
 DECAPx1_ASAP7_75t_R FILLER_81_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_32 ();
 FILLER_ASAP7_75t_R FILLER_81_36 ();
 FILLER_ASAP7_75t_R FILLER_81_44 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_81_54 ();
 FILLER_ASAP7_75t_R FILLER_81_63 ();
 DECAPx10_ASAP7_75t_R FILLER_81_71 ();
 DECAPx6_ASAP7_75t_R FILLER_81_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_107 ();
 FILLER_ASAP7_75t_R FILLER_81_114 ();
 FILLER_ASAP7_75t_R FILLER_81_123 ();
 DECAPx4_ASAP7_75t_R FILLER_81_151 ();
 FILLER_ASAP7_75t_R FILLER_81_161 ();
 DECAPx1_ASAP7_75t_R FILLER_81_173 ();
 DECAPx4_ASAP7_75t_R FILLER_81_183 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_81_193 ();
 FILLER_ASAP7_75t_R FILLER_81_202 ();
 DECAPx10_ASAP7_75t_R FILLER_81_207 ();
 DECAPx4_ASAP7_75t_R FILLER_81_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_239 ();
 DECAPx6_ASAP7_75t_R FILLER_81_246 ();
 DECAPx1_ASAP7_75t_R FILLER_81_260 ();
 FILLER_ASAP7_75t_R FILLER_81_270 ();
 FILLER_ASAP7_75t_R FILLER_81_294 ();
 FILLER_ASAP7_75t_R FILLER_81_302 ();
 DECAPx2_ASAP7_75t_R FILLER_81_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_313 ();
 DECAPx10_ASAP7_75t_R FILLER_81_320 ();
 DECAPx4_ASAP7_75t_R FILLER_81_342 ();
 FILLER_ASAP7_75t_R FILLER_81_352 ();
 DECAPx6_ASAP7_75t_R FILLER_81_362 ();
 DECAPx1_ASAP7_75t_R FILLER_81_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_380 ();
 DECAPx4_ASAP7_75t_R FILLER_81_389 ();
 DECAPx6_ASAP7_75t_R FILLER_81_402 ();
 DECAPx2_ASAP7_75t_R FILLER_81_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_428 ();
 FILLER_ASAP7_75t_R FILLER_81_435 ();
 FILLER_ASAP7_75t_R FILLER_81_443 ();
 DECAPx1_ASAP7_75t_R FILLER_81_451 ();
 DECAPx2_ASAP7_75t_R FILLER_81_481 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_81_487 ();
 DECAPx2_ASAP7_75t_R FILLER_81_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_522 ();
 DECAPx1_ASAP7_75t_R FILLER_81_545 ();
 FILLER_ASAP7_75t_R FILLER_81_555 ();
 FILLER_ASAP7_75t_R FILLER_81_563 ();
 FILLER_ASAP7_75t_R FILLER_81_572 ();
 DECAPx1_ASAP7_75t_R FILLER_81_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_588 ();
 FILLER_ASAP7_75t_R FILLER_81_615 ();
 DECAPx2_ASAP7_75t_R FILLER_81_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_633 ();
 DECAPx1_ASAP7_75t_R FILLER_81_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_645 ();
 DECAPx1_ASAP7_75t_R FILLER_81_649 ();
 DECAPx2_ASAP7_75t_R FILLER_81_673 ();
 FILLER_ASAP7_75t_R FILLER_81_686 ();
 DECAPx6_ASAP7_75t_R FILLER_81_693 ();
 DECAPx1_ASAP7_75t_R FILLER_81_707 ();
 FILLER_ASAP7_75t_R FILLER_81_717 ();
 DECAPx2_ASAP7_75t_R FILLER_81_725 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_81_731 ();
 DECAPx6_ASAP7_75t_R FILLER_81_743 ();
 DECAPx1_ASAP7_75t_R FILLER_81_757 ();
 FILLER_ASAP7_75t_R FILLER_81_768 ();
 DECAPx2_ASAP7_75t_R FILLER_81_778 ();
 FILLER_ASAP7_75t_R FILLER_81_784 ();
 DECAPx2_ASAP7_75t_R FILLER_81_792 ();
 FILLER_ASAP7_75t_R FILLER_81_798 ();
 FILLER_ASAP7_75t_R FILLER_81_808 ();
 FILLER_ASAP7_75t_R FILLER_81_817 ();
 DECAPx10_ASAP7_75t_R FILLER_81_822 ();
 DECAPx10_ASAP7_75t_R FILLER_81_844 ();
 DECAPx4_ASAP7_75t_R FILLER_81_866 ();
 DECAPx2_ASAP7_75t_R FILLER_81_884 ();
 FILLER_ASAP7_75t_R FILLER_81_890 ();
 DECAPx4_ASAP7_75t_R FILLER_81_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_910 ();
 FILLER_ASAP7_75t_R FILLER_81_923 ();
 FILLER_ASAP7_75t_R FILLER_81_927 ();
 FILLER_ASAP7_75t_R FILLER_81_939 ();
 DECAPx1_ASAP7_75t_R FILLER_81_944 ();
 FILLER_ASAP7_75t_R FILLER_81_974 ();
 DECAPx1_ASAP7_75t_R FILLER_81_984 ();
 FILLER_ASAP7_75t_R FILLER_81_994 ();
 DECAPx2_ASAP7_75t_R FILLER_81_1006 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_81_1012 ();
 DECAPx6_ASAP7_75t_R FILLER_81_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_81_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1050 ();
 FILLER_ASAP7_75t_R FILLER_81_1057 ();
 DECAPx6_ASAP7_75t_R FILLER_81_1067 ();
 DECAPx1_ASAP7_75t_R FILLER_81_1081 ();
 FILLER_ASAP7_75t_R FILLER_81_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_81_1098 ();
 DECAPx6_ASAP7_75t_R FILLER_81_1120 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_81_1134 ();
 FILLER_ASAP7_75t_R FILLER_81_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1192 ();
 DECAPx4_ASAP7_75t_R FILLER_81_1214 ();
 FILLER_ASAP7_75t_R FILLER_81_1224 ();
 DECAPx2_ASAP7_75t_R FILLER_81_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_81_1300 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_81_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_81_1312 ();
 FILLER_ASAP7_75t_R FILLER_81_1334 ();
 DECAPx1_ASAP7_75t_R FILLER_81_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_1348 ();
 FILLER_ASAP7_75t_R FILLER_81_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_82_2 ();
 DECAPx2_ASAP7_75t_R FILLER_82_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_40 ();
 DECAPx10_ASAP7_75t_R FILLER_82_47 ();
 DECAPx10_ASAP7_75t_R FILLER_82_69 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_91 ();
 DECAPx4_ASAP7_75t_R FILLER_82_97 ();
 FILLER_ASAP7_75t_R FILLER_82_107 ();
 FILLER_ASAP7_75t_R FILLER_82_116 ();
 DECAPx1_ASAP7_75t_R FILLER_82_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_128 ();
 FILLER_ASAP7_75t_R FILLER_82_139 ();
 DECAPx10_ASAP7_75t_R FILLER_82_144 ();
 DECAPx2_ASAP7_75t_R FILLER_82_166 ();
 FILLER_ASAP7_75t_R FILLER_82_172 ();
 DECAPx2_ASAP7_75t_R FILLER_82_180 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_186 ();
 DECAPx2_ASAP7_75t_R FILLER_82_215 ();
 DECAPx4_ASAP7_75t_R FILLER_82_227 ();
 DECAPx2_ASAP7_75t_R FILLER_82_263 ();
 FILLER_ASAP7_75t_R FILLER_82_269 ();
 DECAPx1_ASAP7_75t_R FILLER_82_277 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_287 ();
 FILLER_ASAP7_75t_R FILLER_82_296 ();
 DECAPx1_ASAP7_75t_R FILLER_82_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_308 ();
 FILLER_ASAP7_75t_R FILLER_82_335 ();
 DECAPx1_ASAP7_75t_R FILLER_82_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_349 ();
 FILLER_ASAP7_75t_R FILLER_82_356 ();
 DECAPx2_ASAP7_75t_R FILLER_82_366 ();
 FILLER_ASAP7_75t_R FILLER_82_372 ();
 FILLER_ASAP7_75t_R FILLER_82_382 ();
 FILLER_ASAP7_75t_R FILLER_82_390 ();
 DECAPx1_ASAP7_75t_R FILLER_82_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_402 ();
 DECAPx1_ASAP7_75t_R FILLER_82_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_413 ();
 DECAPx4_ASAP7_75t_R FILLER_82_417 ();
 DECAPx1_ASAP7_75t_R FILLER_82_453 ();
 FILLER_ASAP7_75t_R FILLER_82_460 ();
 FILLER_ASAP7_75t_R FILLER_82_464 ();
 FILLER_ASAP7_75t_R FILLER_82_472 ();
 FILLER_ASAP7_75t_R FILLER_82_500 ();
 FILLER_ASAP7_75t_R FILLER_82_524 ();
 DECAPx4_ASAP7_75t_R FILLER_82_536 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_546 ();
 FILLER_ASAP7_75t_R FILLER_82_575 ();
 FILLER_ASAP7_75t_R FILLER_82_580 ();
 FILLER_ASAP7_75t_R FILLER_82_593 ();
 FILLER_ASAP7_75t_R FILLER_82_602 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_610 ();
 FILLER_ASAP7_75t_R FILLER_82_620 ();
 DECAPx2_ASAP7_75t_R FILLER_82_625 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_631 ();
 DECAPx6_ASAP7_75t_R FILLER_82_654 ();
 DECAPx2_ASAP7_75t_R FILLER_82_668 ();
 DECAPx4_ASAP7_75t_R FILLER_82_684 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_694 ();
 DECAPx4_ASAP7_75t_R FILLER_82_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_713 ();
 FILLER_ASAP7_75t_R FILLER_82_720 ();
 DECAPx10_ASAP7_75t_R FILLER_82_728 ();
 DECAPx2_ASAP7_75t_R FILLER_82_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_756 ();
 DECAPx6_ASAP7_75t_R FILLER_82_764 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_778 ();
 DECAPx6_ASAP7_75t_R FILLER_82_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_802 ();
 DECAPx6_ASAP7_75t_R FILLER_82_806 ();
 DECAPx2_ASAP7_75t_R FILLER_82_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_826 ();
 DECAPx1_ASAP7_75t_R FILLER_82_833 ();
 DECAPx6_ASAP7_75t_R FILLER_82_840 ();
 DECAPx2_ASAP7_75t_R FILLER_82_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_860 ();
 DECAPx10_ASAP7_75t_R FILLER_82_871 ();
 DECAPx6_ASAP7_75t_R FILLER_82_893 ();
 DECAPx1_ASAP7_75t_R FILLER_82_907 ();
 DECAPx6_ASAP7_75t_R FILLER_82_917 ();
 DECAPx2_ASAP7_75t_R FILLER_82_941 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_947 ();
 DECAPx2_ASAP7_75t_R FILLER_82_956 ();
 DECAPx10_ASAP7_75t_R FILLER_82_965 ();
 DECAPx10_ASAP7_75t_R FILLER_82_987 ();
 FILLER_ASAP7_75t_R FILLER_82_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1035 ();
 FILLER_ASAP7_75t_R FILLER_82_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1069 ();
 FILLER_ASAP7_75t_R FILLER_82_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1103 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_1133 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_1139 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1154 ();
 FILLER_ASAP7_75t_R FILLER_82_1163 ();
 FILLER_ASAP7_75t_R FILLER_82_1171 ();
 FILLER_ASAP7_75t_R FILLER_82_1183 ();
 FILLER_ASAP7_75t_R FILLER_82_1188 ();
 FILLER_ASAP7_75t_R FILLER_82_1200 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1216 ();
 FILLER_ASAP7_75t_R FILLER_82_1223 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1257 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1262 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_82_1274 ();
 DECAPx6_ASAP7_75t_R FILLER_82_1302 ();
 DECAPx1_ASAP7_75t_R FILLER_82_1320 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1324 ();
 DECAPx6_ASAP7_75t_R FILLER_82_1333 ();
 DECAPx2_ASAP7_75t_R FILLER_82_1347 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_1353 ();
 FILLER_ASAP7_75t_R FILLER_82_1360 ();
 FILLER_ASAP7_75t_R FILLER_82_1367 ();
 FILLER_ASAP7_75t_R FILLER_82_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_83_2 ();
 FILLER_ASAP7_75t_R FILLER_83_8 ();
 DECAPx2_ASAP7_75t_R FILLER_83_16 ();
 DECAPx10_ASAP7_75t_R FILLER_83_25 ();
 DECAPx2_ASAP7_75t_R FILLER_83_47 ();
 DECAPx4_ASAP7_75t_R FILLER_83_61 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_71 ();
 DECAPx2_ASAP7_75t_R FILLER_83_80 ();
 FILLER_ASAP7_75t_R FILLER_83_92 ();
 FILLER_ASAP7_75t_R FILLER_83_100 ();
 FILLER_ASAP7_75t_R FILLER_83_108 ();
 DECAPx4_ASAP7_75t_R FILLER_83_117 ();
 DECAPx6_ASAP7_75t_R FILLER_83_133 ();
 DECAPx1_ASAP7_75t_R FILLER_83_147 ();
 FILLER_ASAP7_75t_R FILLER_83_157 ();
 DECAPx2_ASAP7_75t_R FILLER_83_165 ();
 DECAPx2_ASAP7_75t_R FILLER_83_179 ();
 FILLER_ASAP7_75t_R FILLER_83_185 ();
 FILLER_ASAP7_75t_R FILLER_83_193 ();
 DECAPx4_ASAP7_75t_R FILLER_83_201 ();
 DECAPx2_ASAP7_75t_R FILLER_83_237 ();
 FILLER_ASAP7_75t_R FILLER_83_243 ();
 DECAPx2_ASAP7_75t_R FILLER_83_251 ();
 DECAPx1_ASAP7_75t_R FILLER_83_283 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_295 ();
 DECAPx4_ASAP7_75t_R FILLER_83_306 ();
 FILLER_ASAP7_75t_R FILLER_83_316 ();
 DECAPx2_ASAP7_75t_R FILLER_83_324 ();
 FILLER_ASAP7_75t_R FILLER_83_336 ();
 FILLER_ASAP7_75t_R FILLER_83_346 ();
 FILLER_ASAP7_75t_R FILLER_83_354 ();
 DECAPx4_ASAP7_75t_R FILLER_83_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_372 ();
 DECAPx6_ASAP7_75t_R FILLER_83_380 ();
 DECAPx1_ASAP7_75t_R FILLER_83_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_398 ();
 DECAPx4_ASAP7_75t_R FILLER_83_425 ();
 DECAPx1_ASAP7_75t_R FILLER_83_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_461 ();
 FILLER_ASAP7_75t_R FILLER_83_469 ();
 FILLER_ASAP7_75t_R FILLER_83_478 ();
 FILLER_ASAP7_75t_R FILLER_83_487 ();
 DECAPx2_ASAP7_75t_R FILLER_83_495 ();
 DECAPx4_ASAP7_75t_R FILLER_83_504 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_514 ();
 FILLER_ASAP7_75t_R FILLER_83_524 ();
 DECAPx2_ASAP7_75t_R FILLER_83_536 ();
 FILLER_ASAP7_75t_R FILLER_83_542 ();
 FILLER_ASAP7_75t_R FILLER_83_550 ();
 DECAPx2_ASAP7_75t_R FILLER_83_558 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_564 ();
 FILLER_ASAP7_75t_R FILLER_83_573 ();
 DECAPx4_ASAP7_75t_R FILLER_83_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_591 ();
 DECAPx2_ASAP7_75t_R FILLER_83_598 ();
 DECAPx2_ASAP7_75t_R FILLER_83_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_613 ();
 DECAPx4_ASAP7_75t_R FILLER_83_620 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_630 ();
 DECAPx10_ASAP7_75t_R FILLER_83_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_658 ();
 DECAPx6_ASAP7_75t_R FILLER_83_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_678 ();
 FILLER_ASAP7_75t_R FILLER_83_686 ();
 DECAPx1_ASAP7_75t_R FILLER_83_696 ();
 FILLER_ASAP7_75t_R FILLER_83_722 ();
 DECAPx2_ASAP7_75t_R FILLER_83_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_739 ();
 FILLER_ASAP7_75t_R FILLER_83_760 ();
 FILLER_ASAP7_75t_R FILLER_83_771 ();
 DECAPx10_ASAP7_75t_R FILLER_83_779 ();
 DECAPx2_ASAP7_75t_R FILLER_83_801 ();
 FILLER_ASAP7_75t_R FILLER_83_807 ();
 DECAPx1_ASAP7_75t_R FILLER_83_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_821 ();
 DECAPx2_ASAP7_75t_R FILLER_83_848 ();
 FILLER_ASAP7_75t_R FILLER_83_854 ();
 DECAPx10_ASAP7_75t_R FILLER_83_862 ();
 DECAPx2_ASAP7_75t_R FILLER_83_891 ();
 FILLER_ASAP7_75t_R FILLER_83_897 ();
 DECAPx4_ASAP7_75t_R FILLER_83_902 ();
 DECAPx2_ASAP7_75t_R FILLER_83_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_924 ();
 DECAPx10_ASAP7_75t_R FILLER_83_927 ();
 DECAPx2_ASAP7_75t_R FILLER_83_949 ();
 DECAPx2_ASAP7_75t_R FILLER_83_963 ();
 DECAPx2_ASAP7_75t_R FILLER_83_975 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_981 ();
 DECAPx4_ASAP7_75t_R FILLER_83_987 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1023 ();
 FILLER_ASAP7_75t_R FILLER_83_1029 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_1041 ();
 DECAPx1_ASAP7_75t_R FILLER_83_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_83_1060 ();
 FILLER_ASAP7_75t_R FILLER_83_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_83_1097 ();
 FILLER_ASAP7_75t_R FILLER_83_1117 ();
 FILLER_ASAP7_75t_R FILLER_83_1125 ();
 FILLER_ASAP7_75t_R FILLER_83_1137 ();
 DECAPx1_ASAP7_75t_R FILLER_83_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_83_1193 ();
 FILLER_ASAP7_75t_R FILLER_83_1199 ();
 DECAPx4_ASAP7_75t_R FILLER_83_1227 ();
 FILLER_ASAP7_75t_R FILLER_83_1237 ();
 DECAPx6_ASAP7_75t_R FILLER_83_1242 ();
 FILLER_ASAP7_75t_R FILLER_83_1282 ();
 FILLER_ASAP7_75t_R FILLER_83_1290 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_1295 ();
 FILLER_ASAP7_75t_R FILLER_83_1324 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_1329 ();
 FILLER_ASAP7_75t_R FILLER_83_1342 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_1352 ();
 FILLER_ASAP7_75t_R FILLER_83_1361 ();
 FILLER_ASAP7_75t_R FILLER_83_1366 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_1374 ();
 DECAPx10_ASAP7_75t_R FILLER_84_2 ();
 DECAPx2_ASAP7_75t_R FILLER_84_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_30 ();
 FILLER_ASAP7_75t_R FILLER_84_34 ();
 DECAPx2_ASAP7_75t_R FILLER_84_42 ();
 FILLER_ASAP7_75t_R FILLER_84_54 ();
 FILLER_ASAP7_75t_R FILLER_84_64 ();
 FILLER_ASAP7_75t_R FILLER_84_92 ();
 DECAPx2_ASAP7_75t_R FILLER_84_102 ();
 FILLER_ASAP7_75t_R FILLER_84_108 ();
 FILLER_ASAP7_75t_R FILLER_84_117 ();
 FILLER_ASAP7_75t_R FILLER_84_126 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_84_134 ();
 DECAPx1_ASAP7_75t_R FILLER_84_143 ();
 FILLER_ASAP7_75t_R FILLER_84_150 ();
 DECAPx1_ASAP7_75t_R FILLER_84_160 ();
 FILLER_ASAP7_75t_R FILLER_84_170 ();
 DECAPx2_ASAP7_75t_R FILLER_84_175 ();
 FILLER_ASAP7_75t_R FILLER_84_181 ();
 DECAPx2_ASAP7_75t_R FILLER_84_209 ();
 DECAPx1_ASAP7_75t_R FILLER_84_221 ();
 DECAPx10_ASAP7_75t_R FILLER_84_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_250 ();
 DECAPx2_ASAP7_75t_R FILLER_84_254 ();
 FILLER_ASAP7_75t_R FILLER_84_260 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_84_268 ();
 DECAPx2_ASAP7_75t_R FILLER_84_274 ();
 FILLER_ASAP7_75t_R FILLER_84_280 ();
 DECAPx10_ASAP7_75t_R FILLER_84_285 ();
 DECAPx6_ASAP7_75t_R FILLER_84_307 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_84_321 ();
 DECAPx2_ASAP7_75t_R FILLER_84_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_333 ();
 DECAPx10_ASAP7_75t_R FILLER_84_340 ();
 DECAPx4_ASAP7_75t_R FILLER_84_362 ();
 FILLER_ASAP7_75t_R FILLER_84_372 ();
 DECAPx2_ASAP7_75t_R FILLER_84_380 ();
 DECAPx4_ASAP7_75t_R FILLER_84_392 ();
 DECAPx10_ASAP7_75t_R FILLER_84_408 ();
 DECAPx6_ASAP7_75t_R FILLER_84_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_444 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_84_451 ();
 FILLER_ASAP7_75t_R FILLER_84_460 ();
 FILLER_ASAP7_75t_R FILLER_84_464 ();
 FILLER_ASAP7_75t_R FILLER_84_469 ();
 FILLER_ASAP7_75t_R FILLER_84_478 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_84_486 ();
 DECAPx6_ASAP7_75t_R FILLER_84_492 ();
 DECAPx4_ASAP7_75t_R FILLER_84_514 ();
 DECAPx6_ASAP7_75t_R FILLER_84_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_546 ();
 FILLER_ASAP7_75t_R FILLER_84_553 ();
 FILLER_ASAP7_75t_R FILLER_84_561 ();
 DECAPx10_ASAP7_75t_R FILLER_84_566 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_84_588 ();
 DECAPx6_ASAP7_75t_R FILLER_84_597 ();
 DECAPx2_ASAP7_75t_R FILLER_84_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_617 ();
 DECAPx6_ASAP7_75t_R FILLER_84_624 ();
 DECAPx6_ASAP7_75t_R FILLER_84_645 ();
 DECAPx4_ASAP7_75t_R FILLER_84_666 ();
 DECAPx1_ASAP7_75t_R FILLER_84_683 ();
 DECAPx1_ASAP7_75t_R FILLER_84_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_701 ();
 FILLER_ASAP7_75t_R FILLER_84_710 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_84_719 ();
 FILLER_ASAP7_75t_R FILLER_84_730 ();
 DECAPx2_ASAP7_75t_R FILLER_84_743 ();
 FILLER_ASAP7_75t_R FILLER_84_749 ();
 DECAPx4_ASAP7_75t_R FILLER_84_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_773 ();
 DECAPx2_ASAP7_75t_R FILLER_84_780 ();
 DECAPx4_ASAP7_75t_R FILLER_84_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_799 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_84_806 ();
 DECAPx2_ASAP7_75t_R FILLER_84_812 ();
 DECAPx1_ASAP7_75t_R FILLER_84_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_832 ();
 DECAPx1_ASAP7_75t_R FILLER_84_839 ();
 DECAPx2_ASAP7_75t_R FILLER_84_849 ();
 FILLER_ASAP7_75t_R FILLER_84_881 ();
 FILLER_ASAP7_75t_R FILLER_84_909 ();
 DECAPx6_ASAP7_75t_R FILLER_84_937 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_84_951 ();
 FILLER_ASAP7_75t_R FILLER_84_968 ();
 DECAPx6_ASAP7_75t_R FILLER_84_996 ();
 DECAPx1_ASAP7_75t_R FILLER_84_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_84_1042 ();
 FILLER_ASAP7_75t_R FILLER_84_1048 ();
 DECAPx4_ASAP7_75t_R FILLER_84_1061 ();
 FILLER_ASAP7_75t_R FILLER_84_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1089 ();
 DECAPx4_ASAP7_75t_R FILLER_84_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_84_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1147 ();
 FILLER_ASAP7_75t_R FILLER_84_1174 ();
 DECAPx1_ASAP7_75t_R FILLER_84_1184 ();
 DECAPx1_ASAP7_75t_R FILLER_84_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1196 ();
 FILLER_ASAP7_75t_R FILLER_84_1205 ();
 FILLER_ASAP7_75t_R FILLER_84_1215 ();
 DECAPx6_ASAP7_75t_R FILLER_84_1220 ();
 DECAPx1_ASAP7_75t_R FILLER_84_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1238 ();
 DECAPx4_ASAP7_75t_R FILLER_84_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_1256 ();
 FILLER_ASAP7_75t_R FILLER_84_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_84_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_84_1304 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_84_1310 ();
 DECAPx4_ASAP7_75t_R FILLER_84_1339 ();
 FILLER_ASAP7_75t_R FILLER_84_1375 ();
 DECAPx4_ASAP7_75t_R FILLER_85_2 ();
 FILLER_ASAP7_75t_R FILLER_85_12 ();
 DECAPx2_ASAP7_75t_R FILLER_85_20 ();
 FILLER_ASAP7_75t_R FILLER_85_26 ();
 FILLER_ASAP7_75t_R FILLER_85_54 ();
 DECAPx2_ASAP7_75t_R FILLER_85_62 ();
 FILLER_ASAP7_75t_R FILLER_85_68 ();
 DECAPx1_ASAP7_75t_R FILLER_85_76 ();
 FILLER_ASAP7_75t_R FILLER_85_83 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_91 ();
 FILLER_ASAP7_75t_R FILLER_85_100 ();
 DECAPx2_ASAP7_75t_R FILLER_85_128 ();
 FILLER_ASAP7_75t_R FILLER_85_134 ();
 DECAPx6_ASAP7_75t_R FILLER_85_142 ();
 FILLER_ASAP7_75t_R FILLER_85_156 ();
 FILLER_ASAP7_75t_R FILLER_85_164 ();
 DECAPx6_ASAP7_75t_R FILLER_85_173 ();
 DECAPx1_ASAP7_75t_R FILLER_85_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_191 ();
 FILLER_ASAP7_75t_R FILLER_85_198 ();
 DECAPx4_ASAP7_75t_R FILLER_85_203 ();
 FILLER_ASAP7_75t_R FILLER_85_213 ();
 DECAPx2_ASAP7_75t_R FILLER_85_218 ();
 FILLER_ASAP7_75t_R FILLER_85_224 ();
 DECAPx4_ASAP7_75t_R FILLER_85_232 ();
 FILLER_ASAP7_75t_R FILLER_85_242 ();
 DECAPx6_ASAP7_75t_R FILLER_85_250 ();
 DECAPx6_ASAP7_75t_R FILLER_85_267 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_281 ();
 DECAPx6_ASAP7_75t_R FILLER_85_290 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_310 ();
 FILLER_ASAP7_75t_R FILLER_85_319 ();
 DECAPx2_ASAP7_75t_R FILLER_85_327 ();
 DECAPx1_ASAP7_75t_R FILLER_85_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_340 ();
 DECAPx1_ASAP7_75t_R FILLER_85_347 ();
 DECAPx6_ASAP7_75t_R FILLER_85_357 ();
 FILLER_ASAP7_75t_R FILLER_85_371 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_381 ();
 DECAPx2_ASAP7_75t_R FILLER_85_392 ();
 FILLER_ASAP7_75t_R FILLER_85_398 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_426 ();
 DECAPx1_ASAP7_75t_R FILLER_85_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_439 ();
 FILLER_ASAP7_75t_R FILLER_85_443 ();
 DECAPx2_ASAP7_75t_R FILLER_85_453 ();
 FILLER_ASAP7_75t_R FILLER_85_459 ();
 DECAPx4_ASAP7_75t_R FILLER_85_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_497 ();
 FILLER_ASAP7_75t_R FILLER_85_504 ();
 DECAPx2_ASAP7_75t_R FILLER_85_514 ();
 FILLER_ASAP7_75t_R FILLER_85_520 ();
 FILLER_ASAP7_75t_R FILLER_85_528 ();
 DECAPx4_ASAP7_75t_R FILLER_85_536 ();
 FILLER_ASAP7_75t_R FILLER_85_546 ();
 DECAPx2_ASAP7_75t_R FILLER_85_574 ();
 FILLER_ASAP7_75t_R FILLER_85_580 ();
 DECAPx2_ASAP7_75t_R FILLER_85_585 ();
 FILLER_ASAP7_75t_R FILLER_85_591 ();
 DECAPx1_ASAP7_75t_R FILLER_85_599 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_609 ();
 FILLER_ASAP7_75t_R FILLER_85_621 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_649 ();
 FILLER_ASAP7_75t_R FILLER_85_658 ();
 DECAPx1_ASAP7_75t_R FILLER_85_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_671 ();
 DECAPx4_ASAP7_75t_R FILLER_85_684 ();
 DECAPx2_ASAP7_75t_R FILLER_85_714 ();
 FILLER_ASAP7_75t_R FILLER_85_729 ();
 DECAPx10_ASAP7_75t_R FILLER_85_737 ();
 DECAPx4_ASAP7_75t_R FILLER_85_759 ();
 FILLER_ASAP7_75t_R FILLER_85_769 ();
 FILLER_ASAP7_75t_R FILLER_85_797 ();
 DECAPx2_ASAP7_75t_R FILLER_85_825 ();
 FILLER_ASAP7_75t_R FILLER_85_831 ();
 DECAPx1_ASAP7_75t_R FILLER_85_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_843 ();
 DECAPx4_ASAP7_75t_R FILLER_85_850 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_860 ();
 FILLER_ASAP7_75t_R FILLER_85_869 ();
 DECAPx2_ASAP7_75t_R FILLER_85_874 ();
 FILLER_ASAP7_75t_R FILLER_85_890 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_898 ();
 DECAPx2_ASAP7_75t_R FILLER_85_911 ();
 FILLER_ASAP7_75t_R FILLER_85_923 ();
 FILLER_ASAP7_75t_R FILLER_85_927 ();
 DECAPx1_ASAP7_75t_R FILLER_85_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_943 ();
 DECAPx2_ASAP7_75t_R FILLER_85_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_956 ();
 DECAPx6_ASAP7_75t_R FILLER_85_964 ();
 DECAPx1_ASAP7_75t_R FILLER_85_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_982 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_990 ();
 DECAPx6_ASAP7_75t_R FILLER_85_1005 ();
 FILLER_ASAP7_75t_R FILLER_85_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1093 ();
 FILLER_ASAP7_75t_R FILLER_85_1099 ();
 DECAPx4_ASAP7_75t_R FILLER_85_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_85_1143 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_85_1188 ();
 DECAPx4_ASAP7_75t_R FILLER_85_1210 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_1220 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1229 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_1235 ();
 FILLER_ASAP7_75t_R FILLER_85_1246 ();
 DECAPx6_ASAP7_75t_R FILLER_85_1254 ();
 FILLER_ASAP7_75t_R FILLER_85_1268 ();
 DECAPx4_ASAP7_75t_R FILLER_85_1273 ();
 DECAPx4_ASAP7_75t_R FILLER_85_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1296 ();
 DECAPx2_ASAP7_75t_R FILLER_85_1304 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1310 ();
 FILLER_ASAP7_75t_R FILLER_85_1318 ();
 FILLER_ASAP7_75t_R FILLER_85_1326 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_1331 ();
 DECAPx6_ASAP7_75t_R FILLER_85_1337 ();
 FILLER_ASAP7_75t_R FILLER_85_1351 ();
 DECAPx1_ASAP7_75t_R FILLER_85_1360 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_1364 ();
 FILLER_ASAP7_75t_R FILLER_85_1368 ();
 FILLER_ASAP7_75t_R FILLER_85_1375 ();
 FILLER_ASAP7_75t_R FILLER_86_2 ();
 FILLER_ASAP7_75t_R FILLER_86_30 ();
 DECAPx1_ASAP7_75t_R FILLER_86_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_42 ();
 DECAPx10_ASAP7_75t_R FILLER_86_46 ();
 DECAPx10_ASAP7_75t_R FILLER_86_68 ();
 DECAPx4_ASAP7_75t_R FILLER_86_90 ();
 FILLER_ASAP7_75t_R FILLER_86_100 ();
 FILLER_ASAP7_75t_R FILLER_86_108 ();
 FILLER_ASAP7_75t_R FILLER_86_117 ();
 FILLER_ASAP7_75t_R FILLER_86_126 ();
 DECAPx6_ASAP7_75t_R FILLER_86_131 ();
 DECAPx1_ASAP7_75t_R FILLER_86_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_149 ();
 DECAPx10_ASAP7_75t_R FILLER_86_156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_178 ();
 DECAPx4_ASAP7_75t_R FILLER_86_187 ();
 DECAPx1_ASAP7_75t_R FILLER_86_200 ();
 DECAPx2_ASAP7_75t_R FILLER_86_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_216 ();
 FILLER_ASAP7_75t_R FILLER_86_223 ();
 FILLER_ASAP7_75t_R FILLER_86_233 ();
 FILLER_ASAP7_75t_R FILLER_86_261 ();
 DECAPx2_ASAP7_75t_R FILLER_86_266 ();
 FILLER_ASAP7_75t_R FILLER_86_272 ();
 DECAPx2_ASAP7_75t_R FILLER_86_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_306 ();
 FILLER_ASAP7_75t_R FILLER_86_333 ();
 DECAPx2_ASAP7_75t_R FILLER_86_361 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_367 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_396 ();
 FILLER_ASAP7_75t_R FILLER_86_405 ();
 DECAPx2_ASAP7_75t_R FILLER_86_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_419 ();
 FILLER_ASAP7_75t_R FILLER_86_446 ();
 DECAPx4_ASAP7_75t_R FILLER_86_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_461 ();
 FILLER_ASAP7_75t_R FILLER_86_464 ();
 DECAPx1_ASAP7_75t_R FILLER_86_469 ();
 FILLER_ASAP7_75t_R FILLER_86_479 ();
 FILLER_ASAP7_75t_R FILLER_86_507 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_515 ();
 DECAPx4_ASAP7_75t_R FILLER_86_526 ();
 FILLER_ASAP7_75t_R FILLER_86_536 ();
 DECAPx6_ASAP7_75t_R FILLER_86_544 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_558 ();
 FILLER_ASAP7_75t_R FILLER_86_587 ();
 FILLER_ASAP7_75t_R FILLER_86_597 ();
 DECAPx1_ASAP7_75t_R FILLER_86_602 ();
 FILLER_ASAP7_75t_R FILLER_86_614 ();
 FILLER_ASAP7_75t_R FILLER_86_622 ();
 DECAPx4_ASAP7_75t_R FILLER_86_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_637 ();
 DECAPx4_ASAP7_75t_R FILLER_86_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_651 ();
 DECAPx6_ASAP7_75t_R FILLER_86_658 ();
 FILLER_ASAP7_75t_R FILLER_86_672 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_696 ();
 FILLER_ASAP7_75t_R FILLER_86_707 ();
 FILLER_ASAP7_75t_R FILLER_86_729 ();
 FILLER_ASAP7_75t_R FILLER_86_737 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_747 ();
 DECAPx6_ASAP7_75t_R FILLER_86_760 ();
 DECAPx2_ASAP7_75t_R FILLER_86_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_780 ();
 DECAPx6_ASAP7_75t_R FILLER_86_787 ();
 DECAPx2_ASAP7_75t_R FILLER_86_801 ();
 DECAPx6_ASAP7_75t_R FILLER_86_813 ();
 FILLER_ASAP7_75t_R FILLER_86_827 ();
 DECAPx2_ASAP7_75t_R FILLER_86_855 ();
 FILLER_ASAP7_75t_R FILLER_86_861 ();
 DECAPx10_ASAP7_75t_R FILLER_86_869 ();
 DECAPx1_ASAP7_75t_R FILLER_86_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_895 ();
 DECAPx6_ASAP7_75t_R FILLER_86_899 ();
 DECAPx2_ASAP7_75t_R FILLER_86_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_919 ();
 FILLER_ASAP7_75t_R FILLER_86_923 ();
 FILLER_ASAP7_75t_R FILLER_86_930 ();
 FILLER_ASAP7_75t_R FILLER_86_942 ();
 DECAPx1_ASAP7_75t_R FILLER_86_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_958 ();
 FILLER_ASAP7_75t_R FILLER_86_969 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_974 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_1003 ();
 DECAPx6_ASAP7_75t_R FILLER_86_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_86_1037 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_1047 ();
 DECAPx6_ASAP7_75t_R FILLER_86_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1073 ();
 FILLER_ASAP7_75t_R FILLER_86_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1100 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1119 ();
 DECAPx6_ASAP7_75t_R FILLER_86_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1201 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1213 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1217 ();
 FILLER_ASAP7_75t_R FILLER_86_1223 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1232 ();
 FILLER_ASAP7_75t_R FILLER_86_1242 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1252 ();
 FILLER_ASAP7_75t_R FILLER_86_1258 ();
 FILLER_ASAP7_75t_R FILLER_86_1267 ();
 FILLER_ASAP7_75t_R FILLER_86_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_86_1324 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1346 ();
 FILLER_ASAP7_75t_R FILLER_86_1352 ();
 DECAPx1_ASAP7_75t_R FILLER_86_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_1365 ();
 DECAPx2_ASAP7_75t_R FILLER_86_1369 ();
 FILLER_ASAP7_75t_R FILLER_86_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_87_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_8 ();
 DECAPx1_ASAP7_75t_R FILLER_87_15 ();
 DECAPx10_ASAP7_75t_R FILLER_87_22 ();
 DECAPx2_ASAP7_75t_R FILLER_87_44 ();
 FILLER_ASAP7_75t_R FILLER_87_56 ();
 FILLER_ASAP7_75t_R FILLER_87_84 ();
 DECAPx10_ASAP7_75t_R FILLER_87_92 ();
 DECAPx1_ASAP7_75t_R FILLER_87_114 ();
 FILLER_ASAP7_75t_R FILLER_87_124 ();
 DECAPx4_ASAP7_75t_R FILLER_87_132 ();
 FILLER_ASAP7_75t_R FILLER_87_168 ();
 FILLER_ASAP7_75t_R FILLER_87_196 ();
 FILLER_ASAP7_75t_R FILLER_87_204 ();
 DECAPx1_ASAP7_75t_R FILLER_87_214 ();
 DECAPx4_ASAP7_75t_R FILLER_87_226 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_236 ();
 DECAPx1_ASAP7_75t_R FILLER_87_245 ();
 DECAPx6_ASAP7_75t_R FILLER_87_252 ();
 DECAPx1_ASAP7_75t_R FILLER_87_274 ();
 DECAPx1_ASAP7_75t_R FILLER_87_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_288 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_292 ();
 FILLER_ASAP7_75t_R FILLER_87_303 ();
 FILLER_ASAP7_75t_R FILLER_87_327 ();
 DECAPx6_ASAP7_75t_R FILLER_87_332 ();
 DECAPx1_ASAP7_75t_R FILLER_87_346 ();
 DECAPx6_ASAP7_75t_R FILLER_87_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_367 ();
 FILLER_ASAP7_75t_R FILLER_87_374 ();
 FILLER_ASAP7_75t_R FILLER_87_382 ();
 DECAPx10_ASAP7_75t_R FILLER_87_387 ();
 DECAPx1_ASAP7_75t_R FILLER_87_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_413 ();
 DECAPx2_ASAP7_75t_R FILLER_87_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_423 ();
 DECAPx2_ASAP7_75t_R FILLER_87_430 ();
 FILLER_ASAP7_75t_R FILLER_87_442 ();
 DECAPx4_ASAP7_75t_R FILLER_87_450 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_460 ();
 DECAPx2_ASAP7_75t_R FILLER_87_469 ();
 DECAPx2_ASAP7_75t_R FILLER_87_478 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_484 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_493 ();
 DECAPx6_ASAP7_75t_R FILLER_87_499 ();
 DECAPx2_ASAP7_75t_R FILLER_87_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_519 ();
 FILLER_ASAP7_75t_R FILLER_87_528 ();
 FILLER_ASAP7_75t_R FILLER_87_536 ();
 DECAPx4_ASAP7_75t_R FILLER_87_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_574 ();
 DECAPx4_ASAP7_75t_R FILLER_87_578 ();
 DECAPx4_ASAP7_75t_R FILLER_87_604 ();
 DECAPx2_ASAP7_75t_R FILLER_87_620 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_626 ();
 FILLER_ASAP7_75t_R FILLER_87_635 ();
 FILLER_ASAP7_75t_R FILLER_87_647 ();
 DECAPx4_ASAP7_75t_R FILLER_87_655 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_665 ();
 DECAPx2_ASAP7_75t_R FILLER_87_675 ();
 FILLER_ASAP7_75t_R FILLER_87_701 ();
 DECAPx10_ASAP7_75t_R FILLER_87_713 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_735 ();
 FILLER_ASAP7_75t_R FILLER_87_746 ();
 DECAPx2_ASAP7_75t_R FILLER_87_756 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_772 ();
 DECAPx4_ASAP7_75t_R FILLER_87_782 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_800 ();
 DECAPx4_ASAP7_75t_R FILLER_87_811 ();
 DECAPx6_ASAP7_75t_R FILLER_87_829 ();
 DECAPx6_ASAP7_75t_R FILLER_87_846 ();
 DECAPx1_ASAP7_75t_R FILLER_87_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_864 ();
 FILLER_ASAP7_75t_R FILLER_87_875 ();
 DECAPx1_ASAP7_75t_R FILLER_87_885 ();
 FILLER_ASAP7_75t_R FILLER_87_901 ();
 DECAPx1_ASAP7_75t_R FILLER_87_909 ();
 FILLER_ASAP7_75t_R FILLER_87_923 ();
 DECAPx1_ASAP7_75t_R FILLER_87_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_931 ();
 DECAPx6_ASAP7_75t_R FILLER_87_938 ();
 DECAPx2_ASAP7_75t_R FILLER_87_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_958 ();
 DECAPx1_ASAP7_75t_R FILLER_87_985 ();
 FILLER_ASAP7_75t_R FILLER_87_995 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1000 ();
 FILLER_ASAP7_75t_R FILLER_87_1006 ();
 FILLER_ASAP7_75t_R FILLER_87_1018 ();
 DECAPx1_ASAP7_75t_R FILLER_87_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1030 ();
 DECAPx4_ASAP7_75t_R FILLER_87_1039 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1059 ();
 DECAPx6_ASAP7_75t_R FILLER_87_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1089 ();
 FILLER_ASAP7_75t_R FILLER_87_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_87_1103 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_1125 ();
 FILLER_ASAP7_75t_R FILLER_87_1135 ();
 FILLER_ASAP7_75t_R FILLER_87_1140 ();
 DECAPx6_ASAP7_75t_R FILLER_87_1148 ();
 DECAPx1_ASAP7_75t_R FILLER_87_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1193 ();
 FILLER_ASAP7_75t_R FILLER_87_1225 ();
 FILLER_ASAP7_75t_R FILLER_87_1234 ();
 DECAPx4_ASAP7_75t_R FILLER_87_1248 ();
 DECAPx1_ASAP7_75t_R FILLER_87_1284 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_1294 ();
 DECAPx4_ASAP7_75t_R FILLER_87_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_87_1318 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_1324 ();
 DECAPx1_ASAP7_75t_R FILLER_87_1330 ();
 DECAPx1_ASAP7_75t_R FILLER_87_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_1348 ();
 FILLER_ASAP7_75t_R FILLER_87_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_88_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_24 ();
 DECAPx1_ASAP7_75t_R FILLER_88_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_37 ();
 DECAPx1_ASAP7_75t_R FILLER_88_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_68 ();
 DECAPx1_ASAP7_75t_R FILLER_88_75 ();
 FILLER_ASAP7_75t_R FILLER_88_105 ();
 DECAPx2_ASAP7_75t_R FILLER_88_113 ();
 FILLER_ASAP7_75t_R FILLER_88_145 ();
 DECAPx1_ASAP7_75t_R FILLER_88_153 ();
 DECAPx6_ASAP7_75t_R FILLER_88_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_174 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_181 ();
 DECAPx6_ASAP7_75t_R FILLER_88_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_201 ();
 DECAPx4_ASAP7_75t_R FILLER_88_209 ();
 DECAPx10_ASAP7_75t_R FILLER_88_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_247 ();
 DECAPx1_ASAP7_75t_R FILLER_88_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_258 ();
 FILLER_ASAP7_75t_R FILLER_88_265 ();
 DECAPx1_ASAP7_75t_R FILLER_88_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_279 ();
 FILLER_ASAP7_75t_R FILLER_88_286 ();
 FILLER_ASAP7_75t_R FILLER_88_295 ();
 FILLER_ASAP7_75t_R FILLER_88_303 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_327 ();
 DECAPx6_ASAP7_75t_R FILLER_88_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_350 ();
 FILLER_ASAP7_75t_R FILLER_88_357 ();
 DECAPx1_ASAP7_75t_R FILLER_88_365 ();
 FILLER_ASAP7_75t_R FILLER_88_376 ();
 DECAPx4_ASAP7_75t_R FILLER_88_381 ();
 FILLER_ASAP7_75t_R FILLER_88_394 ();
 DECAPx6_ASAP7_75t_R FILLER_88_402 ();
 DECAPx2_ASAP7_75t_R FILLER_88_416 ();
 DECAPx4_ASAP7_75t_R FILLER_88_425 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_435 ();
 FILLER_ASAP7_75t_R FILLER_88_452 ();
 FILLER_ASAP7_75t_R FILLER_88_460 ();
 FILLER_ASAP7_75t_R FILLER_88_464 ();
 DECAPx6_ASAP7_75t_R FILLER_88_472 ();
 DECAPx1_ASAP7_75t_R FILLER_88_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_490 ();
 DECAPx2_ASAP7_75t_R FILLER_88_497 ();
 DECAPx1_ASAP7_75t_R FILLER_88_509 ();
 DECAPx2_ASAP7_75t_R FILLER_88_516 ();
 DECAPx4_ASAP7_75t_R FILLER_88_528 ();
 DECAPx2_ASAP7_75t_R FILLER_88_544 ();
 FILLER_ASAP7_75t_R FILLER_88_550 ();
 DECAPx10_ASAP7_75t_R FILLER_88_555 ();
 DECAPx2_ASAP7_75t_R FILLER_88_577 ();
 DECAPx10_ASAP7_75t_R FILLER_88_586 ();
 DECAPx10_ASAP7_75t_R FILLER_88_608 ();
 DECAPx1_ASAP7_75t_R FILLER_88_630 ();
 DECAPx4_ASAP7_75t_R FILLER_88_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_658 ();
 DECAPx2_ASAP7_75t_R FILLER_88_667 ();
 FILLER_ASAP7_75t_R FILLER_88_673 ();
 FILLER_ASAP7_75t_R FILLER_88_695 ();
 FILLER_ASAP7_75t_R FILLER_88_705 ();
 DECAPx1_ASAP7_75t_R FILLER_88_727 ();
 DECAPx4_ASAP7_75t_R FILLER_88_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_747 ();
 FILLER_ASAP7_75t_R FILLER_88_754 ();
 FILLER_ASAP7_75t_R FILLER_88_776 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_789 ();
 DECAPx1_ASAP7_75t_R FILLER_88_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_805 ();
 DECAPx2_ASAP7_75t_R FILLER_88_816 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_822 ();
 DECAPx2_ASAP7_75t_R FILLER_88_835 ();
 FILLER_ASAP7_75t_R FILLER_88_841 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_853 ();
 DECAPx6_ASAP7_75t_R FILLER_88_862 ();
 DECAPx2_ASAP7_75t_R FILLER_88_876 ();
 DECAPx4_ASAP7_75t_R FILLER_88_894 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_904 ();
 FILLER_ASAP7_75t_R FILLER_88_933 ();
 FILLER_ASAP7_75t_R FILLER_88_945 ();
 DECAPx6_ASAP7_75t_R FILLER_88_953 ();
 DECAPx2_ASAP7_75t_R FILLER_88_967 ();
 DECAPx10_ASAP7_75t_R FILLER_88_976 ();
 DECAPx6_ASAP7_75t_R FILLER_88_998 ();
 FILLER_ASAP7_75t_R FILLER_88_1038 ();
 FILLER_ASAP7_75t_R FILLER_88_1046 ();
 FILLER_ASAP7_75t_R FILLER_88_1074 ();
 FILLER_ASAP7_75t_R FILLER_88_1098 ();
 FILLER_ASAP7_75t_R FILLER_88_1107 ();
 DECAPx4_ASAP7_75t_R FILLER_88_1116 ();
 FILLER_ASAP7_75t_R FILLER_88_1126 ();
 DECAPx6_ASAP7_75t_R FILLER_88_1131 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1149 ();
 FILLER_ASAP7_75t_R FILLER_88_1157 ();
 FILLER_ASAP7_75t_R FILLER_88_1165 ();
 FILLER_ASAP7_75t_R FILLER_88_1179 ();
 FILLER_ASAP7_75t_R FILLER_88_1187 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1192 ();
 FILLER_ASAP7_75t_R FILLER_88_1206 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1214 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_88_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1251 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1258 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_88_1276 ();
 DECAPx1_ASAP7_75t_R FILLER_88_1308 ();
 FILLER_ASAP7_75t_R FILLER_88_1338 ();
 DECAPx4_ASAP7_75t_R FILLER_88_1343 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_1353 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_1362 ();
 FILLER_ASAP7_75t_R FILLER_88_1368 ();
 FILLER_ASAP7_75t_R FILLER_88_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_89_2 ();
 FILLER_ASAP7_75t_R FILLER_89_8 ();
 DECAPx1_ASAP7_75t_R FILLER_89_16 ();
 FILLER_ASAP7_75t_R FILLER_89_46 ();
 FILLER_ASAP7_75t_R FILLER_89_54 ();
 DECAPx1_ASAP7_75t_R FILLER_89_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_63 ();
 FILLER_ASAP7_75t_R FILLER_89_70 ();
 DECAPx2_ASAP7_75t_R FILLER_89_75 ();
 FILLER_ASAP7_75t_R FILLER_89_81 ();
 DECAPx1_ASAP7_75t_R FILLER_89_89 ();
 DECAPx1_ASAP7_75t_R FILLER_89_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_100 ();
 DECAPx2_ASAP7_75t_R FILLER_89_127 ();
 DECAPx10_ASAP7_75t_R FILLER_89_136 ();
 DECAPx1_ASAP7_75t_R FILLER_89_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_162 ();
 FILLER_ASAP7_75t_R FILLER_89_169 ();
 DECAPx10_ASAP7_75t_R FILLER_89_174 ();
 DECAPx10_ASAP7_75t_R FILLER_89_196 ();
 DECAPx2_ASAP7_75t_R FILLER_89_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_224 ();
 DECAPx2_ASAP7_75t_R FILLER_89_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_237 ();
 FILLER_ASAP7_75t_R FILLER_89_264 ();
 DECAPx6_ASAP7_75t_R FILLER_89_272 ();
 FILLER_ASAP7_75t_R FILLER_89_286 ();
 DECAPx4_ASAP7_75t_R FILLER_89_296 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_306 ();
 DECAPx6_ASAP7_75t_R FILLER_89_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_331 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_338 ();
 DECAPx1_ASAP7_75t_R FILLER_89_344 ();
 DECAPx4_ASAP7_75t_R FILLER_89_374 ();
 FILLER_ASAP7_75t_R FILLER_89_390 ();
 DECAPx2_ASAP7_75t_R FILLER_89_400 ();
 FILLER_ASAP7_75t_R FILLER_89_406 ();
 FILLER_ASAP7_75t_R FILLER_89_414 ();
 DECAPx1_ASAP7_75t_R FILLER_89_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_426 ();
 DECAPx4_ASAP7_75t_R FILLER_89_434 ();
 FILLER_ASAP7_75t_R FILLER_89_444 ();
 DECAPx2_ASAP7_75t_R FILLER_89_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_458 ();
 FILLER_ASAP7_75t_R FILLER_89_462 ();
 FILLER_ASAP7_75t_R FILLER_89_486 ();
 DECAPx6_ASAP7_75t_R FILLER_89_514 ();
 DECAPx4_ASAP7_75t_R FILLER_89_534 ();
 FILLER_ASAP7_75t_R FILLER_89_544 ();
 FILLER_ASAP7_75t_R FILLER_89_552 ();
 DECAPx10_ASAP7_75t_R FILLER_89_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_582 ();
 DECAPx4_ASAP7_75t_R FILLER_89_590 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_600 ();
 DECAPx1_ASAP7_75t_R FILLER_89_609 ();
 FILLER_ASAP7_75t_R FILLER_89_621 ();
 DECAPx1_ASAP7_75t_R FILLER_89_626 ();
 DECAPx2_ASAP7_75t_R FILLER_89_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_642 ();
 DECAPx2_ASAP7_75t_R FILLER_89_650 ();
 FILLER_ASAP7_75t_R FILLER_89_656 ();
 DECAPx1_ASAP7_75t_R FILLER_89_666 ();
 FILLER_ASAP7_75t_R FILLER_89_690 ();
 DECAPx1_ASAP7_75t_R FILLER_89_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_702 ();
 FILLER_ASAP7_75t_R FILLER_89_710 ();
 FILLER_ASAP7_75t_R FILLER_89_723 ();
 DECAPx6_ASAP7_75t_R FILLER_89_741 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_755 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_767 ();
 FILLER_ASAP7_75t_R FILLER_89_780 ();
 DECAPx2_ASAP7_75t_R FILLER_89_788 ();
 DECAPx4_ASAP7_75t_R FILLER_89_797 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_807 ();
 FILLER_ASAP7_75t_R FILLER_89_817 ();
 DECAPx1_ASAP7_75t_R FILLER_89_825 ();
 FILLER_ASAP7_75t_R FILLER_89_839 ();
 FILLER_ASAP7_75t_R FILLER_89_855 ();
 DECAPx2_ASAP7_75t_R FILLER_89_871 ();
 FILLER_ASAP7_75t_R FILLER_89_877 ();
 FILLER_ASAP7_75t_R FILLER_89_889 ();
 DECAPx2_ASAP7_75t_R FILLER_89_903 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_909 ();
 DECAPx2_ASAP7_75t_R FILLER_89_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_924 ();
 FILLER_ASAP7_75t_R FILLER_89_927 ();
 FILLER_ASAP7_75t_R FILLER_89_932 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_960 ();
 DECAPx2_ASAP7_75t_R FILLER_89_966 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_972 ();
 DECAPx6_ASAP7_75t_R FILLER_89_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_999 ();
 DECAPx6_ASAP7_75t_R FILLER_89_1006 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_89_1030 ();
 DECAPx6_ASAP7_75t_R FILLER_89_1037 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1057 ();
 FILLER_ASAP7_75t_R FILLER_89_1064 ();
 DECAPx6_ASAP7_75t_R FILLER_89_1069 ();
 FILLER_ASAP7_75t_R FILLER_89_1083 ();
 FILLER_ASAP7_75t_R FILLER_89_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1145 ();
 DECAPx6_ASAP7_75t_R FILLER_89_1172 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_1186 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1196 ();
 FILLER_ASAP7_75t_R FILLER_89_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1218 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_89_1263 ();
 FILLER_ASAP7_75t_R FILLER_89_1292 ();
 FILLER_ASAP7_75t_R FILLER_89_1300 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1305 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_1311 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1318 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_1324 ();
 FILLER_ASAP7_75t_R FILLER_89_1335 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1343 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_1349 ();
 FILLER_ASAP7_75t_R FILLER_89_1355 ();
 DECAPx2_ASAP7_75t_R FILLER_89_1364 ();
 FILLER_ASAP7_75t_R FILLER_89_1375 ();
 FILLER_ASAP7_75t_R FILLER_90_2 ();
 FILLER_ASAP7_75t_R FILLER_90_30 ();
 FILLER_ASAP7_75t_R FILLER_90_38 ();
 DECAPx10_ASAP7_75t_R FILLER_90_43 ();
 DECAPx1_ASAP7_75t_R FILLER_90_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_69 ();
 DECAPx10_ASAP7_75t_R FILLER_90_76 ();
 DECAPx6_ASAP7_75t_R FILLER_90_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_112 ();
 FILLER_ASAP7_75t_R FILLER_90_119 ();
 DECAPx6_ASAP7_75t_R FILLER_90_124 ();
 DECAPx2_ASAP7_75t_R FILLER_90_144 ();
 FILLER_ASAP7_75t_R FILLER_90_150 ();
 FILLER_ASAP7_75t_R FILLER_90_178 ();
 DECAPx4_ASAP7_75t_R FILLER_90_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_196 ();
 FILLER_ASAP7_75t_R FILLER_90_205 ();
 DECAPx1_ASAP7_75t_R FILLER_90_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_217 ();
 DECAPx4_ASAP7_75t_R FILLER_90_224 ();
 FILLER_ASAP7_75t_R FILLER_90_241 ();
 DECAPx1_ASAP7_75t_R FILLER_90_249 ();
 DECAPx6_ASAP7_75t_R FILLER_90_256 ();
 DECAPx1_ASAP7_75t_R FILLER_90_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_274 ();
 DECAPx10_ASAP7_75t_R FILLER_90_281 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_303 ();
 FILLER_ASAP7_75t_R FILLER_90_312 ();
 FILLER_ASAP7_75t_R FILLER_90_325 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_353 ();
 DECAPx1_ASAP7_75t_R FILLER_90_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_382 ();
 FILLER_ASAP7_75t_R FILLER_90_405 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_421 ();
 DECAPx2_ASAP7_75t_R FILLER_90_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_438 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_445 ();
 DECAPx2_ASAP7_75t_R FILLER_90_456 ();
 FILLER_ASAP7_75t_R FILLER_90_464 ();
 FILLER_ASAP7_75t_R FILLER_90_474 ();
 FILLER_ASAP7_75t_R FILLER_90_502 ();
 DECAPx4_ASAP7_75t_R FILLER_90_507 ();
 FILLER_ASAP7_75t_R FILLER_90_517 ();
 FILLER_ASAP7_75t_R FILLER_90_541 ();
 DECAPx6_ASAP7_75t_R FILLER_90_569 ();
 FILLER_ASAP7_75t_R FILLER_90_590 ();
 FILLER_ASAP7_75t_R FILLER_90_606 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_614 ();
 DECAPx6_ASAP7_75t_R FILLER_90_625 ();
 DECAPx1_ASAP7_75t_R FILLER_90_639 ();
 FILLER_ASAP7_75t_R FILLER_90_653 ();
 FILLER_ASAP7_75t_R FILLER_90_663 ();
 FILLER_ASAP7_75t_R FILLER_90_671 ();
 DECAPx2_ASAP7_75t_R FILLER_90_693 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_699 ();
 DECAPx1_ASAP7_75t_R FILLER_90_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_720 ();
 DECAPx10_ASAP7_75t_R FILLER_90_737 ();
 DECAPx6_ASAP7_75t_R FILLER_90_759 ();
 DECAPx1_ASAP7_75t_R FILLER_90_773 ();
 DECAPx10_ASAP7_75t_R FILLER_90_783 ();
 DECAPx10_ASAP7_75t_R FILLER_90_805 ();
 DECAPx2_ASAP7_75t_R FILLER_90_827 ();
 DECAPx10_ASAP7_75t_R FILLER_90_841 ();
 DECAPx1_ASAP7_75t_R FILLER_90_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_867 ();
 FILLER_ASAP7_75t_R FILLER_90_874 ();
 FILLER_ASAP7_75t_R FILLER_90_902 ();
 DECAPx1_ASAP7_75t_R FILLER_90_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_911 ();
 DECAPx10_ASAP7_75t_R FILLER_90_918 ();
 DECAPx1_ASAP7_75t_R FILLER_90_940 ();
 FILLER_ASAP7_75t_R FILLER_90_950 ();
 DECAPx1_ASAP7_75t_R FILLER_90_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_959 ();
 FILLER_ASAP7_75t_R FILLER_90_986 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1018 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1023 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1064 ();
 FILLER_ASAP7_75t_R FILLER_90_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1083 ();
 FILLER_ASAP7_75t_R FILLER_90_1094 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1102 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1123 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_1127 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1185 ();
 FILLER_ASAP7_75t_R FILLER_90_1215 ();
 FILLER_ASAP7_75t_R FILLER_90_1223 ();
 FILLER_ASAP7_75t_R FILLER_90_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_90_1266 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_1272 ();
 DECAPx4_ASAP7_75t_R FILLER_90_1281 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_90_1303 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_1325 ();
 DECAPx1_ASAP7_75t_R FILLER_90_1334 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_1346 ();
 FILLER_ASAP7_75t_R FILLER_90_1375 ();
 DECAPx1_ASAP7_75t_R FILLER_91_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_6 ();
 DECAPx1_ASAP7_75t_R FILLER_91_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_17 ();
 DECAPx4_ASAP7_75t_R FILLER_91_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_31 ();
 DECAPx4_ASAP7_75t_R FILLER_91_35 ();
 FILLER_ASAP7_75t_R FILLER_91_48 ();
 DECAPx2_ASAP7_75t_R FILLER_91_58 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_64 ();
 FILLER_ASAP7_75t_R FILLER_91_75 ();
 DECAPx4_ASAP7_75t_R FILLER_91_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_93 ();
 DECAPx4_ASAP7_75t_R FILLER_91_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_110 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_114 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_123 ();
 FILLER_ASAP7_75t_R FILLER_91_132 ();
 FILLER_ASAP7_75t_R FILLER_91_160 ();
 FILLER_ASAP7_75t_R FILLER_91_168 ();
 FILLER_ASAP7_75t_R FILLER_91_196 ();
 DECAPx4_ASAP7_75t_R FILLER_91_206 ();
 DECAPx2_ASAP7_75t_R FILLER_91_224 ();
 FILLER_ASAP7_75t_R FILLER_91_238 ();
 DECAPx2_ASAP7_75t_R FILLER_91_246 ();
 DECAPx4_ASAP7_75t_R FILLER_91_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_268 ();
 DECAPx10_ASAP7_75t_R FILLER_91_277 ();
 DECAPx2_ASAP7_75t_R FILLER_91_299 ();
 FILLER_ASAP7_75t_R FILLER_91_313 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_321 ();
 DECAPx10_ASAP7_75t_R FILLER_91_335 ();
 DECAPx1_ASAP7_75t_R FILLER_91_357 ();
 FILLER_ASAP7_75t_R FILLER_91_364 ();
 FILLER_ASAP7_75t_R FILLER_91_392 ();
 DECAPx2_ASAP7_75t_R FILLER_91_416 ();
 DECAPx4_ASAP7_75t_R FILLER_91_428 ();
 DECAPx6_ASAP7_75t_R FILLER_91_444 ();
 DECAPx2_ASAP7_75t_R FILLER_91_458 ();
 DECAPx2_ASAP7_75t_R FILLER_91_470 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_476 ();
 FILLER_ASAP7_75t_R FILLER_91_485 ();
 FILLER_ASAP7_75t_R FILLER_91_493 ();
 DECAPx10_ASAP7_75t_R FILLER_91_498 ();
 DECAPx1_ASAP7_75t_R FILLER_91_520 ();
 DECAPx2_ASAP7_75t_R FILLER_91_532 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_538 ();
 FILLER_ASAP7_75t_R FILLER_91_547 ();
 FILLER_ASAP7_75t_R FILLER_91_557 ();
 DECAPx1_ASAP7_75t_R FILLER_91_567 ();
 FILLER_ASAP7_75t_R FILLER_91_597 ();
 DECAPx2_ASAP7_75t_R FILLER_91_602 ();
 DECAPx4_ASAP7_75t_R FILLER_91_614 ();
 DECAPx10_ASAP7_75t_R FILLER_91_634 ();
 DECAPx2_ASAP7_75t_R FILLER_91_656 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_662 ();
 DECAPx1_ASAP7_75t_R FILLER_91_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_675 ();
 FILLER_ASAP7_75t_R FILLER_91_683 ();
 DECAPx1_ASAP7_75t_R FILLER_91_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_697 ();
 FILLER_ASAP7_75t_R FILLER_91_704 ();
 DECAPx10_ASAP7_75t_R FILLER_91_714 ();
 DECAPx1_ASAP7_75t_R FILLER_91_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_740 ();
 DECAPx1_ASAP7_75t_R FILLER_91_747 ();
 DECAPx1_ASAP7_75t_R FILLER_91_766 ();
 FILLER_ASAP7_75t_R FILLER_91_786 ();
 DECAPx4_ASAP7_75t_R FILLER_91_798 ();
 FILLER_ASAP7_75t_R FILLER_91_815 ();
 DECAPx1_ASAP7_75t_R FILLER_91_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_827 ();
 FILLER_ASAP7_75t_R FILLER_91_834 ();
 DECAPx6_ASAP7_75t_R FILLER_91_839 ();
 DECAPx2_ASAP7_75t_R FILLER_91_853 ();
 DECAPx4_ASAP7_75t_R FILLER_91_862 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_872 ();
 DECAPx2_ASAP7_75t_R FILLER_91_882 ();
 FILLER_ASAP7_75t_R FILLER_91_888 ();
 DECAPx1_ASAP7_75t_R FILLER_91_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_897 ();
 DECAPx6_ASAP7_75t_R FILLER_91_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_924 ();
 DECAPx4_ASAP7_75t_R FILLER_91_927 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_937 ();
 DECAPx4_ASAP7_75t_R FILLER_91_946 ();
 FILLER_ASAP7_75t_R FILLER_91_956 ();
 DECAPx2_ASAP7_75t_R FILLER_91_968 ();
 DECAPx2_ASAP7_75t_R FILLER_91_977 ();
 FILLER_ASAP7_75t_R FILLER_91_983 ();
 FILLER_ASAP7_75t_R FILLER_91_992 ();
 FILLER_ASAP7_75t_R FILLER_91_997 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1009 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_1025 ();
 FILLER_ASAP7_75t_R FILLER_91_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1070 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1089 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1101 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1137 ();
 FILLER_ASAP7_75t_R FILLER_91_1143 ();
 FILLER_ASAP7_75t_R FILLER_91_1148 ();
 DECAPx6_ASAP7_75t_R FILLER_91_1153 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_1167 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1184 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_1190 ();
 DECAPx4_ASAP7_75t_R FILLER_91_1199 ();
 FILLER_ASAP7_75t_R FILLER_91_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1243 ();
 DECAPx2_ASAP7_75t_R FILLER_91_1265 ();
 FILLER_ASAP7_75t_R FILLER_91_1282 ();
 FILLER_ASAP7_75t_R FILLER_91_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_91_1302 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1324 ();
 FILLER_ASAP7_75t_R FILLER_91_1328 ();
 FILLER_ASAP7_75t_R FILLER_91_1340 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1348 ();
 FILLER_ASAP7_75t_R FILLER_91_1357 ();
 DECAPx1_ASAP7_75t_R FILLER_91_1365 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_1369 ();
 FILLER_ASAP7_75t_R FILLER_91_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_92_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_8 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_17 ();
 DECAPx10_ASAP7_75t_R FILLER_92_23 ();
 FILLER_ASAP7_75t_R FILLER_92_51 ();
 DECAPx2_ASAP7_75t_R FILLER_92_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_67 ();
 DECAPx2_ASAP7_75t_R FILLER_92_76 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_82 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_111 ();
 FILLER_ASAP7_75t_R FILLER_92_120 ();
 DECAPx1_ASAP7_75t_R FILLER_92_144 ();
 DECAPx10_ASAP7_75t_R FILLER_92_151 ();
 FILLER_ASAP7_75t_R FILLER_92_173 ();
 DECAPx1_ASAP7_75t_R FILLER_92_181 ();
 DECAPx2_ASAP7_75t_R FILLER_92_188 ();
 FILLER_ASAP7_75t_R FILLER_92_200 ();
 FILLER_ASAP7_75t_R FILLER_92_208 ();
 FILLER_ASAP7_75t_R FILLER_92_216 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_240 ();
 FILLER_ASAP7_75t_R FILLER_92_269 ();
 FILLER_ASAP7_75t_R FILLER_92_279 ();
 DECAPx1_ASAP7_75t_R FILLER_92_287 ();
 DECAPx1_ASAP7_75t_R FILLER_92_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_301 ();
 FILLER_ASAP7_75t_R FILLER_92_308 ();
 DECAPx6_ASAP7_75t_R FILLER_92_313 ();
 DECAPx2_ASAP7_75t_R FILLER_92_327 ();
 DECAPx1_ASAP7_75t_R FILLER_92_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_343 ();
 FILLER_ASAP7_75t_R FILLER_92_347 ();
 DECAPx4_ASAP7_75t_R FILLER_92_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_367 ();
 FILLER_ASAP7_75t_R FILLER_92_374 ();
 FILLER_ASAP7_75t_R FILLER_92_382 ();
 DECAPx1_ASAP7_75t_R FILLER_92_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_391 ();
 DECAPx2_ASAP7_75t_R FILLER_92_398 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_404 ();
 DECAPx1_ASAP7_75t_R FILLER_92_413 ();
 DECAPx6_ASAP7_75t_R FILLER_92_420 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_434 ();
 DECAPx2_ASAP7_75t_R FILLER_92_445 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_451 ();
 FILLER_ASAP7_75t_R FILLER_92_460 ();
 FILLER_ASAP7_75t_R FILLER_92_464 ();
 DECAPx1_ASAP7_75t_R FILLER_92_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_476 ();
 DECAPx10_ASAP7_75t_R FILLER_92_483 ();
 DECAPx1_ASAP7_75t_R FILLER_92_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_515 ();
 FILLER_ASAP7_75t_R FILLER_92_522 ();
 FILLER_ASAP7_75t_R FILLER_92_532 ();
 DECAPx4_ASAP7_75t_R FILLER_92_540 ();
 FILLER_ASAP7_75t_R FILLER_92_553 ();
 DECAPx1_ASAP7_75t_R FILLER_92_558 ();
 DECAPx6_ASAP7_75t_R FILLER_92_568 ();
 FILLER_ASAP7_75t_R FILLER_92_582 ();
 FILLER_ASAP7_75t_R FILLER_92_590 ();
 DECAPx10_ASAP7_75t_R FILLER_92_598 ();
 DECAPx1_ASAP7_75t_R FILLER_92_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_624 ();
 DECAPx6_ASAP7_75t_R FILLER_92_631 ();
 FILLER_ASAP7_75t_R FILLER_92_645 ();
 DECAPx2_ASAP7_75t_R FILLER_92_657 ();
 FILLER_ASAP7_75t_R FILLER_92_663 ();
 FILLER_ASAP7_75t_R FILLER_92_671 ();
 DECAPx2_ASAP7_75t_R FILLER_92_679 ();
 FILLER_ASAP7_75t_R FILLER_92_685 ();
 DECAPx4_ASAP7_75t_R FILLER_92_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_707 ();
 DECAPx4_ASAP7_75t_R FILLER_92_717 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_733 ();
 DECAPx2_ASAP7_75t_R FILLER_92_742 ();
 DECAPx10_ASAP7_75t_R FILLER_92_764 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_786 ();
 DECAPx2_ASAP7_75t_R FILLER_92_795 ();
 FILLER_ASAP7_75t_R FILLER_92_801 ();
 DECAPx2_ASAP7_75t_R FILLER_92_806 ();
 FILLER_ASAP7_75t_R FILLER_92_812 ();
 DECAPx4_ASAP7_75t_R FILLER_92_840 ();
 FILLER_ASAP7_75t_R FILLER_92_850 ();
 FILLER_ASAP7_75t_R FILLER_92_861 ();
 DECAPx6_ASAP7_75t_R FILLER_92_869 ();
 FILLER_ASAP7_75t_R FILLER_92_883 ();
 DECAPx2_ASAP7_75t_R FILLER_92_891 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_897 ();
 FILLER_ASAP7_75t_R FILLER_92_926 ();
 FILLER_ASAP7_75t_R FILLER_92_954 ();
 DECAPx10_ASAP7_75t_R FILLER_92_962 ();
 DECAPx2_ASAP7_75t_R FILLER_92_984 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_990 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1003 ();
 FILLER_ASAP7_75t_R FILLER_92_1009 ();
 DECAPx6_ASAP7_75t_R FILLER_92_1014 ();
 DECAPx4_ASAP7_75t_R FILLER_92_1038 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_1055 ();
 FILLER_ASAP7_75t_R FILLER_92_1064 ();
 DECAPx6_ASAP7_75t_R FILLER_92_1069 ();
 FILLER_ASAP7_75t_R FILLER_92_1109 ();
 DECAPx6_ASAP7_75t_R FILLER_92_1114 ();
 DECAPx6_ASAP7_75t_R FILLER_92_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1148 ();
 DECAPx4_ASAP7_75t_R FILLER_92_1157 ();
 FILLER_ASAP7_75t_R FILLER_92_1193 ();
 DECAPx1_ASAP7_75t_R FILLER_92_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1209 ();
 DECAPx4_ASAP7_75t_R FILLER_92_1217 ();
 FILLER_ASAP7_75t_R FILLER_92_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1252 ();
 FILLER_ASAP7_75t_R FILLER_92_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_92_1264 ();
 FILLER_ASAP7_75t_R FILLER_92_1274 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1282 ();
 FILLER_ASAP7_75t_R FILLER_92_1288 ();
 FILLER_ASAP7_75t_R FILLER_92_1296 ();
 DECAPx2_ASAP7_75t_R FILLER_92_1305 ();
 FILLER_ASAP7_75t_R FILLER_92_1311 ();
 DECAPx1_ASAP7_75t_R FILLER_92_1322 ();
 DECAPx1_ASAP7_75t_R FILLER_92_1334 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1338 ();
 DECAPx1_ASAP7_75t_R FILLER_92_1347 ();
 FILLER_ASAP7_75t_R FILLER_92_1356 ();
 DECAPx1_ASAP7_75t_R FILLER_92_1365 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_1369 ();
 FILLER_ASAP7_75t_R FILLER_92_1375 ();
 DECAPx1_ASAP7_75t_R FILLER_93_2 ();
 DECAPx6_ASAP7_75t_R FILLER_93_32 ();
 DECAPx2_ASAP7_75t_R FILLER_93_46 ();
 DECAPx4_ASAP7_75t_R FILLER_93_58 ();
 DECAPx6_ASAP7_75t_R FILLER_93_74 ();
 FILLER_ASAP7_75t_R FILLER_93_88 ();
 DECAPx1_ASAP7_75t_R FILLER_93_96 ();
 DECAPx2_ASAP7_75t_R FILLER_93_103 ();
 FILLER_ASAP7_75t_R FILLER_93_109 ();
 FILLER_ASAP7_75t_R FILLER_93_119 ();
 DECAPx4_ASAP7_75t_R FILLER_93_129 ();
 FILLER_ASAP7_75t_R FILLER_93_139 ();
 DECAPx2_ASAP7_75t_R FILLER_93_167 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_173 ();
 DECAPx10_ASAP7_75t_R FILLER_93_182 ();
 DECAPx2_ASAP7_75t_R FILLER_93_204 ();
 FILLER_ASAP7_75t_R FILLER_93_210 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_215 ();
 DECAPx2_ASAP7_75t_R FILLER_93_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_246 ();
 DECAPx1_ASAP7_75t_R FILLER_93_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_257 ();
 DECAPx2_ASAP7_75t_R FILLER_93_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_267 ();
 DECAPx1_ASAP7_75t_R FILLER_93_274 ();
 FILLER_ASAP7_75t_R FILLER_93_284 ();
 FILLER_ASAP7_75t_R FILLER_93_312 ();
 DECAPx4_ASAP7_75t_R FILLER_93_317 ();
 FILLER_ASAP7_75t_R FILLER_93_333 ();
 FILLER_ASAP7_75t_R FILLER_93_357 ();
 DECAPx6_ASAP7_75t_R FILLER_93_365 ();
 DECAPx2_ASAP7_75t_R FILLER_93_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_385 ();
 FILLER_ASAP7_75t_R FILLER_93_392 ();
 FILLER_ASAP7_75t_R FILLER_93_400 ();
 DECAPx4_ASAP7_75t_R FILLER_93_428 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_438 ();
 DECAPx4_ASAP7_75t_R FILLER_93_449 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_459 ();
 FILLER_ASAP7_75t_R FILLER_93_484 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_489 ();
 FILLER_ASAP7_75t_R FILLER_93_498 ();
 FILLER_ASAP7_75t_R FILLER_93_526 ();
 DECAPx6_ASAP7_75t_R FILLER_93_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_548 ();
 DECAPx2_ASAP7_75t_R FILLER_93_555 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_583 ();
 DECAPx2_ASAP7_75t_R FILLER_93_593 ();
 FILLER_ASAP7_75t_R FILLER_93_606 ();
 DECAPx2_ASAP7_75t_R FILLER_93_618 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_624 ();
 DECAPx2_ASAP7_75t_R FILLER_93_641 ();
 DECAPx2_ASAP7_75t_R FILLER_93_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_668 ();
 DECAPx2_ASAP7_75t_R FILLER_93_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_681 ();
 FILLER_ASAP7_75t_R FILLER_93_688 ();
 DECAPx4_ASAP7_75t_R FILLER_93_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_710 ();
 DECAPx2_ASAP7_75t_R FILLER_93_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_727 ();
 DECAPx1_ASAP7_75t_R FILLER_93_734 ();
 FILLER_ASAP7_75t_R FILLER_93_746 ();
 FILLER_ASAP7_75t_R FILLER_93_756 ();
 DECAPx6_ASAP7_75t_R FILLER_93_768 ();
 DECAPx2_ASAP7_75t_R FILLER_93_782 ();
 DECAPx2_ASAP7_75t_R FILLER_93_814 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_820 ();
 DECAPx1_ASAP7_75t_R FILLER_93_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_833 ();
 FILLER_ASAP7_75t_R FILLER_93_843 ();
 DECAPx2_ASAP7_75t_R FILLER_93_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_857 ();
 DECAPx2_ASAP7_75t_R FILLER_93_867 ();
 FILLER_ASAP7_75t_R FILLER_93_873 ();
 DECAPx6_ASAP7_75t_R FILLER_93_901 ();
 DECAPx2_ASAP7_75t_R FILLER_93_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_924 ();
 FILLER_ASAP7_75t_R FILLER_93_927 ();
 DECAPx1_ASAP7_75t_R FILLER_93_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_939 ();
 DECAPx4_ASAP7_75t_R FILLER_93_946 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_956 ();
 FILLER_ASAP7_75t_R FILLER_93_969 ();
 FILLER_ASAP7_75t_R FILLER_93_981 ();
 DECAPx4_ASAP7_75t_R FILLER_93_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_996 ();
 FILLER_ASAP7_75t_R FILLER_93_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_93_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1070 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_1077 ();
 DECAPx4_ASAP7_75t_R FILLER_93_1090 ();
 FILLER_ASAP7_75t_R FILLER_93_1100 ();
 FILLER_ASAP7_75t_R FILLER_93_1110 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_1124 ();
 FILLER_ASAP7_75t_R FILLER_93_1137 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_1142 ();
 FILLER_ASAP7_75t_R FILLER_93_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1167 ();
 FILLER_ASAP7_75t_R FILLER_93_1173 ();
 DECAPx4_ASAP7_75t_R FILLER_93_1181 ();
 FILLER_ASAP7_75t_R FILLER_93_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1203 ();
 DECAPx4_ASAP7_75t_R FILLER_93_1225 ();
 DECAPx2_ASAP7_75t_R FILLER_93_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1249 ();
 FILLER_ASAP7_75t_R FILLER_93_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_93_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_1291 ();
 FILLER_ASAP7_75t_R FILLER_93_1302 ();
 FILLER_ASAP7_75t_R FILLER_93_1310 ();
 DECAPx1_ASAP7_75t_R FILLER_93_1338 ();
 FILLER_ASAP7_75t_R FILLER_93_1347 ();
 FILLER_ASAP7_75t_R FILLER_93_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_94_2 ();
 DECAPx2_ASAP7_75t_R FILLER_94_14 ();
 DECAPx2_ASAP7_75t_R FILLER_94_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_32 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_36 ();
 DECAPx2_ASAP7_75t_R FILLER_94_47 ();
 DECAPx10_ASAP7_75t_R FILLER_94_59 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_81 ();
 DECAPx2_ASAP7_75t_R FILLER_94_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_96 ();
 DECAPx10_ASAP7_75t_R FILLER_94_100 ();
 DECAPx6_ASAP7_75t_R FILLER_94_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_136 ();
 FILLER_ASAP7_75t_R FILLER_94_143 ();
 DECAPx2_ASAP7_75t_R FILLER_94_151 ();
 FILLER_ASAP7_75t_R FILLER_94_157 ();
 FILLER_ASAP7_75t_R FILLER_94_185 ();
 DECAPx4_ASAP7_75t_R FILLER_94_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_200 ();
 FILLER_ASAP7_75t_R FILLER_94_207 ();
 FILLER_ASAP7_75t_R FILLER_94_215 ();
 DECAPx10_ASAP7_75t_R FILLER_94_243 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_265 ();
 FILLER_ASAP7_75t_R FILLER_94_290 ();
 DECAPx1_ASAP7_75t_R FILLER_94_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_302 ();
 FILLER_ASAP7_75t_R FILLER_94_309 ();
 FILLER_ASAP7_75t_R FILLER_94_317 ();
 DECAPx1_ASAP7_75t_R FILLER_94_329 ();
 FILLER_ASAP7_75t_R FILLER_94_339 ();
 DECAPx2_ASAP7_75t_R FILLER_94_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_373 ();
 DECAPx1_ASAP7_75t_R FILLER_94_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_404 ();
 DECAPx2_ASAP7_75t_R FILLER_94_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_433 ();
 DECAPx1_ASAP7_75t_R FILLER_94_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_441 ();
 DECAPx2_ASAP7_75t_R FILLER_94_448 ();
 FILLER_ASAP7_75t_R FILLER_94_460 ();
 DECAPx2_ASAP7_75t_R FILLER_94_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_470 ();
 DECAPx2_ASAP7_75t_R FILLER_94_497 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_503 ();
 DECAPx1_ASAP7_75t_R FILLER_94_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_516 ();
 FILLER_ASAP7_75t_R FILLER_94_520 ();
 DECAPx6_ASAP7_75t_R FILLER_94_525 ();
 DECAPx2_ASAP7_75t_R FILLER_94_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_545 ();
 DECAPx6_ASAP7_75t_R FILLER_94_572 ();
 FILLER_ASAP7_75t_R FILLER_94_592 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_597 ();
 FILLER_ASAP7_75t_R FILLER_94_626 ();
 FILLER_ASAP7_75t_R FILLER_94_654 ();
 DECAPx2_ASAP7_75t_R FILLER_94_659 ();
 FILLER_ASAP7_75t_R FILLER_94_665 ();
 DECAPx2_ASAP7_75t_R FILLER_94_683 ();
 FILLER_ASAP7_75t_R FILLER_94_689 ();
 DECAPx4_ASAP7_75t_R FILLER_94_699 ();
 FILLER_ASAP7_75t_R FILLER_94_709 ();
 DECAPx10_ASAP7_75t_R FILLER_94_721 ();
 FILLER_ASAP7_75t_R FILLER_94_751 ();
 DECAPx2_ASAP7_75t_R FILLER_94_759 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_765 ();
 DECAPx2_ASAP7_75t_R FILLER_94_774 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_780 ();
 FILLER_ASAP7_75t_R FILLER_94_790 ();
 DECAPx6_ASAP7_75t_R FILLER_94_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_812 ();
 DECAPx6_ASAP7_75t_R FILLER_94_820 ();
 DECAPx6_ASAP7_75t_R FILLER_94_843 ();
 FILLER_ASAP7_75t_R FILLER_94_865 ();
 DECAPx2_ASAP7_75t_R FILLER_94_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_879 ();
 DECAPx1_ASAP7_75t_R FILLER_94_886 ();
 DECAPx10_ASAP7_75t_R FILLER_94_893 ();
 DECAPx2_ASAP7_75t_R FILLER_94_915 ();
 FILLER_ASAP7_75t_R FILLER_94_921 ();
 DECAPx2_ASAP7_75t_R FILLER_94_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_935 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_939 ();
 FILLER_ASAP7_75t_R FILLER_94_954 ();
 FILLER_ASAP7_75t_R FILLER_94_982 ();
 DECAPx6_ASAP7_75t_R FILLER_94_991 ();
 FILLER_ASAP7_75t_R FILLER_94_1005 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1017 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1038 ();
 FILLER_ASAP7_75t_R FILLER_94_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1059 ();
 FILLER_ASAP7_75t_R FILLER_94_1070 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1082 ();
 FILLER_ASAP7_75t_R FILLER_94_1090 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1106 ();
 FILLER_ASAP7_75t_R FILLER_94_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_94_1144 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_1166 ();
 DECAPx6_ASAP7_75t_R FILLER_94_1176 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1205 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_1220 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1224 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_1234 ();
 FILLER_ASAP7_75t_R FILLER_94_1243 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1248 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_1254 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_94_1276 ();
 FILLER_ASAP7_75t_R FILLER_94_1294 ();
 DECAPx4_ASAP7_75t_R FILLER_94_1299 ();
 FILLER_ASAP7_75t_R FILLER_94_1309 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1318 ();
 FILLER_ASAP7_75t_R FILLER_94_1325 ();
 FILLER_ASAP7_75t_R FILLER_94_1332 ();
 FILLER_ASAP7_75t_R FILLER_94_1339 ();
 FILLER_ASAP7_75t_R FILLER_94_1346 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1356 ();
 DECAPx1_ASAP7_75t_R FILLER_94_1366 ();
 FILLER_ASAP7_75t_R FILLER_94_1375 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_95_2 ();
 DECAPx2_ASAP7_75t_R FILLER_95_31 ();
 FILLER_ASAP7_75t_R FILLER_95_37 ();
 DECAPx10_ASAP7_75t_R FILLER_95_47 ();
 DECAPx1_ASAP7_75t_R FILLER_95_69 ();
 DECAPx1_ASAP7_75t_R FILLER_95_99 ();
 FILLER_ASAP7_75t_R FILLER_95_111 ();
 DECAPx1_ASAP7_75t_R FILLER_95_119 ();
 DECAPx2_ASAP7_75t_R FILLER_95_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_139 ();
 DECAPx2_ASAP7_75t_R FILLER_95_146 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_95_152 ();
 DECAPx6_ASAP7_75t_R FILLER_95_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_172 ();
 FILLER_ASAP7_75t_R FILLER_95_179 ();
 DECAPx1_ASAP7_75t_R FILLER_95_184 ();
 DECAPx2_ASAP7_75t_R FILLER_95_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_220 ();
 DECAPx1_ASAP7_75t_R FILLER_95_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_231 ();
 DECAPx10_ASAP7_75t_R FILLER_95_235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_95_263 ();
 DECAPx2_ASAP7_75t_R FILLER_95_269 ();
 DECAPx6_ASAP7_75t_R FILLER_95_301 ();
 DECAPx2_ASAP7_75t_R FILLER_95_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_321 ();
 DECAPx4_ASAP7_75t_R FILLER_95_330 ();
 FILLER_ASAP7_75t_R FILLER_95_340 ();
 DECAPx2_ASAP7_75t_R FILLER_95_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_354 ();
 DECAPx4_ASAP7_75t_R FILLER_95_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_368 ();
 DECAPx1_ASAP7_75t_R FILLER_95_375 ();
 FILLER_ASAP7_75t_R FILLER_95_385 ();
 FILLER_ASAP7_75t_R FILLER_95_390 ();
 DECAPx4_ASAP7_75t_R FILLER_95_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_408 ();
 DECAPx2_ASAP7_75t_R FILLER_95_435 ();
 DECAPx1_ASAP7_75t_R FILLER_95_447 ();
 FILLER_ASAP7_75t_R FILLER_95_477 ();
 DECAPx2_ASAP7_75t_R FILLER_95_485 ();
 DECAPx2_ASAP7_75t_R FILLER_95_517 ();
 FILLER_ASAP7_75t_R FILLER_95_523 ();
 FILLER_ASAP7_75t_R FILLER_95_531 ();
 DECAPx2_ASAP7_75t_R FILLER_95_539 ();
 FILLER_ASAP7_75t_R FILLER_95_545 ();
 DECAPx2_ASAP7_75t_R FILLER_95_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_559 ();
 FILLER_ASAP7_75t_R FILLER_95_563 ();
 DECAPx2_ASAP7_75t_R FILLER_95_571 ();
 DECAPx10_ASAP7_75t_R FILLER_95_580 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_95_602 ();
 DECAPx1_ASAP7_75t_R FILLER_95_612 ();
 DECAPx4_ASAP7_75t_R FILLER_95_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_629 ();
 DECAPx2_ASAP7_75t_R FILLER_95_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_643 ();
 DECAPx10_ASAP7_75t_R FILLER_95_655 ();
 DECAPx10_ASAP7_75t_R FILLER_95_677 ();
 DECAPx2_ASAP7_75t_R FILLER_95_699 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_95_705 ();
 DECAPx10_ASAP7_75t_R FILLER_95_716 ();
 DECAPx4_ASAP7_75t_R FILLER_95_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_748 ();
 DECAPx2_ASAP7_75t_R FILLER_95_759 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_95_765 ();
 FILLER_ASAP7_75t_R FILLER_95_778 ();
 DECAPx6_ASAP7_75t_R FILLER_95_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_800 ();
 FILLER_ASAP7_75t_R FILLER_95_808 ();
 FILLER_ASAP7_75t_R FILLER_95_820 ();
 DECAPx10_ASAP7_75t_R FILLER_95_829 ();
 DECAPx1_ASAP7_75t_R FILLER_95_851 ();
 DECAPx10_ASAP7_75t_R FILLER_95_869 ();
 DECAPx1_ASAP7_75t_R FILLER_95_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_895 ();
 DECAPx1_ASAP7_75t_R FILLER_95_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_906 ();
 DECAPx4_ASAP7_75t_R FILLER_95_913 ();
 FILLER_ASAP7_75t_R FILLER_95_923 ();
 DECAPx1_ASAP7_75t_R FILLER_95_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_931 ();
 DECAPx10_ASAP7_75t_R FILLER_95_938 ();
 DECAPx4_ASAP7_75t_R FILLER_95_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_970 ();
 DECAPx1_ASAP7_75t_R FILLER_95_974 ();
 FILLER_ASAP7_75t_R FILLER_95_984 ();
 DECAPx10_ASAP7_75t_R FILLER_95_996 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1018 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_95_1024 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1040 ();
 FILLER_ASAP7_75t_R FILLER_95_1044 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1090 ();
 FILLER_ASAP7_75t_R FILLER_95_1094 ();
 DECAPx4_ASAP7_75t_R FILLER_95_1110 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_95_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1130 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_1151 ();
 DECAPx4_ASAP7_75t_R FILLER_95_1158 ();
 FILLER_ASAP7_75t_R FILLER_95_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1177 ();
 DECAPx6_ASAP7_75t_R FILLER_95_1193 ();
 FILLER_ASAP7_75t_R FILLER_95_1233 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1245 ();
 DECAPx2_ASAP7_75t_R FILLER_95_1255 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_95_1261 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_95_1300 ();
 DECAPx1_ASAP7_75t_R FILLER_95_1322 ();
 FILLER_ASAP7_75t_R FILLER_95_1331 ();
 FILLER_ASAP7_75t_R FILLER_95_1338 ();
 FILLER_ASAP7_75t_R FILLER_95_1345 ();
 FILLER_ASAP7_75t_R FILLER_95_1352 ();
 FILLER_ASAP7_75t_R FILLER_95_1359 ();
 FILLER_ASAP7_75t_R FILLER_95_1366 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_95_1374 ();
 DECAPx4_ASAP7_75t_R FILLER_96_2 ();
 FILLER_ASAP7_75t_R FILLER_96_12 ();
 FILLER_ASAP7_75t_R FILLER_96_20 ();
 DECAPx4_ASAP7_75t_R FILLER_96_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_35 ();
 FILLER_ASAP7_75t_R FILLER_96_42 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_50 ();
 FILLER_ASAP7_75t_R FILLER_96_59 ();
 FILLER_ASAP7_75t_R FILLER_96_67 ();
 DECAPx1_ASAP7_75t_R FILLER_96_75 ();
 FILLER_ASAP7_75t_R FILLER_96_85 ();
 DECAPx2_ASAP7_75t_R FILLER_96_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_96 ();
 FILLER_ASAP7_75t_R FILLER_96_103 ();
 DECAPx6_ASAP7_75t_R FILLER_96_113 ();
 FILLER_ASAP7_75t_R FILLER_96_127 ();
 DECAPx10_ASAP7_75t_R FILLER_96_137 ();
 DECAPx10_ASAP7_75t_R FILLER_96_159 ();
 DECAPx4_ASAP7_75t_R FILLER_96_181 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_191 ();
 FILLER_ASAP7_75t_R FILLER_96_200 ();
 DECAPx2_ASAP7_75t_R FILLER_96_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_211 ();
 DECAPx2_ASAP7_75t_R FILLER_96_224 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_230 ();
 DECAPx1_ASAP7_75t_R FILLER_96_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_243 ();
 DECAPx4_ASAP7_75t_R FILLER_96_270 ();
 FILLER_ASAP7_75t_R FILLER_96_302 ();
 DECAPx2_ASAP7_75t_R FILLER_96_307 ();
 DECAPx4_ASAP7_75t_R FILLER_96_323 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_333 ();
 DECAPx1_ASAP7_75t_R FILLER_96_342 ();
 DECAPx2_ASAP7_75t_R FILLER_96_352 ();
 DECAPx4_ASAP7_75t_R FILLER_96_384 ();
 DECAPx6_ASAP7_75t_R FILLER_96_400 ();
 DECAPx1_ASAP7_75t_R FILLER_96_420 ();
 FILLER_ASAP7_75t_R FILLER_96_430 ();
 DECAPx6_ASAP7_75t_R FILLER_96_435 ();
 DECAPx1_ASAP7_75t_R FILLER_96_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_453 ();
 FILLER_ASAP7_75t_R FILLER_96_460 ();
 FILLER_ASAP7_75t_R FILLER_96_464 ();
 DECAPx10_ASAP7_75t_R FILLER_96_469 ();
 FILLER_ASAP7_75t_R FILLER_96_491 ();
 DECAPx1_ASAP7_75t_R FILLER_96_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_503 ();
 FILLER_ASAP7_75t_R FILLER_96_507 ();
 DECAPx4_ASAP7_75t_R FILLER_96_515 ();
 DECAPx4_ASAP7_75t_R FILLER_96_551 ();
 FILLER_ASAP7_75t_R FILLER_96_561 ();
 DECAPx2_ASAP7_75t_R FILLER_96_589 ();
 FILLER_ASAP7_75t_R FILLER_96_602 ();
 DECAPx4_ASAP7_75t_R FILLER_96_610 ();
 FILLER_ASAP7_75t_R FILLER_96_620 ();
 DECAPx10_ASAP7_75t_R FILLER_96_632 ();
 DECAPx6_ASAP7_75t_R FILLER_96_654 ();
 DECAPx1_ASAP7_75t_R FILLER_96_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_672 ();
 FILLER_ASAP7_75t_R FILLER_96_682 ();
 DECAPx10_ASAP7_75t_R FILLER_96_695 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_717 ();
 FILLER_ASAP7_75t_R FILLER_96_732 ();
 DECAPx2_ASAP7_75t_R FILLER_96_740 ();
 FILLER_ASAP7_75t_R FILLER_96_746 ();
 DECAPx6_ASAP7_75t_R FILLER_96_754 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_768 ();
 DECAPx2_ASAP7_75t_R FILLER_96_778 ();
 DECAPx2_ASAP7_75t_R FILLER_96_794 ();
 DECAPx10_ASAP7_75t_R FILLER_96_806 ();
 DECAPx2_ASAP7_75t_R FILLER_96_835 ();
 DECAPx2_ASAP7_75t_R FILLER_96_849 ();
 FILLER_ASAP7_75t_R FILLER_96_875 ();
 DECAPx4_ASAP7_75t_R FILLER_96_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_893 ();
 DECAPx2_ASAP7_75t_R FILLER_96_900 ();
 FILLER_ASAP7_75t_R FILLER_96_906 ();
 FILLER_ASAP7_75t_R FILLER_96_930 ();
 FILLER_ASAP7_75t_R FILLER_96_938 ();
 FILLER_ASAP7_75t_R FILLER_96_946 ();
 DECAPx10_ASAP7_75t_R FILLER_96_954 ();
 DECAPx2_ASAP7_75t_R FILLER_96_976 ();
 FILLER_ASAP7_75t_R FILLER_96_982 ();
 DECAPx4_ASAP7_75t_R FILLER_96_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1008 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_1014 ();
 FILLER_ASAP7_75t_R FILLER_96_1023 ();
 FILLER_ASAP7_75t_R FILLER_96_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_96_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1045 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1052 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1064 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1086 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1114 ();
 FILLER_ASAP7_75t_R FILLER_96_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1128 ();
 FILLER_ASAP7_75t_R FILLER_96_1134 ();
 FILLER_ASAP7_75t_R FILLER_96_1139 ();
 FILLER_ASAP7_75t_R FILLER_96_1167 ();
 FILLER_ASAP7_75t_R FILLER_96_1195 ();
 DECAPx1_ASAP7_75t_R FILLER_96_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_96_1220 ();
 DECAPx4_ASAP7_75t_R FILLER_96_1242 ();
 FILLER_ASAP7_75t_R FILLER_96_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_96_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1275 ();
 FILLER_ASAP7_75t_R FILLER_96_1282 ();
 DECAPx6_ASAP7_75t_R FILLER_96_1287 ();
 DECAPx2_ASAP7_75t_R FILLER_96_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_1307 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_1318 ();
 FILLER_ASAP7_75t_R FILLER_96_1326 ();
 DECAPx1_ASAP7_75t_R FILLER_96_1335 ();
 FILLER_ASAP7_75t_R FILLER_96_1351 ();
 FILLER_ASAP7_75t_R FILLER_96_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_97_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_16 ();
 DECAPx6_ASAP7_75t_R FILLER_97_25 ();
 DECAPx2_ASAP7_75t_R FILLER_97_39 ();
 FILLER_ASAP7_75t_R FILLER_97_53 ();
 DECAPx2_ASAP7_75t_R FILLER_97_63 ();
 DECAPx6_ASAP7_75t_R FILLER_97_80 ();
 DECAPx2_ASAP7_75t_R FILLER_97_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_100 ();
 DECAPx6_ASAP7_75t_R FILLER_97_107 ();
 DECAPx1_ASAP7_75t_R FILLER_97_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_125 ();
 FILLER_ASAP7_75t_R FILLER_97_129 ();
 FILLER_ASAP7_75t_R FILLER_97_137 ();
 DECAPx6_ASAP7_75t_R FILLER_97_145 ();
 FILLER_ASAP7_75t_R FILLER_97_159 ();
 DECAPx10_ASAP7_75t_R FILLER_97_167 ();
 DECAPx1_ASAP7_75t_R FILLER_97_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_193 ();
 DECAPx2_ASAP7_75t_R FILLER_97_200 ();
 DECAPx6_ASAP7_75t_R FILLER_97_209 ();
 FILLER_ASAP7_75t_R FILLER_97_223 ();
 FILLER_ASAP7_75t_R FILLER_97_251 ();
 FILLER_ASAP7_75t_R FILLER_97_259 ();
 DECAPx6_ASAP7_75t_R FILLER_97_264 ();
 DECAPx1_ASAP7_75t_R FILLER_97_278 ();
 FILLER_ASAP7_75t_R FILLER_97_288 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_293 ();
 FILLER_ASAP7_75t_R FILLER_97_303 ();
 DECAPx4_ASAP7_75t_R FILLER_97_320 ();
 FILLER_ASAP7_75t_R FILLER_97_330 ();
 DECAPx1_ASAP7_75t_R FILLER_97_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_362 ();
 DECAPx1_ASAP7_75t_R FILLER_97_369 ();
 DECAPx6_ASAP7_75t_R FILLER_97_376 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_390 ();
 DECAPx6_ASAP7_75t_R FILLER_97_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_425 ();
 DECAPx2_ASAP7_75t_R FILLER_97_436 ();
 FILLER_ASAP7_75t_R FILLER_97_442 ();
 DECAPx10_ASAP7_75t_R FILLER_97_450 ();
 FILLER_ASAP7_75t_R FILLER_97_472 ();
 DECAPx1_ASAP7_75t_R FILLER_97_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_484 ();
 DECAPx2_ASAP7_75t_R FILLER_97_491 ();
 DECAPx2_ASAP7_75t_R FILLER_97_510 ();
 FILLER_ASAP7_75t_R FILLER_97_538 ();
 DECAPx6_ASAP7_75t_R FILLER_97_543 ();
 FILLER_ASAP7_75t_R FILLER_97_557 ();
 FILLER_ASAP7_75t_R FILLER_97_562 ();
 DECAPx10_ASAP7_75t_R FILLER_97_570 ();
 DECAPx6_ASAP7_75t_R FILLER_97_618 ();
 FILLER_ASAP7_75t_R FILLER_97_638 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_646 ();
 DECAPx2_ASAP7_75t_R FILLER_97_657 ();
 FILLER_ASAP7_75t_R FILLER_97_663 ();
 FILLER_ASAP7_75t_R FILLER_97_671 ();
 FILLER_ASAP7_75t_R FILLER_97_679 ();
 FILLER_ASAP7_75t_R FILLER_97_689 ();
 DECAPx1_ASAP7_75t_R FILLER_97_701 ();
 DECAPx1_ASAP7_75t_R FILLER_97_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_720 ();
 FILLER_ASAP7_75t_R FILLER_97_737 ();
 FILLER_ASAP7_75t_R FILLER_97_753 ();
 DECAPx2_ASAP7_75t_R FILLER_97_764 ();
 FILLER_ASAP7_75t_R FILLER_97_770 ();
 DECAPx2_ASAP7_75t_R FILLER_97_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_784 ();
 FILLER_ASAP7_75t_R FILLER_97_795 ();
 FILLER_ASAP7_75t_R FILLER_97_807 ();
 DECAPx2_ASAP7_75t_R FILLER_97_819 ();
 FILLER_ASAP7_75t_R FILLER_97_825 ();
 FILLER_ASAP7_75t_R FILLER_97_835 ();
 FILLER_ASAP7_75t_R FILLER_97_845 ();
 FILLER_ASAP7_75t_R FILLER_97_867 ();
 FILLER_ASAP7_75t_R FILLER_97_889 ();
 FILLER_ASAP7_75t_R FILLER_97_903 ();
 DECAPx2_ASAP7_75t_R FILLER_97_917 ();
 FILLER_ASAP7_75t_R FILLER_97_923 ();
 FILLER_ASAP7_75t_R FILLER_97_927 ();
 DECAPx2_ASAP7_75t_R FILLER_97_935 ();
 FILLER_ASAP7_75t_R FILLER_97_941 ();
 FILLER_ASAP7_75t_R FILLER_97_955 ();
 FILLER_ASAP7_75t_R FILLER_97_969 ();
 DECAPx2_ASAP7_75t_R FILLER_97_979 ();
 FILLER_ASAP7_75t_R FILLER_97_985 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_994 ();
 FILLER_ASAP7_75t_R FILLER_97_1003 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1013 ();
 FILLER_ASAP7_75t_R FILLER_97_1025 ();
 DECAPx6_ASAP7_75t_R FILLER_97_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1051 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1104 ();
 DECAPx4_ASAP7_75t_R FILLER_97_1134 ();
 FILLER_ASAP7_75t_R FILLER_97_1144 ();
 FILLER_ASAP7_75t_R FILLER_97_1153 ();
 FILLER_ASAP7_75t_R FILLER_97_1161 ();
 DECAPx4_ASAP7_75t_R FILLER_97_1166 ();
 FILLER_ASAP7_75t_R FILLER_97_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_97_1187 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1220 ();
 FILLER_ASAP7_75t_R FILLER_97_1232 ();
 DECAPx2_ASAP7_75t_R FILLER_97_1237 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_1243 ();
 FILLER_ASAP7_75t_R FILLER_97_1249 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_1257 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_1267 ();
 DECAPx6_ASAP7_75t_R FILLER_97_1276 ();
 DECAPx1_ASAP7_75t_R FILLER_97_1290 ();
 DECAPx4_ASAP7_75t_R FILLER_97_1297 ();
 FILLER_ASAP7_75t_R FILLER_97_1310 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_1318 ();
 FILLER_ASAP7_75t_R FILLER_97_1347 ();
 FILLER_ASAP7_75t_R FILLER_97_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_98_2 ();
 FILLER_ASAP7_75t_R FILLER_98_34 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_39 ();
 FILLER_ASAP7_75t_R FILLER_98_48 ();
 FILLER_ASAP7_75t_R FILLER_98_56 ();
 DECAPx10_ASAP7_75t_R FILLER_98_64 ();
 DECAPx2_ASAP7_75t_R FILLER_98_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_92 ();
 DECAPx6_ASAP7_75t_R FILLER_98_99 ();
 DECAPx1_ASAP7_75t_R FILLER_98_113 ();
 DECAPx4_ASAP7_75t_R FILLER_98_123 ();
 FILLER_ASAP7_75t_R FILLER_98_139 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_151 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_180 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_189 ();
 DECAPx2_ASAP7_75t_R FILLER_98_218 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_224 ();
 DECAPx2_ASAP7_75t_R FILLER_98_233 ();
 FILLER_ASAP7_75t_R FILLER_98_242 ();
 DECAPx10_ASAP7_75t_R FILLER_98_247 ();
 FILLER_ASAP7_75t_R FILLER_98_275 ();
 DECAPx2_ASAP7_75t_R FILLER_98_283 ();
 FILLER_ASAP7_75t_R FILLER_98_295 ();
 DECAPx2_ASAP7_75t_R FILLER_98_305 ();
 DECAPx10_ASAP7_75t_R FILLER_98_317 ();
 DECAPx2_ASAP7_75t_R FILLER_98_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_345 ();
 DECAPx10_ASAP7_75t_R FILLER_98_349 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_371 ();
 DECAPx2_ASAP7_75t_R FILLER_98_380 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_386 ();
 FILLER_ASAP7_75t_R FILLER_98_395 ();
 FILLER_ASAP7_75t_R FILLER_98_405 ();
 FILLER_ASAP7_75t_R FILLER_98_413 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_421 ();
 DECAPx1_ASAP7_75t_R FILLER_98_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_431 ();
 DECAPx1_ASAP7_75t_R FILLER_98_458 ();
 DECAPx1_ASAP7_75t_R FILLER_98_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_468 ();
 DECAPx2_ASAP7_75t_R FILLER_98_495 ();
 FILLER_ASAP7_75t_R FILLER_98_501 ();
 FILLER_ASAP7_75t_R FILLER_98_529 ();
 FILLER_ASAP7_75t_R FILLER_98_537 ();
 FILLER_ASAP7_75t_R FILLER_98_545 ();
 DECAPx1_ASAP7_75t_R FILLER_98_553 ();
 DECAPx4_ASAP7_75t_R FILLER_98_565 ();
 FILLER_ASAP7_75t_R FILLER_98_575 ();
 DECAPx10_ASAP7_75t_R FILLER_98_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_605 ();
 DECAPx6_ASAP7_75t_R FILLER_98_609 ();
 FILLER_ASAP7_75t_R FILLER_98_629 ();
 DECAPx2_ASAP7_75t_R FILLER_98_637 ();
 FILLER_ASAP7_75t_R FILLER_98_643 ();
 FILLER_ASAP7_75t_R FILLER_98_651 ();
 FILLER_ASAP7_75t_R FILLER_98_659 ();
 DECAPx6_ASAP7_75t_R FILLER_98_667 ();
 DECAPx2_ASAP7_75t_R FILLER_98_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_687 ();
 DECAPx4_ASAP7_75t_R FILLER_98_698 ();
 DECAPx6_ASAP7_75t_R FILLER_98_718 ();
 DECAPx1_ASAP7_75t_R FILLER_98_732 ();
 DECAPx6_ASAP7_75t_R FILLER_98_742 ();
 DECAPx2_ASAP7_75t_R FILLER_98_756 ();
 DECAPx4_ASAP7_75t_R FILLER_98_772 ();
 FILLER_ASAP7_75t_R FILLER_98_782 ();
 DECAPx1_ASAP7_75t_R FILLER_98_793 ();
 DECAPx4_ASAP7_75t_R FILLER_98_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_815 ();
 FILLER_ASAP7_75t_R FILLER_98_822 ();
 DECAPx2_ASAP7_75t_R FILLER_98_832 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_838 ();
 FILLER_ASAP7_75t_R FILLER_98_848 ();
 DECAPx2_ASAP7_75t_R FILLER_98_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_863 ();
 DECAPx2_ASAP7_75t_R FILLER_98_874 ();
 FILLER_ASAP7_75t_R FILLER_98_880 ();
 DECAPx2_ASAP7_75t_R FILLER_98_902 ();
 FILLER_ASAP7_75t_R FILLER_98_915 ();
 FILLER_ASAP7_75t_R FILLER_98_923 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_931 ();
 FILLER_ASAP7_75t_R FILLER_98_941 ();
 FILLER_ASAP7_75t_R FILLER_98_949 ();
 DECAPx2_ASAP7_75t_R FILLER_98_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_963 ();
 FILLER_ASAP7_75t_R FILLER_98_970 ();
 DECAPx2_ASAP7_75t_R FILLER_98_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_988 ();
 DECAPx4_ASAP7_75t_R FILLER_98_995 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_98_1015 ();
 FILLER_ASAP7_75t_R FILLER_98_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1038 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_1044 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1056 ();
 FILLER_ASAP7_75t_R FILLER_98_1086 ();
 FILLER_ASAP7_75t_R FILLER_98_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_1109 ();
 FILLER_ASAP7_75t_R FILLER_98_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_98_1147 ();
 FILLER_ASAP7_75t_R FILLER_98_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1180 ();
 FILLER_ASAP7_75t_R FILLER_98_1193 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_98_1207 ();
 FILLER_ASAP7_75t_R FILLER_98_1239 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1244 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_1257 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1267 ();
 DECAPx4_ASAP7_75t_R FILLER_98_1280 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_1290 ();
 FILLER_ASAP7_75t_R FILLER_98_1299 ();
 DECAPx1_ASAP7_75t_R FILLER_98_1307 ();
 FILLER_ASAP7_75t_R FILLER_98_1318 ();
 FILLER_ASAP7_75t_R FILLER_98_1326 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_1331 ();
 FILLER_ASAP7_75t_R FILLER_98_1340 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_1345 ();
 FILLER_ASAP7_75t_R FILLER_98_1353 ();
 FILLER_ASAP7_75t_R FILLER_98_1362 ();
 FILLER_ASAP7_75t_R FILLER_98_1370 ();
 FILLER_ASAP7_75t_R FILLER_98_1375 ();
 DECAPx4_ASAP7_75t_R FILLER_99_2 ();
 DECAPx1_ASAP7_75t_R FILLER_99_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_22 ();
 DECAPx2_ASAP7_75t_R FILLER_99_26 ();
 DECAPx10_ASAP7_75t_R FILLER_99_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_80 ();
 FILLER_ASAP7_75t_R FILLER_99_107 ();
 DECAPx6_ASAP7_75t_R FILLER_99_135 ();
 DECAPx2_ASAP7_75t_R FILLER_99_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_155 ();
 DECAPx2_ASAP7_75t_R FILLER_99_162 ();
 DECAPx2_ASAP7_75t_R FILLER_99_171 ();
 DECAPx1_ASAP7_75t_R FILLER_99_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_207 ();
 FILLER_ASAP7_75t_R FILLER_99_214 ();
 FILLER_ASAP7_75t_R FILLER_99_224 ();
 DECAPx4_ASAP7_75t_R FILLER_99_229 ();
 FILLER_ASAP7_75t_R FILLER_99_239 ();
 DECAPx4_ASAP7_75t_R FILLER_99_247 ();
 FILLER_ASAP7_75t_R FILLER_99_263 ();
 DECAPx1_ASAP7_75t_R FILLER_99_291 ();
 DECAPx6_ASAP7_75t_R FILLER_99_301 ();
 FILLER_ASAP7_75t_R FILLER_99_315 ();
 DECAPx6_ASAP7_75t_R FILLER_99_320 ();
 FILLER_ASAP7_75t_R FILLER_99_334 ();
 FILLER_ASAP7_75t_R FILLER_99_342 ();
 DECAPx2_ASAP7_75t_R FILLER_99_347 ();
 DECAPx1_ASAP7_75t_R FILLER_99_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_363 ();
 DECAPx1_ASAP7_75t_R FILLER_99_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_394 ();
 DECAPx2_ASAP7_75t_R FILLER_99_403 ();
 FILLER_ASAP7_75t_R FILLER_99_435 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_443 ();
 DECAPx1_ASAP7_75t_R FILLER_99_449 ();
 FILLER_ASAP7_75t_R FILLER_99_456 ();
 DECAPx1_ASAP7_75t_R FILLER_99_466 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_480 ();
 DECAPx2_ASAP7_75t_R FILLER_99_486 ();
 FILLER_ASAP7_75t_R FILLER_99_495 ();
 FILLER_ASAP7_75t_R FILLER_99_519 ();
 FILLER_ASAP7_75t_R FILLER_99_527 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_537 ();
 FILLER_ASAP7_75t_R FILLER_99_548 ();
 FILLER_ASAP7_75t_R FILLER_99_556 ();
 DECAPx2_ASAP7_75t_R FILLER_99_566 ();
 FILLER_ASAP7_75t_R FILLER_99_572 ();
 DECAPx1_ASAP7_75t_R FILLER_99_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_604 ();
 FILLER_ASAP7_75t_R FILLER_99_631 ();
 FILLER_ASAP7_75t_R FILLER_99_641 ();
 DECAPx4_ASAP7_75t_R FILLER_99_646 ();
 DECAPx1_ASAP7_75t_R FILLER_99_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_666 ();
 DECAPx2_ASAP7_75t_R FILLER_99_673 ();
 FILLER_ASAP7_75t_R FILLER_99_679 ();
 DECAPx1_ASAP7_75t_R FILLER_99_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_691 ();
 FILLER_ASAP7_75t_R FILLER_99_698 ();
 FILLER_ASAP7_75t_R FILLER_99_706 ();
 DECAPx10_ASAP7_75t_R FILLER_99_718 ();
 DECAPx2_ASAP7_75t_R FILLER_99_740 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_746 ();
 DECAPx4_ASAP7_75t_R FILLER_99_755 ();
 FILLER_ASAP7_75t_R FILLER_99_772 ();
 DECAPx6_ASAP7_75t_R FILLER_99_780 ();
 DECAPx1_ASAP7_75t_R FILLER_99_794 ();
 DECAPx6_ASAP7_75t_R FILLER_99_806 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_820 ();
 DECAPx10_ASAP7_75t_R FILLER_99_829 ();
 DECAPx10_ASAP7_75t_R FILLER_99_851 ();
 FILLER_ASAP7_75t_R FILLER_99_879 ();
 FILLER_ASAP7_75t_R FILLER_99_888 ();
 FILLER_ASAP7_75t_R FILLER_99_910 ();
 DECAPx2_ASAP7_75t_R FILLER_99_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_924 ();
 DECAPx10_ASAP7_75t_R FILLER_99_927 ();
 DECAPx6_ASAP7_75t_R FILLER_99_949 ();
 DECAPx1_ASAP7_75t_R FILLER_99_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_967 ();
 DECAPx1_ASAP7_75t_R FILLER_99_974 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_986 ();
 FILLER_ASAP7_75t_R FILLER_99_999 ();
 FILLER_ASAP7_75t_R FILLER_99_1013 ();
 FILLER_ASAP7_75t_R FILLER_99_1023 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_1033 ();
 FILLER_ASAP7_75t_R FILLER_99_1046 ();
 FILLER_ASAP7_75t_R FILLER_99_1057 ();
 FILLER_ASAP7_75t_R FILLER_99_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_99_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1080 ();
 FILLER_ASAP7_75t_R FILLER_99_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_99_1096 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_1106 ();
 DECAPx4_ASAP7_75t_R FILLER_99_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1126 ();
 FILLER_ASAP7_75t_R FILLER_99_1137 ();
 DECAPx1_ASAP7_75t_R FILLER_99_1145 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_99_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1212 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_1220 ();
 DECAPx1_ASAP7_75t_R FILLER_99_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1246 ();
 FILLER_ASAP7_75t_R FILLER_99_1252 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_1269 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1279 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_1285 ();
 FILLER_ASAP7_75t_R FILLER_99_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_99_1302 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_1308 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_1337 ();
 FILLER_ASAP7_75t_R FILLER_99_1345 ();
 FILLER_ASAP7_75t_R FILLER_99_1352 ();
 FILLER_ASAP7_75t_R FILLER_99_1361 ();
 FILLER_ASAP7_75t_R FILLER_99_1368 ();
 FILLER_ASAP7_75t_R FILLER_99_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_100_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_8 ();
 DECAPx6_ASAP7_75t_R FILLER_100_15 ();
 DECAPx2_ASAP7_75t_R FILLER_100_29 ();
 DECAPx1_ASAP7_75t_R FILLER_100_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_45 ();
 DECAPx10_ASAP7_75t_R FILLER_100_49 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_71 ();
 DECAPx2_ASAP7_75t_R FILLER_100_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_86 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_93 ();
 DECAPx4_ASAP7_75t_R FILLER_100_99 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_109 ();
 DECAPx1_ASAP7_75t_R FILLER_100_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_122 ();
 DECAPx2_ASAP7_75t_R FILLER_100_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_132 ();
 DECAPx6_ASAP7_75t_R FILLER_100_139 ();
 DECAPx2_ASAP7_75t_R FILLER_100_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_159 ();
 FILLER_ASAP7_75t_R FILLER_100_166 ();
 DECAPx2_ASAP7_75t_R FILLER_100_171 ();
 FILLER_ASAP7_75t_R FILLER_100_177 ();
 DECAPx2_ASAP7_75t_R FILLER_100_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_191 ();
 DECAPx1_ASAP7_75t_R FILLER_100_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_199 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_206 ();
 FILLER_ASAP7_75t_R FILLER_100_215 ();
 DECAPx1_ASAP7_75t_R FILLER_100_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_229 ();
 FILLER_ASAP7_75t_R FILLER_100_236 ();
 DECAPx2_ASAP7_75t_R FILLER_100_246 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_252 ();
 FILLER_ASAP7_75t_R FILLER_100_281 ();
 DECAPx10_ASAP7_75t_R FILLER_100_286 ();
 DECAPx2_ASAP7_75t_R FILLER_100_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_314 ();
 FILLER_ASAP7_75t_R FILLER_100_321 ();
 FILLER_ASAP7_75t_R FILLER_100_326 ();
 FILLER_ASAP7_75t_R FILLER_100_354 ();
 FILLER_ASAP7_75t_R FILLER_100_362 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_367 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_376 ();
 DECAPx2_ASAP7_75t_R FILLER_100_382 ();
 FILLER_ASAP7_75t_R FILLER_100_388 ();
 DECAPx6_ASAP7_75t_R FILLER_100_396 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_410 ();
 FILLER_ASAP7_75t_R FILLER_100_419 ();
 DECAPx10_ASAP7_75t_R FILLER_100_424 ();
 DECAPx2_ASAP7_75t_R FILLER_100_446 ();
 FILLER_ASAP7_75t_R FILLER_100_452 ();
 FILLER_ASAP7_75t_R FILLER_100_460 ();
 DECAPx2_ASAP7_75t_R FILLER_100_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_470 ();
 DECAPx6_ASAP7_75t_R FILLER_100_483 ();
 FILLER_ASAP7_75t_R FILLER_100_497 ();
 DECAPx4_ASAP7_75t_R FILLER_100_505 ();
 FILLER_ASAP7_75t_R FILLER_100_515 ();
 DECAPx2_ASAP7_75t_R FILLER_100_520 ();
 FILLER_ASAP7_75t_R FILLER_100_529 ();
 DECAPx10_ASAP7_75t_R FILLER_100_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_559 ();
 DECAPx2_ASAP7_75t_R FILLER_100_566 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_572 ();
 DECAPx2_ASAP7_75t_R FILLER_100_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_587 ();
 DECAPx6_ASAP7_75t_R FILLER_100_591 ();
 DECAPx2_ASAP7_75t_R FILLER_100_605 ();
 FILLER_ASAP7_75t_R FILLER_100_617 ();
 DECAPx10_ASAP7_75t_R FILLER_100_622 ();
 DECAPx10_ASAP7_75t_R FILLER_100_644 ();
 DECAPx6_ASAP7_75t_R FILLER_100_666 ();
 DECAPx2_ASAP7_75t_R FILLER_100_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_686 ();
 FILLER_ASAP7_75t_R FILLER_100_697 ();
 DECAPx1_ASAP7_75t_R FILLER_100_705 ();
 DECAPx4_ASAP7_75t_R FILLER_100_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_725 ();
 DECAPx2_ASAP7_75t_R FILLER_100_729 ();
 DECAPx4_ASAP7_75t_R FILLER_100_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_752 ();
 DECAPx2_ASAP7_75t_R FILLER_100_761 ();
 FILLER_ASAP7_75t_R FILLER_100_767 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_783 ();
 FILLER_ASAP7_75t_R FILLER_100_794 ();
 DECAPx4_ASAP7_75t_R FILLER_100_803 ();
 FILLER_ASAP7_75t_R FILLER_100_813 ();
 DECAPx1_ASAP7_75t_R FILLER_100_822 ();
 DECAPx1_ASAP7_75t_R FILLER_100_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_837 ();
 FILLER_ASAP7_75t_R FILLER_100_846 ();
 FILLER_ASAP7_75t_R FILLER_100_854 ();
 DECAPx2_ASAP7_75t_R FILLER_100_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_871 ();
 FILLER_ASAP7_75t_R FILLER_100_892 ();
 FILLER_ASAP7_75t_R FILLER_100_914 ();
 DECAPx2_ASAP7_75t_R FILLER_100_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_928 ();
 DECAPx2_ASAP7_75t_R FILLER_100_935 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_941 ();
 DECAPx4_ASAP7_75t_R FILLER_100_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_963 ();
 DECAPx2_ASAP7_75t_R FILLER_100_974 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_980 ();
 FILLER_ASAP7_75t_R FILLER_100_989 ();
 DECAPx4_ASAP7_75t_R FILLER_100_1005 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_1015 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1026 ();
 DECAPx4_ASAP7_75t_R FILLER_100_1042 ();
 FILLER_ASAP7_75t_R FILLER_100_1052 ();
 DECAPx6_ASAP7_75t_R FILLER_100_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1100 ();
 FILLER_ASAP7_75t_R FILLER_100_1132 ();
 FILLER_ASAP7_75t_R FILLER_100_1160 ();
 FILLER_ASAP7_75t_R FILLER_100_1169 ();
 FILLER_ASAP7_75t_R FILLER_100_1177 ();
 DECAPx4_ASAP7_75t_R FILLER_100_1182 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_1192 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_100_1237 ();
 DECAPx6_ASAP7_75t_R FILLER_100_1259 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1273 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1282 ();
 FILLER_ASAP7_75t_R FILLER_100_1293 ();
 DECAPx4_ASAP7_75t_R FILLER_100_1301 ();
 DECAPx1_ASAP7_75t_R FILLER_100_1317 ();
 FILLER_ASAP7_75t_R FILLER_100_1324 ();
 DECAPx2_ASAP7_75t_R FILLER_100_1329 ();
 FILLER_ASAP7_75t_R FILLER_100_1340 ();
 FILLER_ASAP7_75t_R FILLER_100_1347 ();
 FILLER_ASAP7_75t_R FILLER_100_1375 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_2 ();
 DECAPx10_ASAP7_75t_R FILLER_101_31 ();
 DECAPx4_ASAP7_75t_R FILLER_101_53 ();
 FILLER_ASAP7_75t_R FILLER_101_63 ();
 FILLER_ASAP7_75t_R FILLER_101_91 ();
 DECAPx4_ASAP7_75t_R FILLER_101_96 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_106 ();
 DECAPx2_ASAP7_75t_R FILLER_101_117 ();
 FILLER_ASAP7_75t_R FILLER_101_149 ();
 DECAPx2_ASAP7_75t_R FILLER_101_177 ();
 FILLER_ASAP7_75t_R FILLER_101_183 ();
 DECAPx10_ASAP7_75t_R FILLER_101_191 ();
 DECAPx4_ASAP7_75t_R FILLER_101_213 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_223 ();
 FILLER_ASAP7_75t_R FILLER_101_232 ();
 FILLER_ASAP7_75t_R FILLER_101_242 ();
 DECAPx2_ASAP7_75t_R FILLER_101_250 ();
 FILLER_ASAP7_75t_R FILLER_101_256 ();
 DECAPx2_ASAP7_75t_R FILLER_101_264 ();
 DECAPx6_ASAP7_75t_R FILLER_101_273 ();
 DECAPx1_ASAP7_75t_R FILLER_101_287 ();
 FILLER_ASAP7_75t_R FILLER_101_297 ();
 DECAPx2_ASAP7_75t_R FILLER_101_302 ();
 FILLER_ASAP7_75t_R FILLER_101_334 ();
 DECAPx4_ASAP7_75t_R FILLER_101_342 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_352 ();
 FILLER_ASAP7_75t_R FILLER_101_361 ();
 DECAPx6_ASAP7_75t_R FILLER_101_369 ();
 DECAPx1_ASAP7_75t_R FILLER_101_383 ();
 FILLER_ASAP7_75t_R FILLER_101_390 ();
 DECAPx10_ASAP7_75t_R FILLER_101_398 ();
 DECAPx1_ASAP7_75t_R FILLER_101_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_424 ();
 DECAPx1_ASAP7_75t_R FILLER_101_428 ();
 DECAPx1_ASAP7_75t_R FILLER_101_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_442 ();
 DECAPx2_ASAP7_75t_R FILLER_101_465 ();
 FILLER_ASAP7_75t_R FILLER_101_471 ();
 DECAPx2_ASAP7_75t_R FILLER_101_481 ();
 FILLER_ASAP7_75t_R FILLER_101_493 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_503 ();
 FILLER_ASAP7_75t_R FILLER_101_509 ();
 DECAPx2_ASAP7_75t_R FILLER_101_519 ();
 DECAPx6_ASAP7_75t_R FILLER_101_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_547 ();
 DECAPx10_ASAP7_75t_R FILLER_101_554 ();
 DECAPx10_ASAP7_75t_R FILLER_101_576 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_598 ();
 DECAPx2_ASAP7_75t_R FILLER_101_609 ();
 DECAPx2_ASAP7_75t_R FILLER_101_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_631 ();
 DECAPx1_ASAP7_75t_R FILLER_101_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_642 ();
 DECAPx2_ASAP7_75t_R FILLER_101_646 ();
 FILLER_ASAP7_75t_R FILLER_101_658 ();
 DECAPx1_ASAP7_75t_R FILLER_101_668 ();
 DECAPx4_ASAP7_75t_R FILLER_101_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_689 ();
 DECAPx2_ASAP7_75t_R FILLER_101_698 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_704 ();
 DECAPx2_ASAP7_75t_R FILLER_101_713 ();
 DECAPx2_ASAP7_75t_R FILLER_101_725 ();
 DECAPx1_ASAP7_75t_R FILLER_101_745 ();
 FILLER_ASAP7_75t_R FILLER_101_759 ();
 FILLER_ASAP7_75t_R FILLER_101_771 ();
 DECAPx2_ASAP7_75t_R FILLER_101_780 ();
 FILLER_ASAP7_75t_R FILLER_101_786 ();
 DECAPx2_ASAP7_75t_R FILLER_101_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_804 ();
 FILLER_ASAP7_75t_R FILLER_101_819 ();
 DECAPx2_ASAP7_75t_R FILLER_101_829 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_835 ();
 FILLER_ASAP7_75t_R FILLER_101_847 ();
 FILLER_ASAP7_75t_R FILLER_101_856 ();
 FILLER_ASAP7_75t_R FILLER_101_869 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_877 ();
 DECAPx1_ASAP7_75t_R FILLER_101_887 ();
 FILLER_ASAP7_75t_R FILLER_101_899 ();
 DECAPx1_ASAP7_75t_R FILLER_101_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_915 ();
 FILLER_ASAP7_75t_R FILLER_101_923 ();
 FILLER_ASAP7_75t_R FILLER_101_927 ();
 DECAPx2_ASAP7_75t_R FILLER_101_937 ();
 FILLER_ASAP7_75t_R FILLER_101_943 ();
 FILLER_ASAP7_75t_R FILLER_101_955 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_964 ();
 DECAPx10_ASAP7_75t_R FILLER_101_973 ();
 FILLER_ASAP7_75t_R FILLER_101_995 ();
 DECAPx6_ASAP7_75t_R FILLER_101_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1048 ();
 DECAPx6_ASAP7_75t_R FILLER_101_1077 ();
 FILLER_ASAP7_75t_R FILLER_101_1091 ();
 DECAPx6_ASAP7_75t_R FILLER_101_1099 ();
 FILLER_ASAP7_75t_R FILLER_101_1119 ();
 DECAPx2_ASAP7_75t_R FILLER_101_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1130 ();
 DECAPx2_ASAP7_75t_R FILLER_101_1138 ();
 DECAPx6_ASAP7_75t_R FILLER_101_1147 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_101_1189 ();
 FILLER_ASAP7_75t_R FILLER_101_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_101_1200 ();
 DECAPx1_ASAP7_75t_R FILLER_101_1222 ();
 DECAPx4_ASAP7_75t_R FILLER_101_1229 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_1239 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_1249 ();
 DECAPx6_ASAP7_75t_R FILLER_101_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_101_1276 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1282 ();
 DECAPx1_ASAP7_75t_R FILLER_101_1309 ();
 DECAPx2_ASAP7_75t_R FILLER_101_1320 ();
 FILLER_ASAP7_75t_R FILLER_101_1326 ();
 DECAPx1_ASAP7_75t_R FILLER_101_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_1340 ();
 FILLER_ASAP7_75t_R FILLER_101_1346 ();
 FILLER_ASAP7_75t_R FILLER_101_1356 ();
 DECAPx1_ASAP7_75t_R FILLER_101_1364 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_1374 ();
 DECAPx1_ASAP7_75t_R FILLER_102_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_6 ();
 DECAPx2_ASAP7_75t_R FILLER_102_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_19 ();
 DECAPx1_ASAP7_75t_R FILLER_102_23 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_33 ();
 DECAPx2_ASAP7_75t_R FILLER_102_39 ();
 FILLER_ASAP7_75t_R FILLER_102_45 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_55 ();
 DECAPx1_ASAP7_75t_R FILLER_102_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_68 ();
 DECAPx1_ASAP7_75t_R FILLER_102_75 ();
 DECAPx10_ASAP7_75t_R FILLER_102_82 ();
 DECAPx2_ASAP7_75t_R FILLER_102_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_110 ();
 DECAPx4_ASAP7_75t_R FILLER_102_119 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_135 ();
 DECAPx4_ASAP7_75t_R FILLER_102_141 ();
 FILLER_ASAP7_75t_R FILLER_102_151 ();
 DECAPx2_ASAP7_75t_R FILLER_102_159 ();
 DECAPx4_ASAP7_75t_R FILLER_102_168 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_178 ();
 DECAPx10_ASAP7_75t_R FILLER_102_207 ();
 DECAPx10_ASAP7_75t_R FILLER_102_229 ();
 DECAPx10_ASAP7_75t_R FILLER_102_251 ();
 DECAPx2_ASAP7_75t_R FILLER_102_273 ();
 FILLER_ASAP7_75t_R FILLER_102_279 ();
 DECAPx1_ASAP7_75t_R FILLER_102_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_311 ();
 FILLER_ASAP7_75t_R FILLER_102_318 ();
 DECAPx10_ASAP7_75t_R FILLER_102_342 ();
 DECAPx4_ASAP7_75t_R FILLER_102_364 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_374 ();
 FILLER_ASAP7_75t_R FILLER_102_383 ();
 DECAPx1_ASAP7_75t_R FILLER_102_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_392 ();
 FILLER_ASAP7_75t_R FILLER_102_401 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_409 ();
 FILLER_ASAP7_75t_R FILLER_102_418 ();
 FILLER_ASAP7_75t_R FILLER_102_426 ();
 FILLER_ASAP7_75t_R FILLER_102_454 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_459 ();
 FILLER_ASAP7_75t_R FILLER_102_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_473 ();
 FILLER_ASAP7_75t_R FILLER_102_502 ();
 FILLER_ASAP7_75t_R FILLER_102_512 ();
 FILLER_ASAP7_75t_R FILLER_102_536 ();
 DECAPx6_ASAP7_75t_R FILLER_102_545 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_585 ();
 FILLER_ASAP7_75t_R FILLER_102_614 ();
 DECAPx1_ASAP7_75t_R FILLER_102_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_625 ();
 DECAPx2_ASAP7_75t_R FILLER_102_635 ();
 FILLER_ASAP7_75t_R FILLER_102_647 ();
 FILLER_ASAP7_75t_R FILLER_102_655 ();
 FILLER_ASAP7_75t_R FILLER_102_664 ();
 FILLER_ASAP7_75t_R FILLER_102_674 ();
 DECAPx2_ASAP7_75t_R FILLER_102_682 ();
 DECAPx4_ASAP7_75t_R FILLER_102_699 ();
 FILLER_ASAP7_75t_R FILLER_102_715 ();
 DECAPx1_ASAP7_75t_R FILLER_102_727 ();
 DECAPx6_ASAP7_75t_R FILLER_102_737 ();
 FILLER_ASAP7_75t_R FILLER_102_751 ();
 DECAPx2_ASAP7_75t_R FILLER_102_759 ();
 FILLER_ASAP7_75t_R FILLER_102_765 ();
 DECAPx1_ASAP7_75t_R FILLER_102_774 ();
 DECAPx1_ASAP7_75t_R FILLER_102_786 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_796 ();
 DECAPx4_ASAP7_75t_R FILLER_102_805 ();
 FILLER_ASAP7_75t_R FILLER_102_815 ();
 DECAPx10_ASAP7_75t_R FILLER_102_824 ();
 DECAPx2_ASAP7_75t_R FILLER_102_846 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_852 ();
 FILLER_ASAP7_75t_R FILLER_102_861 ();
 DECAPx1_ASAP7_75t_R FILLER_102_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_873 ();
 FILLER_ASAP7_75t_R FILLER_102_880 ();
 DECAPx1_ASAP7_75t_R FILLER_102_889 ();
 DECAPx2_ASAP7_75t_R FILLER_102_901 ();
 FILLER_ASAP7_75t_R FILLER_102_914 ();
 DECAPx2_ASAP7_75t_R FILLER_102_919 ();
 FILLER_ASAP7_75t_R FILLER_102_931 ();
 FILLER_ASAP7_75t_R FILLER_102_939 ();
 DECAPx2_ASAP7_75t_R FILLER_102_947 ();
 DECAPx2_ASAP7_75t_R FILLER_102_959 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_965 ();
 DECAPx2_ASAP7_75t_R FILLER_102_988 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_994 ();
 DECAPx1_ASAP7_75t_R FILLER_102_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1009 ();
 DECAPx4_ASAP7_75t_R FILLER_102_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1028 ();
 DECAPx4_ASAP7_75t_R FILLER_102_1039 ();
 FILLER_ASAP7_75t_R FILLER_102_1049 ();
 FILLER_ASAP7_75t_R FILLER_102_1058 ();
 FILLER_ASAP7_75t_R FILLER_102_1066 ();
 FILLER_ASAP7_75t_R FILLER_102_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1148 ();
 FILLER_ASAP7_75t_R FILLER_102_1155 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1163 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_102_1187 ();
 FILLER_ASAP7_75t_R FILLER_102_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_102_1199 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1221 ();
 FILLER_ASAP7_75t_R FILLER_102_1235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_1263 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_1273 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1279 ();
 DECAPx1_ASAP7_75t_R FILLER_102_1293 ();
 DECAPx6_ASAP7_75t_R FILLER_102_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1314 ();
 FILLER_ASAP7_75t_R FILLER_102_1341 ();
 DECAPx1_ASAP7_75t_R FILLER_102_1351 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_1355 ();
 FILLER_ASAP7_75t_R FILLER_102_1361 ();
 FILLER_ASAP7_75t_R FILLER_102_1368 ();
 FILLER_ASAP7_75t_R FILLER_102_1375 ();
 DECAPx4_ASAP7_75t_R FILLER_103_2 ();
 FILLER_ASAP7_75t_R FILLER_103_12 ();
 DECAPx1_ASAP7_75t_R FILLER_103_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_44 ();
 FILLER_ASAP7_75t_R FILLER_103_53 ();
 DECAPx6_ASAP7_75t_R FILLER_103_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_75 ();
 DECAPx1_ASAP7_75t_R FILLER_103_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_86 ();
 FILLER_ASAP7_75t_R FILLER_103_93 ();
 FILLER_ASAP7_75t_R FILLER_103_103 ();
 FILLER_ASAP7_75t_R FILLER_103_111 ();
 DECAPx2_ASAP7_75t_R FILLER_103_119 ();
 FILLER_ASAP7_75t_R FILLER_103_125 ();
 DECAPx6_ASAP7_75t_R FILLER_103_133 ();
 DECAPx1_ASAP7_75t_R FILLER_103_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_151 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_155 ();
 FILLER_ASAP7_75t_R FILLER_103_164 ();
 DECAPx4_ASAP7_75t_R FILLER_103_172 ();
 DECAPx2_ASAP7_75t_R FILLER_103_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_194 ();
 DECAPx4_ASAP7_75t_R FILLER_103_198 ();
 FILLER_ASAP7_75t_R FILLER_103_208 ();
 FILLER_ASAP7_75t_R FILLER_103_220 ();
 DECAPx4_ASAP7_75t_R FILLER_103_228 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_238 ();
 DECAPx2_ASAP7_75t_R FILLER_103_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_255 ();
 FILLER_ASAP7_75t_R FILLER_103_262 ();
 DECAPx2_ASAP7_75t_R FILLER_103_267 ();
 DECAPx2_ASAP7_75t_R FILLER_103_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_285 ();
 FILLER_ASAP7_75t_R FILLER_103_292 ();
 DECAPx2_ASAP7_75t_R FILLER_103_297 ();
 FILLER_ASAP7_75t_R FILLER_103_303 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_331 ();
 FILLER_ASAP7_75t_R FILLER_103_340 ();
 DECAPx2_ASAP7_75t_R FILLER_103_345 ();
 FILLER_ASAP7_75t_R FILLER_103_351 ();
 FILLER_ASAP7_75t_R FILLER_103_361 ();
 FILLER_ASAP7_75t_R FILLER_103_369 ();
 FILLER_ASAP7_75t_R FILLER_103_397 ();
 DECAPx1_ASAP7_75t_R FILLER_103_407 ();
 FILLER_ASAP7_75t_R FILLER_103_437 ();
 DECAPx2_ASAP7_75t_R FILLER_103_445 ();
 FILLER_ASAP7_75t_R FILLER_103_457 ();
 DECAPx2_ASAP7_75t_R FILLER_103_469 ();
 FILLER_ASAP7_75t_R FILLER_103_481 ();
 FILLER_ASAP7_75t_R FILLER_103_489 ();
 DECAPx6_ASAP7_75t_R FILLER_103_494 ();
 DECAPx2_ASAP7_75t_R FILLER_103_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_514 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_522 ();
 FILLER_ASAP7_75t_R FILLER_103_551 ();
 FILLER_ASAP7_75t_R FILLER_103_556 ();
 DECAPx2_ASAP7_75t_R FILLER_103_565 ();
 FILLER_ASAP7_75t_R FILLER_103_571 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_599 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_605 ();
 DECAPx10_ASAP7_75t_R FILLER_103_612 ();
 DECAPx2_ASAP7_75t_R FILLER_103_634 ();
 DECAPx10_ASAP7_75t_R FILLER_103_648 ();
 FILLER_ASAP7_75t_R FILLER_103_678 ();
 DECAPx10_ASAP7_75t_R FILLER_103_690 ();
 DECAPx6_ASAP7_75t_R FILLER_103_712 ();
 DECAPx6_ASAP7_75t_R FILLER_103_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_749 ();
 FILLER_ASAP7_75t_R FILLER_103_756 ();
 DECAPx2_ASAP7_75t_R FILLER_103_765 ();
 FILLER_ASAP7_75t_R FILLER_103_799 ();
 DECAPx10_ASAP7_75t_R FILLER_103_807 ();
 DECAPx10_ASAP7_75t_R FILLER_103_829 ();
 DECAPx10_ASAP7_75t_R FILLER_103_851 ();
 DECAPx2_ASAP7_75t_R FILLER_103_873 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_879 ();
 DECAPx10_ASAP7_75t_R FILLER_103_890 ();
 DECAPx4_ASAP7_75t_R FILLER_103_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_922 ();
 DECAPx2_ASAP7_75t_R FILLER_103_927 ();
 FILLER_ASAP7_75t_R FILLER_103_933 ();
 DECAPx6_ASAP7_75t_R FILLER_103_943 ();
 DECAPx2_ASAP7_75t_R FILLER_103_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_963 ();
 DECAPx2_ASAP7_75t_R FILLER_103_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_977 ();
 DECAPx2_ASAP7_75t_R FILLER_103_984 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_990 ();
 FILLER_ASAP7_75t_R FILLER_103_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_103_1019 ();
 FILLER_ASAP7_75t_R FILLER_103_1041 ();
 DECAPx1_ASAP7_75t_R FILLER_103_1046 ();
 FILLER_ASAP7_75t_R FILLER_103_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_103_1084 ();
 FILLER_ASAP7_75t_R FILLER_103_1114 ();
 FILLER_ASAP7_75t_R FILLER_103_1123 ();
 DECAPx4_ASAP7_75t_R FILLER_103_1131 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_1141 ();
 DECAPx1_ASAP7_75t_R FILLER_103_1154 ();
 DECAPx4_ASAP7_75t_R FILLER_103_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1175 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1202 ();
 FILLER_ASAP7_75t_R FILLER_103_1216 ();
 FILLER_ASAP7_75t_R FILLER_103_1225 ();
 FILLER_ASAP7_75t_R FILLER_103_1233 ();
 DECAPx4_ASAP7_75t_R FILLER_103_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1248 ();
 FILLER_ASAP7_75t_R FILLER_103_1255 ();
 FILLER_ASAP7_75t_R FILLER_103_1260 ();
 DECAPx6_ASAP7_75t_R FILLER_103_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1302 ();
 DECAPx6_ASAP7_75t_R FILLER_103_1310 ();
 DECAPx1_ASAP7_75t_R FILLER_103_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_1328 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_1332 ();
 DECAPx2_ASAP7_75t_R FILLER_103_1338 ();
 FILLER_ASAP7_75t_R FILLER_103_1352 ();
 FILLER_ASAP7_75t_R FILLER_103_1361 ();
 FILLER_ASAP7_75t_R FILLER_103_1366 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_1374 ();
 DECAPx6_ASAP7_75t_R FILLER_104_2 ();
 DECAPx1_ASAP7_75t_R FILLER_104_16 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_26 ();
 DECAPx4_ASAP7_75t_R FILLER_104_32 ();
 DECAPx2_ASAP7_75t_R FILLER_104_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_54 ();
 DECAPx2_ASAP7_75t_R FILLER_104_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_67 ();
 FILLER_ASAP7_75t_R FILLER_104_94 ();
 DECAPx6_ASAP7_75t_R FILLER_104_104 ();
 DECAPx2_ASAP7_75t_R FILLER_104_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_124 ();
 FILLER_ASAP7_75t_R FILLER_104_151 ();
 FILLER_ASAP7_75t_R FILLER_104_159 ();
 DECAPx6_ASAP7_75t_R FILLER_104_169 ();
 DECAPx1_ASAP7_75t_R FILLER_104_183 ();
 DECAPx1_ASAP7_75t_R FILLER_104_193 ();
 FILLER_ASAP7_75t_R FILLER_104_203 ();
 DECAPx1_ASAP7_75t_R FILLER_104_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_215 ();
 FILLER_ASAP7_75t_R FILLER_104_219 ();
 FILLER_ASAP7_75t_R FILLER_104_229 ();
 DECAPx2_ASAP7_75t_R FILLER_104_237 ();
 FILLER_ASAP7_75t_R FILLER_104_269 ();
 DECAPx1_ASAP7_75t_R FILLER_104_297 ();
 FILLER_ASAP7_75t_R FILLER_104_304 ();
 FILLER_ASAP7_75t_R FILLER_104_313 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_322 ();
 FILLER_ASAP7_75t_R FILLER_104_351 ();
 FILLER_ASAP7_75t_R FILLER_104_361 ();
 DECAPx1_ASAP7_75t_R FILLER_104_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_373 ();
 DECAPx4_ASAP7_75t_R FILLER_104_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_390 ();
 DECAPx6_ASAP7_75t_R FILLER_104_398 ();
 DECAPx2_ASAP7_75t_R FILLER_104_412 ();
 DECAPx2_ASAP7_75t_R FILLER_104_440 ();
 DECAPx4_ASAP7_75t_R FILLER_104_452 ();
 FILLER_ASAP7_75t_R FILLER_104_464 ();
 DECAPx10_ASAP7_75t_R FILLER_104_469 ();
 DECAPx10_ASAP7_75t_R FILLER_104_491 ();
 DECAPx6_ASAP7_75t_R FILLER_104_519 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_533 ();
 FILLER_ASAP7_75t_R FILLER_104_539 ();
 FILLER_ASAP7_75t_R FILLER_104_563 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_568 ();
 FILLER_ASAP7_75t_R FILLER_104_578 ();
 DECAPx2_ASAP7_75t_R FILLER_104_586 ();
 FILLER_ASAP7_75t_R FILLER_104_595 ();
 DECAPx2_ASAP7_75t_R FILLER_104_600 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_606 ();
 DECAPx4_ASAP7_75t_R FILLER_104_615 ();
 FILLER_ASAP7_75t_R FILLER_104_631 ();
 DECAPx4_ASAP7_75t_R FILLER_104_640 ();
 DECAPx10_ASAP7_75t_R FILLER_104_656 ();
 DECAPx6_ASAP7_75t_R FILLER_104_678 ();
 DECAPx1_ASAP7_75t_R FILLER_104_692 ();
 DECAPx10_ASAP7_75t_R FILLER_104_708 ();
 DECAPx6_ASAP7_75t_R FILLER_104_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_751 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_761 ();
 FILLER_ASAP7_75t_R FILLER_104_774 ();
 FILLER_ASAP7_75t_R FILLER_104_788 ();
 DECAPx2_ASAP7_75t_R FILLER_104_796 ();
 FILLER_ASAP7_75t_R FILLER_104_802 ();
 DECAPx6_ASAP7_75t_R FILLER_104_813 ();
 DECAPx2_ASAP7_75t_R FILLER_104_834 ();
 DECAPx1_ASAP7_75t_R FILLER_104_847 ();
 FILLER_ASAP7_75t_R FILLER_104_857 ();
 DECAPx1_ASAP7_75t_R FILLER_104_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_866 ();
 FILLER_ASAP7_75t_R FILLER_104_874 ();
 DECAPx6_ASAP7_75t_R FILLER_104_883 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_897 ();
 DECAPx6_ASAP7_75t_R FILLER_104_910 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_924 ();
 FILLER_ASAP7_75t_R FILLER_104_935 ();
 DECAPx1_ASAP7_75t_R FILLER_104_946 ();
 DECAPx2_ASAP7_75t_R FILLER_104_956 ();
 DECAPx2_ASAP7_75t_R FILLER_104_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_974 ();
 DECAPx4_ASAP7_75t_R FILLER_104_984 ();
 DECAPx4_ASAP7_75t_R FILLER_104_1000 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_1010 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_1021 ();
 FILLER_ASAP7_75t_R FILLER_104_1030 ();
 DECAPx6_ASAP7_75t_R FILLER_104_1038 ();
 FILLER_ASAP7_75t_R FILLER_104_1052 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_1062 ();
 DECAPx6_ASAP7_75t_R FILLER_104_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1101 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1105 ();
 FILLER_ASAP7_75t_R FILLER_104_1135 ();
 DECAPx4_ASAP7_75t_R FILLER_104_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_1157 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_1184 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1193 ();
 FILLER_ASAP7_75t_R FILLER_104_1199 ();
 FILLER_ASAP7_75t_R FILLER_104_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_104_1237 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1259 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_1265 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_104_1280 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1294 ();
 FILLER_ASAP7_75t_R FILLER_104_1300 ();
 DECAPx2_ASAP7_75t_R FILLER_104_1309 ();
 FILLER_ASAP7_75t_R FILLER_104_1315 ();
 FILLER_ASAP7_75t_R FILLER_104_1327 ();
 DECAPx4_ASAP7_75t_R FILLER_104_1336 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_1346 ();
 FILLER_ASAP7_75t_R FILLER_104_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_105_2 ();
 DECAPx2_ASAP7_75t_R FILLER_105_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_22 ();
 DECAPx10_ASAP7_75t_R FILLER_105_29 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_51 ();
 FILLER_ASAP7_75t_R FILLER_105_60 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_68 ();
 DECAPx1_ASAP7_75t_R FILLER_105_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_81 ();
 DECAPx2_ASAP7_75t_R FILLER_105_85 ();
 DECAPx2_ASAP7_75t_R FILLER_105_97 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_103 ();
 DECAPx6_ASAP7_75t_R FILLER_105_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_127 ();
 DECAPx1_ASAP7_75t_R FILLER_105_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_138 ();
 FILLER_ASAP7_75t_R FILLER_105_142 ();
 DECAPx6_ASAP7_75t_R FILLER_105_150 ();
 DECAPx1_ASAP7_75t_R FILLER_105_164 ();
 DECAPx1_ASAP7_75t_R FILLER_105_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_180 ();
 FILLER_ASAP7_75t_R FILLER_105_207 ();
 DECAPx4_ASAP7_75t_R FILLER_105_212 ();
 FILLER_ASAP7_75t_R FILLER_105_222 ();
 DECAPx2_ASAP7_75t_R FILLER_105_230 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_236 ();
 FILLER_ASAP7_75t_R FILLER_105_245 ();
 DECAPx2_ASAP7_75t_R FILLER_105_253 ();
 FILLER_ASAP7_75t_R FILLER_105_259 ();
 DECAPx2_ASAP7_75t_R FILLER_105_264 ();
 FILLER_ASAP7_75t_R FILLER_105_270 ();
 DECAPx4_ASAP7_75t_R FILLER_105_278 ();
 DECAPx1_ASAP7_75t_R FILLER_105_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_298 ();
 FILLER_ASAP7_75t_R FILLER_105_305 ();
 FILLER_ASAP7_75t_R FILLER_105_313 ();
 FILLER_ASAP7_75t_R FILLER_105_322 ();
 FILLER_ASAP7_75t_R FILLER_105_331 ();
 FILLER_ASAP7_75t_R FILLER_105_339 ();
 DECAPx2_ASAP7_75t_R FILLER_105_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_350 ();
 FILLER_ASAP7_75t_R FILLER_105_357 ();
 DECAPx2_ASAP7_75t_R FILLER_105_365 ();
 FILLER_ASAP7_75t_R FILLER_105_371 ();
 DECAPx1_ASAP7_75t_R FILLER_105_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_383 ();
 DECAPx6_ASAP7_75t_R FILLER_105_390 ();
 DECAPx1_ASAP7_75t_R FILLER_105_404 ();
 DECAPx1_ASAP7_75t_R FILLER_105_414 ();
 DECAPx6_ASAP7_75t_R FILLER_105_421 ();
 DECAPx1_ASAP7_75t_R FILLER_105_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_439 ();
 FILLER_ASAP7_75t_R FILLER_105_466 ();
 DECAPx6_ASAP7_75t_R FILLER_105_475 ();
 DECAPx1_ASAP7_75t_R FILLER_105_489 ();
 FILLER_ASAP7_75t_R FILLER_105_499 ();
 DECAPx1_ASAP7_75t_R FILLER_105_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_511 ();
 DECAPx4_ASAP7_75t_R FILLER_105_518 ();
 FILLER_ASAP7_75t_R FILLER_105_528 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_537 ();
 DECAPx4_ASAP7_75t_R FILLER_105_546 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_556 ();
 DECAPx2_ASAP7_75t_R FILLER_105_565 ();
 FILLER_ASAP7_75t_R FILLER_105_571 ();
 DECAPx6_ASAP7_75t_R FILLER_105_576 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_590 ();
 FILLER_ASAP7_75t_R FILLER_105_619 ();
 FILLER_ASAP7_75t_R FILLER_105_628 ();
 DECAPx4_ASAP7_75t_R FILLER_105_636 ();
 FILLER_ASAP7_75t_R FILLER_105_646 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_656 ();
 FILLER_ASAP7_75t_R FILLER_105_667 ();
 DECAPx2_ASAP7_75t_R FILLER_105_676 ();
 FILLER_ASAP7_75t_R FILLER_105_694 ();
 FILLER_ASAP7_75t_R FILLER_105_703 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_711 ();
 FILLER_ASAP7_75t_R FILLER_105_726 ();
 DECAPx4_ASAP7_75t_R FILLER_105_734 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_744 ();
 DECAPx6_ASAP7_75t_R FILLER_105_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_789 ();
 DECAPx4_ASAP7_75t_R FILLER_105_800 ();
 DECAPx2_ASAP7_75t_R FILLER_105_819 ();
 DECAPx2_ASAP7_75t_R FILLER_105_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_841 ();
 FILLER_ASAP7_75t_R FILLER_105_854 ();
 DECAPx1_ASAP7_75t_R FILLER_105_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_868 ();
 DECAPx6_ASAP7_75t_R FILLER_105_877 ();
 DECAPx2_ASAP7_75t_R FILLER_105_891 ();
 FILLER_ASAP7_75t_R FILLER_105_903 ();
 DECAPx1_ASAP7_75t_R FILLER_105_913 ();
 FILLER_ASAP7_75t_R FILLER_105_923 ();
 FILLER_ASAP7_75t_R FILLER_105_927 ();
 DECAPx4_ASAP7_75t_R FILLER_105_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_947 ();
 DECAPx2_ASAP7_75t_R FILLER_105_955 ();
 FILLER_ASAP7_75t_R FILLER_105_968 ();
 DECAPx10_ASAP7_75t_R FILLER_105_985 ();
 DECAPx6_ASAP7_75t_R FILLER_105_1007 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1078 ();
 DECAPx6_ASAP7_75t_R FILLER_105_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1120 ();
 DECAPx4_ASAP7_75t_R FILLER_105_1131 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1147 ();
 DECAPx1_ASAP7_75t_R FILLER_105_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1176 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1186 ();
 FILLER_ASAP7_75t_R FILLER_105_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1225 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_105_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_1293 ();
 DECAPx4_ASAP7_75t_R FILLER_105_1320 ();
 FILLER_ASAP7_75t_R FILLER_105_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_105_1364 ();
 FILLER_ASAP7_75t_R FILLER_105_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_106_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_16 ();
 FILLER_ASAP7_75t_R FILLER_106_43 ();
 DECAPx2_ASAP7_75t_R FILLER_106_48 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_54 ();
 FILLER_ASAP7_75t_R FILLER_106_63 ();
 DECAPx2_ASAP7_75t_R FILLER_106_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_77 ();
 DECAPx6_ASAP7_75t_R FILLER_106_84 ();
 DECAPx1_ASAP7_75t_R FILLER_106_98 ();
 DECAPx1_ASAP7_75t_R FILLER_106_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_112 ();
 DECAPx1_ASAP7_75t_R FILLER_106_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_125 ();
 DECAPx2_ASAP7_75t_R FILLER_106_152 ();
 FILLER_ASAP7_75t_R FILLER_106_158 ();
 DECAPx2_ASAP7_75t_R FILLER_106_166 ();
 DECAPx1_ASAP7_75t_R FILLER_106_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_182 ();
 DECAPx2_ASAP7_75t_R FILLER_106_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_195 ();
 DECAPx10_ASAP7_75t_R FILLER_106_199 ();
 DECAPx10_ASAP7_75t_R FILLER_106_221 ();
 DECAPx6_ASAP7_75t_R FILLER_106_243 ();
 DECAPx1_ASAP7_75t_R FILLER_106_257 ();
 DECAPx6_ASAP7_75t_R FILLER_106_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_283 ();
 DECAPx1_ASAP7_75t_R FILLER_106_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_314 ();
 FILLER_ASAP7_75t_R FILLER_106_322 ();
 DECAPx10_ASAP7_75t_R FILLER_106_330 ();
 DECAPx6_ASAP7_75t_R FILLER_106_352 ();
 DECAPx4_ASAP7_75t_R FILLER_106_392 ();
 FILLER_ASAP7_75t_R FILLER_106_402 ();
 DECAPx4_ASAP7_75t_R FILLER_106_430 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_440 ();
 DECAPx1_ASAP7_75t_R FILLER_106_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_453 ();
 DECAPx1_ASAP7_75t_R FILLER_106_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_461 ();
 DECAPx1_ASAP7_75t_R FILLER_106_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_468 ();
 DECAPx1_ASAP7_75t_R FILLER_106_475 ();
 FILLER_ASAP7_75t_R FILLER_106_485 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_493 ();
 DECAPx2_ASAP7_75t_R FILLER_106_522 ();
 DECAPx6_ASAP7_75t_R FILLER_106_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_568 ();
 DECAPx10_ASAP7_75t_R FILLER_106_575 ();
 DECAPx4_ASAP7_75t_R FILLER_106_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_607 ();
 FILLER_ASAP7_75t_R FILLER_106_611 ();
 DECAPx4_ASAP7_75t_R FILLER_106_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_626 ();
 DECAPx4_ASAP7_75t_R FILLER_106_636 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_646 ();
 FILLER_ASAP7_75t_R FILLER_106_655 ();
 DECAPx1_ASAP7_75t_R FILLER_106_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_670 ();
 DECAPx4_ASAP7_75t_R FILLER_106_677 ();
 DECAPx2_ASAP7_75t_R FILLER_106_701 ();
 DECAPx4_ASAP7_75t_R FILLER_106_713 ();
 FILLER_ASAP7_75t_R FILLER_106_723 ();
 FILLER_ASAP7_75t_R FILLER_106_733 ();
 DECAPx1_ASAP7_75t_R FILLER_106_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_745 ();
 FILLER_ASAP7_75t_R FILLER_106_752 ();
 DECAPx1_ASAP7_75t_R FILLER_106_766 ();
 DECAPx10_ASAP7_75t_R FILLER_106_777 ();
 DECAPx2_ASAP7_75t_R FILLER_106_799 ();
 FILLER_ASAP7_75t_R FILLER_106_809 ();
 DECAPx4_ASAP7_75t_R FILLER_106_814 ();
 FILLER_ASAP7_75t_R FILLER_106_831 ();
 DECAPx10_ASAP7_75t_R FILLER_106_839 ();
 FILLER_ASAP7_75t_R FILLER_106_861 ();
 FILLER_ASAP7_75t_R FILLER_106_877 ();
 FILLER_ASAP7_75t_R FILLER_106_887 ();
 FILLER_ASAP7_75t_R FILLER_106_897 ();
 FILLER_ASAP7_75t_R FILLER_106_905 ();
 DECAPx1_ASAP7_75t_R FILLER_106_913 ();
 DECAPx4_ASAP7_75t_R FILLER_106_923 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_933 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_944 ();
 FILLER_ASAP7_75t_R FILLER_106_953 ();
 FILLER_ASAP7_75t_R FILLER_106_963 ();
 DECAPx1_ASAP7_75t_R FILLER_106_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_977 ();
 FILLER_ASAP7_75t_R FILLER_106_986 ();
 FILLER_ASAP7_75t_R FILLER_106_995 ();
 FILLER_ASAP7_75t_R FILLER_106_1004 ();
 FILLER_ASAP7_75t_R FILLER_106_1012 ();
 DECAPx4_ASAP7_75t_R FILLER_106_1022 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_106_1045 ();
 DECAPx4_ASAP7_75t_R FILLER_106_1059 ();
 FILLER_ASAP7_75t_R FILLER_106_1083 ();
 FILLER_ASAP7_75t_R FILLER_106_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1103 ();
 FILLER_ASAP7_75t_R FILLER_106_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1137 ();
 FILLER_ASAP7_75t_R FILLER_106_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_106_1171 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1193 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_1217 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_1224 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_1239 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_1249 ();
 FILLER_ASAP7_75t_R FILLER_106_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1269 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1287 ();
 FILLER_ASAP7_75t_R FILLER_106_1293 ();
 FILLER_ASAP7_75t_R FILLER_106_1302 ();
 FILLER_ASAP7_75t_R FILLER_106_1310 ();
 DECAPx6_ASAP7_75t_R FILLER_106_1315 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1335 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_1341 ();
 FILLER_ASAP7_75t_R FILLER_106_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_106_1371 ();
 DECAPx6_ASAP7_75t_R FILLER_107_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_107_16 ();
 DECAPx2_ASAP7_75t_R FILLER_107_25 ();
 FILLER_ASAP7_75t_R FILLER_107_37 ();
 DECAPx10_ASAP7_75t_R FILLER_107_42 ();
 DECAPx2_ASAP7_75t_R FILLER_107_64 ();
 FILLER_ASAP7_75t_R FILLER_107_70 ();
 FILLER_ASAP7_75t_R FILLER_107_98 ();
 DECAPx6_ASAP7_75t_R FILLER_107_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_122 ();
 DECAPx4_ASAP7_75t_R FILLER_107_129 ();
 FILLER_ASAP7_75t_R FILLER_107_139 ();
 DECAPx4_ASAP7_75t_R FILLER_107_144 ();
 FILLER_ASAP7_75t_R FILLER_107_160 ();
 FILLER_ASAP7_75t_R FILLER_107_170 ();
 DECAPx6_ASAP7_75t_R FILLER_107_180 ();
 DECAPx2_ASAP7_75t_R FILLER_107_194 ();
 DECAPx6_ASAP7_75t_R FILLER_107_206 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_107_220 ();
 DECAPx4_ASAP7_75t_R FILLER_107_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_239 ();
 FILLER_ASAP7_75t_R FILLER_107_248 ();
 DECAPx1_ASAP7_75t_R FILLER_107_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_260 ();
 FILLER_ASAP7_75t_R FILLER_107_269 ();
 DECAPx2_ASAP7_75t_R FILLER_107_277 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_107_283 ();
 DECAPx2_ASAP7_75t_R FILLER_107_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_298 ();
 FILLER_ASAP7_75t_R FILLER_107_302 ();
 DECAPx1_ASAP7_75t_R FILLER_107_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_334 ();
 DECAPx2_ASAP7_75t_R FILLER_107_341 ();
 DECAPx10_ASAP7_75t_R FILLER_107_353 ();
 DECAPx2_ASAP7_75t_R FILLER_107_375 ();
 DECAPx2_ASAP7_75t_R FILLER_107_384 ();
 DECAPx4_ASAP7_75t_R FILLER_107_393 ();
 FILLER_ASAP7_75t_R FILLER_107_403 ();
 DECAPx2_ASAP7_75t_R FILLER_107_411 ();
 FILLER_ASAP7_75t_R FILLER_107_423 ();
 FILLER_ASAP7_75t_R FILLER_107_431 ();
 DECAPx10_ASAP7_75t_R FILLER_107_436 ();
 FILLER_ASAP7_75t_R FILLER_107_458 ();
 FILLER_ASAP7_75t_R FILLER_107_466 ();
 FILLER_ASAP7_75t_R FILLER_107_476 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_107_504 ();
 FILLER_ASAP7_75t_R FILLER_107_510 ();
 FILLER_ASAP7_75t_R FILLER_107_520 ();
 FILLER_ASAP7_75t_R FILLER_107_528 ();
 DECAPx1_ASAP7_75t_R FILLER_107_536 ();
 FILLER_ASAP7_75t_R FILLER_107_543 ();
 DECAPx2_ASAP7_75t_R FILLER_107_555 ();
 FILLER_ASAP7_75t_R FILLER_107_567 ();
 FILLER_ASAP7_75t_R FILLER_107_577 ();
 FILLER_ASAP7_75t_R FILLER_107_586 ();
 FILLER_ASAP7_75t_R FILLER_107_594 ();
 DECAPx1_ASAP7_75t_R FILLER_107_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_607 ();
 DECAPx6_ASAP7_75t_R FILLER_107_611 ();
 DECAPx2_ASAP7_75t_R FILLER_107_625 ();
 FILLER_ASAP7_75t_R FILLER_107_637 ();
 DECAPx10_ASAP7_75t_R FILLER_107_645 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_107_667 ();
 DECAPx4_ASAP7_75t_R FILLER_107_682 ();
 FILLER_ASAP7_75t_R FILLER_107_698 ();
 FILLER_ASAP7_75t_R FILLER_107_720 ();
 DECAPx6_ASAP7_75t_R FILLER_107_729 ();
 FILLER_ASAP7_75t_R FILLER_107_743 ();
 DECAPx6_ASAP7_75t_R FILLER_107_748 ();
 FILLER_ASAP7_75t_R FILLER_107_762 ();
 FILLER_ASAP7_75t_R FILLER_107_767 ();
 DECAPx1_ASAP7_75t_R FILLER_107_777 ();
 DECAPx6_ASAP7_75t_R FILLER_107_789 ();
 DECAPx2_ASAP7_75t_R FILLER_107_803 ();
 DECAPx2_ASAP7_75t_R FILLER_107_818 ();
 FILLER_ASAP7_75t_R FILLER_107_824 ();
 FILLER_ASAP7_75t_R FILLER_107_833 ();
 DECAPx6_ASAP7_75t_R FILLER_107_844 ();
 DECAPx1_ASAP7_75t_R FILLER_107_858 ();
 DECAPx2_ASAP7_75t_R FILLER_107_870 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_107_876 ();
 FILLER_ASAP7_75t_R FILLER_107_887 ();
 DECAPx6_ASAP7_75t_R FILLER_107_897 ();
 FILLER_ASAP7_75t_R FILLER_107_911 ();
 FILLER_ASAP7_75t_R FILLER_107_923 ();
 DECAPx10_ASAP7_75t_R FILLER_107_927 ();
 DECAPx10_ASAP7_75t_R FILLER_107_949 ();
 DECAPx1_ASAP7_75t_R FILLER_107_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_975 ();
 FILLER_ASAP7_75t_R FILLER_107_983 ();
 FILLER_ASAP7_75t_R FILLER_107_992 ();
 FILLER_ASAP7_75t_R FILLER_107_1001 ();
 FILLER_ASAP7_75t_R FILLER_107_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1021 ();
 FILLER_ASAP7_75t_R FILLER_107_1035 ();
 FILLER_ASAP7_75t_R FILLER_107_1043 ();
 DECAPx4_ASAP7_75t_R FILLER_107_1071 ();
 FILLER_ASAP7_75t_R FILLER_107_1081 ();
 FILLER_ASAP7_75t_R FILLER_107_1109 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1114 ();
 FILLER_ASAP7_75t_R FILLER_107_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_107_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_1178 ();
 FILLER_ASAP7_75t_R FILLER_107_1186 ();
 FILLER_ASAP7_75t_R FILLER_107_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1199 ();
 FILLER_ASAP7_75t_R FILLER_107_1205 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_107_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1262 ();
 FILLER_ASAP7_75t_R FILLER_107_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_107_1296 ();
 DECAPx6_ASAP7_75t_R FILLER_107_1318 ();
 DECAPx2_ASAP7_75t_R FILLER_107_1352 ();
 FILLER_ASAP7_75t_R FILLER_107_1363 ();
 FILLER_ASAP7_75t_R FILLER_107_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_108_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_24 ();
 DECAPx1_ASAP7_75t_R FILLER_108_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_38 ();
 FILLER_ASAP7_75t_R FILLER_108_45 ();
 FILLER_ASAP7_75t_R FILLER_108_53 ();
 DECAPx1_ASAP7_75t_R FILLER_108_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_62 ();
 DECAPx1_ASAP7_75t_R FILLER_108_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_73 ();
 DECAPx2_ASAP7_75t_R FILLER_108_77 ();
 FILLER_ASAP7_75t_R FILLER_108_89 ();
 FILLER_ASAP7_75t_R FILLER_108_94 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_99 ();
 DECAPx2_ASAP7_75t_R FILLER_108_110 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_116 ();
 DECAPx10_ASAP7_75t_R FILLER_108_145 ();
 DECAPx4_ASAP7_75t_R FILLER_108_167 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_177 ();
 FILLER_ASAP7_75t_R FILLER_108_186 ();
 FILLER_ASAP7_75t_R FILLER_108_214 ();
 DECAPx1_ASAP7_75t_R FILLER_108_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_246 ();
 DECAPx2_ASAP7_75t_R FILLER_108_255 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_261 ();
 FILLER_ASAP7_75t_R FILLER_108_270 ();
 DECAPx6_ASAP7_75t_R FILLER_108_294 ();
 FILLER_ASAP7_75t_R FILLER_108_308 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_316 ();
 DECAPx2_ASAP7_75t_R FILLER_108_322 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_328 ();
 DECAPx6_ASAP7_75t_R FILLER_108_357 ();
 DECAPx6_ASAP7_75t_R FILLER_108_377 ();
 FILLER_ASAP7_75t_R FILLER_108_391 ();
 DECAPx2_ASAP7_75t_R FILLER_108_401 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_407 ();
 FILLER_ASAP7_75t_R FILLER_108_418 ();
 DECAPx1_ASAP7_75t_R FILLER_108_428 ();
 DECAPx1_ASAP7_75t_R FILLER_108_458 ();
 FILLER_ASAP7_75t_R FILLER_108_464 ();
 FILLER_ASAP7_75t_R FILLER_108_472 ();
 FILLER_ASAP7_75t_R FILLER_108_496 ();
 DECAPx1_ASAP7_75t_R FILLER_108_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_505 ();
 DECAPx10_ASAP7_75t_R FILLER_108_509 ();
 DECAPx2_ASAP7_75t_R FILLER_108_531 ();
 FILLER_ASAP7_75t_R FILLER_108_537 ();
 FILLER_ASAP7_75t_R FILLER_108_542 ();
 DECAPx2_ASAP7_75t_R FILLER_108_554 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_560 ();
 FILLER_ASAP7_75t_R FILLER_108_571 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_579 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_590 ();
 DECAPx1_ASAP7_75t_R FILLER_108_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_623 ();
 DECAPx2_ASAP7_75t_R FILLER_108_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_637 ();
 FILLER_ASAP7_75t_R FILLER_108_653 ();
 DECAPx1_ASAP7_75t_R FILLER_108_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_665 ();
 DECAPx6_ASAP7_75t_R FILLER_108_673 ();
 FILLER_ASAP7_75t_R FILLER_108_687 ();
 FILLER_ASAP7_75t_R FILLER_108_695 ();
 FILLER_ASAP7_75t_R FILLER_108_717 ();
 DECAPx6_ASAP7_75t_R FILLER_108_739 ();
 DECAPx10_ASAP7_75t_R FILLER_108_759 ();
 DECAPx1_ASAP7_75t_R FILLER_108_781 ();
 DECAPx2_ASAP7_75t_R FILLER_108_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_797 ();
 DECAPx10_ASAP7_75t_R FILLER_108_801 ();
 FILLER_ASAP7_75t_R FILLER_108_823 ();
 DECAPx1_ASAP7_75t_R FILLER_108_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_835 ();
 DECAPx1_ASAP7_75t_R FILLER_108_844 ();
 DECAPx2_ASAP7_75t_R FILLER_108_854 ();
 FILLER_ASAP7_75t_R FILLER_108_860 ();
 DECAPx10_ASAP7_75t_R FILLER_108_870 ();
 DECAPx6_ASAP7_75t_R FILLER_108_892 ();
 FILLER_ASAP7_75t_R FILLER_108_906 ();
 DECAPx2_ASAP7_75t_R FILLER_108_914 ();
 FILLER_ASAP7_75t_R FILLER_108_920 ();
 DECAPx2_ASAP7_75t_R FILLER_108_928 ();
 DECAPx2_ASAP7_75t_R FILLER_108_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_946 ();
 DECAPx4_ASAP7_75t_R FILLER_108_953 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_963 ();
 DECAPx10_ASAP7_75t_R FILLER_108_972 ();
 DECAPx1_ASAP7_75t_R FILLER_108_994 ();
 DECAPx6_ASAP7_75t_R FILLER_108_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1022 ();
 FILLER_ASAP7_75t_R FILLER_108_1035 ();
 FILLER_ASAP7_75t_R FILLER_108_1045 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1054 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1093 ();
 DECAPx4_ASAP7_75t_R FILLER_108_1109 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_1119 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1133 ();
 DECAPx4_ASAP7_75t_R FILLER_108_1137 ();
 FILLER_ASAP7_75t_R FILLER_108_1147 ();
 FILLER_ASAP7_75t_R FILLER_108_1156 ();
 FILLER_ASAP7_75t_R FILLER_108_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1170 ();
 DECAPx4_ASAP7_75t_R FILLER_108_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1210 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_108_1224 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1246 ();
 FILLER_ASAP7_75t_R FILLER_108_1256 ();
 DECAPx4_ASAP7_75t_R FILLER_108_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_1271 ();
 FILLER_ASAP7_75t_R FILLER_108_1279 ();
 FILLER_ASAP7_75t_R FILLER_108_1287 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_1292 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1301 ();
 FILLER_ASAP7_75t_R FILLER_108_1313 ();
 DECAPx2_ASAP7_75t_R FILLER_108_1321 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_1327 ();
 DECAPx1_ASAP7_75t_R FILLER_108_1336 ();
 FILLER_ASAP7_75t_R FILLER_108_1366 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_1374 ();
 DECAPx4_ASAP7_75t_R FILLER_109_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_12 ();
 DECAPx2_ASAP7_75t_R FILLER_109_19 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_25 ();
 DECAPx2_ASAP7_75t_R FILLER_109_54 ();
 DECAPx2_ASAP7_75t_R FILLER_109_86 ();
 FILLER_ASAP7_75t_R FILLER_109_92 ();
 FILLER_ASAP7_75t_R FILLER_109_100 ();
 DECAPx6_ASAP7_75t_R FILLER_109_108 ();
 DECAPx2_ASAP7_75t_R FILLER_109_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_128 ();
 FILLER_ASAP7_75t_R FILLER_109_135 ();
 DECAPx2_ASAP7_75t_R FILLER_109_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_146 ();
 DECAPx10_ASAP7_75t_R FILLER_109_150 ();
 DECAPx2_ASAP7_75t_R FILLER_109_172 ();
 FILLER_ASAP7_75t_R FILLER_109_184 ();
 FILLER_ASAP7_75t_R FILLER_109_193 ();
 FILLER_ASAP7_75t_R FILLER_109_201 ();
 FILLER_ASAP7_75t_R FILLER_109_209 ();
 DECAPx1_ASAP7_75t_R FILLER_109_214 ();
 DECAPx2_ASAP7_75t_R FILLER_109_224 ();
 DECAPx1_ASAP7_75t_R FILLER_109_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_237 ();
 FILLER_ASAP7_75t_R FILLER_109_244 ();
 FILLER_ASAP7_75t_R FILLER_109_252 ();
 DECAPx1_ASAP7_75t_R FILLER_109_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_264 ();
 FILLER_ASAP7_75t_R FILLER_109_268 ();
 FILLER_ASAP7_75t_R FILLER_109_276 ();
 DECAPx10_ASAP7_75t_R FILLER_109_304 ();
 DECAPx6_ASAP7_75t_R FILLER_109_326 ();
 DECAPx1_ASAP7_75t_R FILLER_109_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_344 ();
 DECAPx1_ASAP7_75t_R FILLER_109_348 ();
 DECAPx2_ASAP7_75t_R FILLER_109_355 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_361 ();
 DECAPx1_ASAP7_75t_R FILLER_109_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_394 ();
 FILLER_ASAP7_75t_R FILLER_109_403 ();
 DECAPx10_ASAP7_75t_R FILLER_109_411 ();
 DECAPx1_ASAP7_75t_R FILLER_109_433 ();
 DECAPx1_ASAP7_75t_R FILLER_109_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_447 ();
 DECAPx4_ASAP7_75t_R FILLER_109_474 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_484 ();
 DECAPx1_ASAP7_75t_R FILLER_109_497 ();
 FILLER_ASAP7_75t_R FILLER_109_523 ();
 DECAPx10_ASAP7_75t_R FILLER_109_535 ();
 DECAPx10_ASAP7_75t_R FILLER_109_557 ();
 DECAPx1_ASAP7_75t_R FILLER_109_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_583 ();
 DECAPx4_ASAP7_75t_R FILLER_109_591 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_601 ();
 DECAPx6_ASAP7_75t_R FILLER_109_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_624 ();
 DECAPx10_ASAP7_75t_R FILLER_109_637 ();
 DECAPx6_ASAP7_75t_R FILLER_109_659 ();
 FILLER_ASAP7_75t_R FILLER_109_682 ();
 DECAPx2_ASAP7_75t_R FILLER_109_691 ();
 DECAPx2_ASAP7_75t_R FILLER_109_706 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_712 ();
 DECAPx2_ASAP7_75t_R FILLER_109_722 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_728 ();
 FILLER_ASAP7_75t_R FILLER_109_742 ();
 FILLER_ASAP7_75t_R FILLER_109_753 ();
 FILLER_ASAP7_75t_R FILLER_109_761 ();
 DECAPx6_ASAP7_75t_R FILLER_109_769 ();
 DECAPx6_ASAP7_75t_R FILLER_109_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_823 ();
 DECAPx4_ASAP7_75t_R FILLER_109_834 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_854 ();
 DECAPx4_ASAP7_75t_R FILLER_109_864 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_874 ();
 FILLER_ASAP7_75t_R FILLER_109_884 ();
 DECAPx2_ASAP7_75t_R FILLER_109_894 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_900 ();
 FILLER_ASAP7_75t_R FILLER_109_911 ();
 FILLER_ASAP7_75t_R FILLER_109_923 ();
 FILLER_ASAP7_75t_R FILLER_109_927 ();
 DECAPx1_ASAP7_75t_R FILLER_109_936 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_947 ();
 DECAPx2_ASAP7_75t_R FILLER_109_957 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_963 ();
 DECAPx10_ASAP7_75t_R FILLER_109_980 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1024 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_109_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1055 ();
 FILLER_ASAP7_75t_R FILLER_109_1065 ();
 DECAPx4_ASAP7_75t_R FILLER_109_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1091 ();
 FILLER_ASAP7_75t_R FILLER_109_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1121 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1143 ();
 FILLER_ASAP7_75t_R FILLER_109_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_109_1185 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1192 ();
 FILLER_ASAP7_75t_R FILLER_109_1206 ();
 DECAPx6_ASAP7_75t_R FILLER_109_1214 ();
 FILLER_ASAP7_75t_R FILLER_109_1228 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1237 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_109_1274 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_1296 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1309 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1315 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1330 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1337 ();
 FILLER_ASAP7_75t_R FILLER_109_1343 ();
 FILLER_ASAP7_75t_R FILLER_109_1348 ();
 FILLER_ASAP7_75t_R FILLER_109_1355 ();
 DECAPx2_ASAP7_75t_R FILLER_109_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_1369 ();
 FILLER_ASAP7_75t_R FILLER_109_1375 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_2 ();
 FILLER_ASAP7_75t_R FILLER_110_31 ();
 DECAPx2_ASAP7_75t_R FILLER_110_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_46 ();
 DECAPx2_ASAP7_75t_R FILLER_110_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_61 ();
 DECAPx10_ASAP7_75t_R FILLER_110_68 ();
 DECAPx2_ASAP7_75t_R FILLER_110_90 ();
 DECAPx10_ASAP7_75t_R FILLER_110_102 ();
 DECAPx2_ASAP7_75t_R FILLER_110_124 ();
 FILLER_ASAP7_75t_R FILLER_110_130 ();
 DECAPx2_ASAP7_75t_R FILLER_110_138 ();
 FILLER_ASAP7_75t_R FILLER_110_144 ();
 FILLER_ASAP7_75t_R FILLER_110_152 ();
 FILLER_ASAP7_75t_R FILLER_110_162 ();
 FILLER_ASAP7_75t_R FILLER_110_172 ();
 DECAPx1_ASAP7_75t_R FILLER_110_182 ();
 FILLER_ASAP7_75t_R FILLER_110_193 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_202 ();
 DECAPx10_ASAP7_75t_R FILLER_110_211 ();
 DECAPx4_ASAP7_75t_R FILLER_110_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_243 ();
 DECAPx2_ASAP7_75t_R FILLER_110_255 ();
 FILLER_ASAP7_75t_R FILLER_110_261 ();
 FILLER_ASAP7_75t_R FILLER_110_285 ();
 FILLER_ASAP7_75t_R FILLER_110_293 ();
 DECAPx2_ASAP7_75t_R FILLER_110_298 ();
 FILLER_ASAP7_75t_R FILLER_110_304 ();
 DECAPx4_ASAP7_75t_R FILLER_110_312 ();
 DECAPx2_ASAP7_75t_R FILLER_110_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_335 ();
 FILLER_ASAP7_75t_R FILLER_110_342 ();
 DECAPx4_ASAP7_75t_R FILLER_110_350 ();
 FILLER_ASAP7_75t_R FILLER_110_366 ();
 DECAPx1_ASAP7_75t_R FILLER_110_374 ();
 FILLER_ASAP7_75t_R FILLER_110_385 ();
 FILLER_ASAP7_75t_R FILLER_110_394 ();
 DECAPx2_ASAP7_75t_R FILLER_110_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_409 ();
 FILLER_ASAP7_75t_R FILLER_110_418 ();
 DECAPx1_ASAP7_75t_R FILLER_110_426 ();
 FILLER_ASAP7_75t_R FILLER_110_433 ();
 DECAPx2_ASAP7_75t_R FILLER_110_441 ();
 FILLER_ASAP7_75t_R FILLER_110_450 ();
 DECAPx1_ASAP7_75t_R FILLER_110_458 ();
 FILLER_ASAP7_75t_R FILLER_110_464 ();
 DECAPx1_ASAP7_75t_R FILLER_110_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_473 ();
 FILLER_ASAP7_75t_R FILLER_110_486 ();
 FILLER_ASAP7_75t_R FILLER_110_514 ();
 DECAPx1_ASAP7_75t_R FILLER_110_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_527 ();
 DECAPx2_ASAP7_75t_R FILLER_110_538 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_544 ();
 DECAPx4_ASAP7_75t_R FILLER_110_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_569 ();
 DECAPx1_ASAP7_75t_R FILLER_110_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_580 ();
 FILLER_ASAP7_75t_R FILLER_110_603 ();
 FILLER_ASAP7_75t_R FILLER_110_611 ();
 DECAPx2_ASAP7_75t_R FILLER_110_616 ();
 DECAPx6_ASAP7_75t_R FILLER_110_628 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_642 ();
 FILLER_ASAP7_75t_R FILLER_110_651 ();
 FILLER_ASAP7_75t_R FILLER_110_660 ();
 FILLER_ASAP7_75t_R FILLER_110_669 ();
 FILLER_ASAP7_75t_R FILLER_110_691 ();
 DECAPx2_ASAP7_75t_R FILLER_110_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_707 ();
 FILLER_ASAP7_75t_R FILLER_110_714 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_730 ();
 DECAPx6_ASAP7_75t_R FILLER_110_739 ();
 FILLER_ASAP7_75t_R FILLER_110_753 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_762 ();
 FILLER_ASAP7_75t_R FILLER_110_773 ();
 DECAPx2_ASAP7_75t_R FILLER_110_781 ();
 FILLER_ASAP7_75t_R FILLER_110_787 ();
 FILLER_ASAP7_75t_R FILLER_110_795 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_800 ();
 FILLER_ASAP7_75t_R FILLER_110_809 ();
 DECAPx1_ASAP7_75t_R FILLER_110_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_825 ();
 DECAPx6_ASAP7_75t_R FILLER_110_836 ();
 FILLER_ASAP7_75t_R FILLER_110_850 ();
 DECAPx6_ASAP7_75t_R FILLER_110_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_878 ();
 FILLER_ASAP7_75t_R FILLER_110_885 ();
 DECAPx2_ASAP7_75t_R FILLER_110_893 ();
 FILLER_ASAP7_75t_R FILLER_110_899 ();
 FILLER_ASAP7_75t_R FILLER_110_907 ();
 FILLER_ASAP7_75t_R FILLER_110_915 ();
 DECAPx4_ASAP7_75t_R FILLER_110_923 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_933 ();
 DECAPx2_ASAP7_75t_R FILLER_110_942 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_948 ();
 DECAPx2_ASAP7_75t_R FILLER_110_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_964 ();
 FILLER_ASAP7_75t_R FILLER_110_971 ();
 DECAPx2_ASAP7_75t_R FILLER_110_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_987 ();
 DECAPx6_ASAP7_75t_R FILLER_110_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1010 ();
 FILLER_ASAP7_75t_R FILLER_110_1019 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_110_1042 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1064 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1094 ();
 FILLER_ASAP7_75t_R FILLER_110_1104 ();
 FILLER_ASAP7_75t_R FILLER_110_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_110_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1158 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1183 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1190 ();
 FILLER_ASAP7_75t_R FILLER_110_1204 ();
 FILLER_ASAP7_75t_R FILLER_110_1226 ();
 DECAPx4_ASAP7_75t_R FILLER_110_1254 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1274 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1280 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1307 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_1313 ();
 DECAPx6_ASAP7_75t_R FILLER_110_1322 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1342 ();
 DECAPx2_ASAP7_75t_R FILLER_110_1351 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_1357 ();
 FILLER_ASAP7_75t_R FILLER_110_1368 ();
 FILLER_ASAP7_75t_R FILLER_110_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_111_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_8 ();
 DECAPx1_ASAP7_75t_R FILLER_111_15 ();
 DECAPx1_ASAP7_75t_R FILLER_111_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_26 ();
 FILLER_ASAP7_75t_R FILLER_111_34 ();
 DECAPx2_ASAP7_75t_R FILLER_111_43 ();
 FILLER_ASAP7_75t_R FILLER_111_49 ();
 DECAPx6_ASAP7_75t_R FILLER_111_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_73 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_81 ();
 FILLER_ASAP7_75t_R FILLER_111_110 ();
 FILLER_ASAP7_75t_R FILLER_111_122 ();
 DECAPx1_ASAP7_75t_R FILLER_111_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_154 ();
 FILLER_ASAP7_75t_R FILLER_111_158 ();
 DECAPx2_ASAP7_75t_R FILLER_111_168 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_174 ();
 FILLER_ASAP7_75t_R FILLER_111_184 ();
 DECAPx1_ASAP7_75t_R FILLER_111_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_197 ();
 FILLER_ASAP7_75t_R FILLER_111_224 ();
 DECAPx6_ASAP7_75t_R FILLER_111_232 ();
 DECAPx1_ASAP7_75t_R FILLER_111_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_250 ();
 DECAPx2_ASAP7_75t_R FILLER_111_259 ();
 FILLER_ASAP7_75t_R FILLER_111_265 ();
 DECAPx6_ASAP7_75t_R FILLER_111_273 ();
 DECAPx2_ASAP7_75t_R FILLER_111_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_293 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_320 ();
 FILLER_ASAP7_75t_R FILLER_111_331 ();
 DECAPx1_ASAP7_75t_R FILLER_111_336 ();
 FILLER_ASAP7_75t_R FILLER_111_366 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_375 ();
 DECAPx2_ASAP7_75t_R FILLER_111_381 ();
 FILLER_ASAP7_75t_R FILLER_111_394 ();
 FILLER_ASAP7_75t_R FILLER_111_403 ();
 FILLER_ASAP7_75t_R FILLER_111_412 ();
 DECAPx10_ASAP7_75t_R FILLER_111_422 ();
 DECAPx6_ASAP7_75t_R FILLER_111_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_458 ();
 FILLER_ASAP7_75t_R FILLER_111_474 ();
 DECAPx2_ASAP7_75t_R FILLER_111_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_492 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_503 ();
 FILLER_ASAP7_75t_R FILLER_111_512 ();
 DECAPx2_ASAP7_75t_R FILLER_111_524 ();
 DECAPx6_ASAP7_75t_R FILLER_111_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_556 ();
 DECAPx2_ASAP7_75t_R FILLER_111_567 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_573 ();
 FILLER_ASAP7_75t_R FILLER_111_588 ();
 FILLER_ASAP7_75t_R FILLER_111_596 ();
 DECAPx1_ASAP7_75t_R FILLER_111_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_628 ();
 FILLER_ASAP7_75t_R FILLER_111_635 ();
 FILLER_ASAP7_75t_R FILLER_111_645 ();
 DECAPx6_ASAP7_75t_R FILLER_111_653 ();
 FILLER_ASAP7_75t_R FILLER_111_667 ();
 DECAPx6_ASAP7_75t_R FILLER_111_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_690 ();
 FILLER_ASAP7_75t_R FILLER_111_698 ();
 DECAPx4_ASAP7_75t_R FILLER_111_706 ();
 FILLER_ASAP7_75t_R FILLER_111_716 ();
 DECAPx4_ASAP7_75t_R FILLER_111_724 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_734 ();
 DECAPx6_ASAP7_75t_R FILLER_111_745 ();
 DECAPx6_ASAP7_75t_R FILLER_111_765 ();
 DECAPx1_ASAP7_75t_R FILLER_111_779 ();
 DECAPx2_ASAP7_75t_R FILLER_111_794 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_800 ();
 FILLER_ASAP7_75t_R FILLER_111_807 ();
 DECAPx10_ASAP7_75t_R FILLER_111_815 ();
 DECAPx1_ASAP7_75t_R FILLER_111_837 ();
 DECAPx6_ASAP7_75t_R FILLER_111_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_861 ();
 FILLER_ASAP7_75t_R FILLER_111_866 ();
 FILLER_ASAP7_75t_R FILLER_111_875 ();
 DECAPx10_ASAP7_75t_R FILLER_111_883 ();
 DECAPx6_ASAP7_75t_R FILLER_111_905 ();
 DECAPx2_ASAP7_75t_R FILLER_111_919 ();
 DECAPx2_ASAP7_75t_R FILLER_111_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_933 ();
 DECAPx10_ASAP7_75t_R FILLER_111_940 ();
 DECAPx2_ASAP7_75t_R FILLER_111_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_968 ();
 DECAPx1_ASAP7_75t_R FILLER_111_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_979 ();
 FILLER_ASAP7_75t_R FILLER_111_988 ();
 DECAPx2_ASAP7_75t_R FILLER_111_1005 ();
 FILLER_ASAP7_75t_R FILLER_111_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_111_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1036 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_1043 ();
 FILLER_ASAP7_75t_R FILLER_111_1058 ();
 FILLER_ASAP7_75t_R FILLER_111_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1094 ();
 FILLER_ASAP7_75t_R FILLER_111_1115 ();
 FILLER_ASAP7_75t_R FILLER_111_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_111_1128 ();
 FILLER_ASAP7_75t_R FILLER_111_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1150 ();
 FILLER_ASAP7_75t_R FILLER_111_1157 ();
 FILLER_ASAP7_75t_R FILLER_111_1185 ();
 FILLER_ASAP7_75t_R FILLER_111_1194 ();
 FILLER_ASAP7_75t_R FILLER_111_1216 ();
 FILLER_ASAP7_75t_R FILLER_111_1224 ();
 DECAPx4_ASAP7_75t_R FILLER_111_1232 ();
 DECAPx2_ASAP7_75t_R FILLER_111_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1251 ();
 FILLER_ASAP7_75t_R FILLER_111_1278 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_1283 ();
 FILLER_ASAP7_75t_R FILLER_111_1294 ();
 DECAPx6_ASAP7_75t_R FILLER_111_1299 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1313 ();
 DECAPx2_ASAP7_75t_R FILLER_111_1327 ();
 FILLER_ASAP7_75t_R FILLER_111_1339 ();
 DECAPx1_ASAP7_75t_R FILLER_111_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_1348 ();
 FILLER_ASAP7_75t_R FILLER_111_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_112_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_16 ();
 DECAPx1_ASAP7_75t_R FILLER_112_23 ();
 FILLER_ASAP7_75t_R FILLER_112_34 ();
 DECAPx1_ASAP7_75t_R FILLER_112_39 ();
 FILLER_ASAP7_75t_R FILLER_112_49 ();
 FILLER_ASAP7_75t_R FILLER_112_57 ();
 DECAPx4_ASAP7_75t_R FILLER_112_65 ();
 DECAPx2_ASAP7_75t_R FILLER_112_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_89 ();
 FILLER_ASAP7_75t_R FILLER_112_96 ();
 DECAPx4_ASAP7_75t_R FILLER_112_101 ();
 FILLER_ASAP7_75t_R FILLER_112_111 ();
 DECAPx2_ASAP7_75t_R FILLER_112_120 ();
 DECAPx2_ASAP7_75t_R FILLER_112_132 ();
 DECAPx6_ASAP7_75t_R FILLER_112_141 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_155 ();
 DECAPx1_ASAP7_75t_R FILLER_112_164 ();
 FILLER_ASAP7_75t_R FILLER_112_174 ();
 FILLER_ASAP7_75t_R FILLER_112_182 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_210 ();
 FILLER_ASAP7_75t_R FILLER_112_219 ();
 FILLER_ASAP7_75t_R FILLER_112_235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_245 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_260 ();
 FILLER_ASAP7_75t_R FILLER_112_289 ();
 DECAPx1_ASAP7_75t_R FILLER_112_297 ();
 FILLER_ASAP7_75t_R FILLER_112_307 ();
 DECAPx4_ASAP7_75t_R FILLER_112_312 ();
 FILLER_ASAP7_75t_R FILLER_112_328 ();
 DECAPx1_ASAP7_75t_R FILLER_112_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_340 ();
 FILLER_ASAP7_75t_R FILLER_112_349 ();
 FILLER_ASAP7_75t_R FILLER_112_357 ();
 DECAPx2_ASAP7_75t_R FILLER_112_362 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_368 ();
 DECAPx4_ASAP7_75t_R FILLER_112_377 ();
 FILLER_ASAP7_75t_R FILLER_112_393 ();
 FILLER_ASAP7_75t_R FILLER_112_406 ();
 FILLER_ASAP7_75t_R FILLER_112_414 ();
 DECAPx1_ASAP7_75t_R FILLER_112_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_426 ();
 DECAPx2_ASAP7_75t_R FILLER_112_433 ();
 FILLER_ASAP7_75t_R FILLER_112_439 ();
 DECAPx6_ASAP7_75t_R FILLER_112_444 ();
 DECAPx1_ASAP7_75t_R FILLER_112_458 ();
 DECAPx2_ASAP7_75t_R FILLER_112_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_470 ();
 DECAPx2_ASAP7_75t_R FILLER_112_495 ();
 FILLER_ASAP7_75t_R FILLER_112_501 ();
 DECAPx2_ASAP7_75t_R FILLER_112_506 ();
 DECAPx6_ASAP7_75t_R FILLER_112_515 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_529 ();
 DECAPx4_ASAP7_75t_R FILLER_112_535 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_545 ();
 DECAPx4_ASAP7_75t_R FILLER_112_554 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_564 ();
 DECAPx1_ASAP7_75t_R FILLER_112_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_581 ();
 DECAPx1_ASAP7_75t_R FILLER_112_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_598 ();
 DECAPx10_ASAP7_75t_R FILLER_112_606 ();
 DECAPx10_ASAP7_75t_R FILLER_112_634 ();
 DECAPx6_ASAP7_75t_R FILLER_112_656 ();
 DECAPx2_ASAP7_75t_R FILLER_112_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_676 ();
 DECAPx4_ASAP7_75t_R FILLER_112_683 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_693 ();
 DECAPx1_ASAP7_75t_R FILLER_112_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_715 ();
 FILLER_ASAP7_75t_R FILLER_112_724 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_734 ();
 DECAPx4_ASAP7_75t_R FILLER_112_749 ();
 DECAPx4_ASAP7_75t_R FILLER_112_767 ();
 FILLER_ASAP7_75t_R FILLER_112_777 ();
 DECAPx10_ASAP7_75t_R FILLER_112_785 ();
 DECAPx6_ASAP7_75t_R FILLER_112_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_821 ();
 DECAPx2_ASAP7_75t_R FILLER_112_825 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_831 ();
 FILLER_ASAP7_75t_R FILLER_112_840 ();
 DECAPx4_ASAP7_75t_R FILLER_112_852 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_862 ();
 DECAPx10_ASAP7_75t_R FILLER_112_871 ();
 DECAPx6_ASAP7_75t_R FILLER_112_893 ();
 DECAPx2_ASAP7_75t_R FILLER_112_913 ();
 DECAPx6_ASAP7_75t_R FILLER_112_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_945 ();
 FILLER_ASAP7_75t_R FILLER_112_954 ();
 DECAPx2_ASAP7_75t_R FILLER_112_962 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_968 ();
 DECAPx6_ASAP7_75t_R FILLER_112_977 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_991 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_1001 ();
 FILLER_ASAP7_75t_R FILLER_112_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1040 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1049 ();
 FILLER_ASAP7_75t_R FILLER_112_1073 ();
 FILLER_ASAP7_75t_R FILLER_112_1085 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_1095 ();
 DECAPx4_ASAP7_75t_R FILLER_112_1104 ();
 FILLER_ASAP7_75t_R FILLER_112_1114 ();
 FILLER_ASAP7_75t_R FILLER_112_1122 ();
 FILLER_ASAP7_75t_R FILLER_112_1130 ();
 FILLER_ASAP7_75t_R FILLER_112_1142 ();
 DECAPx4_ASAP7_75t_R FILLER_112_1147 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_1157 ();
 FILLER_ASAP7_75t_R FILLER_112_1168 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_1180 ();
 FILLER_ASAP7_75t_R FILLER_112_1191 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1199 ();
 DECAPx2_ASAP7_75t_R FILLER_112_1215 ();
 DECAPx6_ASAP7_75t_R FILLER_112_1247 ();
 FILLER_ASAP7_75t_R FILLER_112_1267 ();
 FILLER_ASAP7_75t_R FILLER_112_1277 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1282 ();
 DECAPx4_ASAP7_75t_R FILLER_112_1292 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_112_1314 ();
 FILLER_ASAP7_75t_R FILLER_112_1336 ();
 FILLER_ASAP7_75t_R FILLER_112_1347 ();
 DECAPx1_ASAP7_75t_R FILLER_112_1357 ();
 FILLER_ASAP7_75t_R FILLER_112_1369 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_1374 ();
 FILLER_ASAP7_75t_R FILLER_113_2 ();
 DECAPx2_ASAP7_75t_R FILLER_113_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_36 ();
 DECAPx1_ASAP7_75t_R FILLER_113_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_49 ();
 FILLER_ASAP7_75t_R FILLER_113_56 ();
 FILLER_ASAP7_75t_R FILLER_113_64 ();
 DECAPx2_ASAP7_75t_R FILLER_113_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_78 ();
 DECAPx10_ASAP7_75t_R FILLER_113_91 ();
 DECAPx10_ASAP7_75t_R FILLER_113_113 ();
 DECAPx2_ASAP7_75t_R FILLER_113_135 ();
 FILLER_ASAP7_75t_R FILLER_113_141 ();
 DECAPx4_ASAP7_75t_R FILLER_113_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_159 ();
 FILLER_ASAP7_75t_R FILLER_113_163 ();
 FILLER_ASAP7_75t_R FILLER_113_173 ();
 DECAPx2_ASAP7_75t_R FILLER_113_181 ();
 FILLER_ASAP7_75t_R FILLER_113_187 ();
 DECAPx1_ASAP7_75t_R FILLER_113_195 ();
 DECAPx4_ASAP7_75t_R FILLER_113_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_212 ();
 DECAPx2_ASAP7_75t_R FILLER_113_216 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_222 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_231 ();
 FILLER_ASAP7_75t_R FILLER_113_240 ();
 FILLER_ASAP7_75t_R FILLER_113_264 ();
 FILLER_ASAP7_75t_R FILLER_113_272 ();
 FILLER_ASAP7_75t_R FILLER_113_277 ();
 FILLER_ASAP7_75t_R FILLER_113_285 ();
 DECAPx10_ASAP7_75t_R FILLER_113_293 ();
 DECAPx10_ASAP7_75t_R FILLER_113_315 ();
 DECAPx10_ASAP7_75t_R FILLER_113_337 ();
 DECAPx6_ASAP7_75t_R FILLER_113_359 ();
 FILLER_ASAP7_75t_R FILLER_113_389 ();
 DECAPx4_ASAP7_75t_R FILLER_113_405 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_415 ();
 FILLER_ASAP7_75t_R FILLER_113_424 ();
 FILLER_ASAP7_75t_R FILLER_113_452 ();
 DECAPx4_ASAP7_75t_R FILLER_113_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_467 ();
 FILLER_ASAP7_75t_R FILLER_113_480 ();
 DECAPx6_ASAP7_75t_R FILLER_113_490 ();
 DECAPx10_ASAP7_75t_R FILLER_113_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_533 ();
 DECAPx1_ASAP7_75t_R FILLER_113_540 ();
 FILLER_ASAP7_75t_R FILLER_113_550 ();
 FILLER_ASAP7_75t_R FILLER_113_560 ();
 DECAPx10_ASAP7_75t_R FILLER_113_568 ();
 FILLER_ASAP7_75t_R FILLER_113_596 ();
 DECAPx2_ASAP7_75t_R FILLER_113_624 ();
 DECAPx2_ASAP7_75t_R FILLER_113_640 ();
 DECAPx2_ASAP7_75t_R FILLER_113_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_659 ();
 DECAPx4_ASAP7_75t_R FILLER_113_666 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_676 ();
 DECAPx2_ASAP7_75t_R FILLER_113_687 ();
 FILLER_ASAP7_75t_R FILLER_113_693 ();
 FILLER_ASAP7_75t_R FILLER_113_715 ();
 FILLER_ASAP7_75t_R FILLER_113_727 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_735 ();
 DECAPx2_ASAP7_75t_R FILLER_113_750 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_756 ();
 DECAPx4_ASAP7_75t_R FILLER_113_768 ();
 FILLER_ASAP7_75t_R FILLER_113_787 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_795 ();
 DECAPx4_ASAP7_75t_R FILLER_113_808 ();
 FILLER_ASAP7_75t_R FILLER_113_827 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_835 ();
 DECAPx6_ASAP7_75t_R FILLER_113_841 ();
 FILLER_ASAP7_75t_R FILLER_113_855 ();
 FILLER_ASAP7_75t_R FILLER_113_883 ();
 FILLER_ASAP7_75t_R FILLER_113_894 ();
 FILLER_ASAP7_75t_R FILLER_113_899 ();
 DECAPx4_ASAP7_75t_R FILLER_113_915 ();
 FILLER_ASAP7_75t_R FILLER_113_927 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_936 ();
 FILLER_ASAP7_75t_R FILLER_113_951 ();
 DECAPx2_ASAP7_75t_R FILLER_113_959 ();
 FILLER_ASAP7_75t_R FILLER_113_965 ();
 DECAPx4_ASAP7_75t_R FILLER_113_979 ();
 DECAPx2_ASAP7_75t_R FILLER_113_996 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1008 ();
 FILLER_ASAP7_75t_R FILLER_113_1018 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1049 ();
 FILLER_ASAP7_75t_R FILLER_113_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1067 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_1073 ();
 FILLER_ASAP7_75t_R FILLER_113_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1120 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_1126 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1165 ();
 FILLER_ASAP7_75t_R FILLER_113_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_113_1198 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_1220 ();
 DECAPx1_ASAP7_75t_R FILLER_113_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1235 ();
 DECAPx6_ASAP7_75t_R FILLER_113_1239 ();
 DECAPx6_ASAP7_75t_R FILLER_113_1259 ();
 DECAPx6_ASAP7_75t_R FILLER_113_1276 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1290 ();
 FILLER_ASAP7_75t_R FILLER_113_1299 ();
 FILLER_ASAP7_75t_R FILLER_113_1307 ();
 FILLER_ASAP7_75t_R FILLER_113_1335 ();
 DECAPx4_ASAP7_75t_R FILLER_113_1347 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_1357 ();
 DECAPx2_ASAP7_75t_R FILLER_113_1364 ();
 FILLER_ASAP7_75t_R FILLER_113_1375 ();
 DECAPx4_ASAP7_75t_R FILLER_114_2 ();
 FILLER_ASAP7_75t_R FILLER_114_18 ();
 DECAPx2_ASAP7_75t_R FILLER_114_23 ();
 FILLER_ASAP7_75t_R FILLER_114_35 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_45 ();
 DECAPx10_ASAP7_75t_R FILLER_114_54 ();
 DECAPx6_ASAP7_75t_R FILLER_114_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_90 ();
 DECAPx2_ASAP7_75t_R FILLER_114_97 ();
 FILLER_ASAP7_75t_R FILLER_114_103 ();
 DECAPx1_ASAP7_75t_R FILLER_114_131 ();
 DECAPx10_ASAP7_75t_R FILLER_114_161 ();
 DECAPx10_ASAP7_75t_R FILLER_114_183 ();
 DECAPx10_ASAP7_75t_R FILLER_114_205 ();
 DECAPx2_ASAP7_75t_R FILLER_114_227 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_233 ();
 FILLER_ASAP7_75t_R FILLER_114_242 ();
 DECAPx6_ASAP7_75t_R FILLER_114_251 ();
 DECAPx1_ASAP7_75t_R FILLER_114_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_269 ();
 DECAPx2_ASAP7_75t_R FILLER_114_276 ();
 DECAPx4_ASAP7_75t_R FILLER_114_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_298 ();
 DECAPx10_ASAP7_75t_R FILLER_114_305 ();
 FILLER_ASAP7_75t_R FILLER_114_327 ();
 DECAPx6_ASAP7_75t_R FILLER_114_339 ();
 DECAPx2_ASAP7_75t_R FILLER_114_353 ();
 DECAPx2_ASAP7_75t_R FILLER_114_365 ();
 FILLER_ASAP7_75t_R FILLER_114_371 ();
 FILLER_ASAP7_75t_R FILLER_114_376 ();
 DECAPx10_ASAP7_75t_R FILLER_114_388 ();
 DECAPx10_ASAP7_75t_R FILLER_114_410 ();
 FILLER_ASAP7_75t_R FILLER_114_432 ();
 FILLER_ASAP7_75t_R FILLER_114_460 ();
 FILLER_ASAP7_75t_R FILLER_114_464 ();
 DECAPx4_ASAP7_75t_R FILLER_114_469 ();
 FILLER_ASAP7_75t_R FILLER_114_479 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_487 ();
 FILLER_ASAP7_75t_R FILLER_114_516 ();
 DECAPx1_ASAP7_75t_R FILLER_114_521 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_537 ();
 FILLER_ASAP7_75t_R FILLER_114_546 ();
 FILLER_ASAP7_75t_R FILLER_114_570 ();
 DECAPx4_ASAP7_75t_R FILLER_114_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_588 ();
 FILLER_ASAP7_75t_R FILLER_114_595 ();
 DECAPx2_ASAP7_75t_R FILLER_114_603 ();
 FILLER_ASAP7_75t_R FILLER_114_609 ();
 FILLER_ASAP7_75t_R FILLER_114_614 ();
 DECAPx6_ASAP7_75t_R FILLER_114_622 ();
 DECAPx1_ASAP7_75t_R FILLER_114_636 ();
 FILLER_ASAP7_75t_R FILLER_114_646 ();
 DECAPx2_ASAP7_75t_R FILLER_114_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_662 ();
 FILLER_ASAP7_75t_R FILLER_114_669 ();
 FILLER_ASAP7_75t_R FILLER_114_677 ();
 DECAPx1_ASAP7_75t_R FILLER_114_691 ();
 DECAPx2_ASAP7_75t_R FILLER_114_709 ();
 FILLER_ASAP7_75t_R FILLER_114_715 ();
 DECAPx4_ASAP7_75t_R FILLER_114_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_734 ();
 DECAPx1_ASAP7_75t_R FILLER_114_742 ();
 DECAPx2_ASAP7_75t_R FILLER_114_752 ();
 FILLER_ASAP7_75t_R FILLER_114_758 ();
 DECAPx6_ASAP7_75t_R FILLER_114_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_780 ();
 DECAPx1_ASAP7_75t_R FILLER_114_793 ();
 FILLER_ASAP7_75t_R FILLER_114_817 ();
 FILLER_ASAP7_75t_R FILLER_114_828 ();
 DECAPx4_ASAP7_75t_R FILLER_114_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_848 ();
 FILLER_ASAP7_75t_R FILLER_114_855 ();
 DECAPx1_ASAP7_75t_R FILLER_114_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_864 ();
 FILLER_ASAP7_75t_R FILLER_114_871 ();
 DECAPx4_ASAP7_75t_R FILLER_114_876 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_886 ();
 FILLER_ASAP7_75t_R FILLER_114_897 ();
 DECAPx2_ASAP7_75t_R FILLER_114_905 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_911 ();
 DECAPx1_ASAP7_75t_R FILLER_114_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_925 ();
 DECAPx6_ASAP7_75t_R FILLER_114_932 ();
 FILLER_ASAP7_75t_R FILLER_114_946 ();
 FILLER_ASAP7_75t_R FILLER_114_954 ();
 FILLER_ASAP7_75t_R FILLER_114_959 ();
 FILLER_ASAP7_75t_R FILLER_114_967 ();
 FILLER_ASAP7_75t_R FILLER_114_976 ();
 FILLER_ASAP7_75t_R FILLER_114_988 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1014 ();
 FILLER_ASAP7_75t_R FILLER_114_1040 ();
 FILLER_ASAP7_75t_R FILLER_114_1047 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1079 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1099 ();
 FILLER_ASAP7_75t_R FILLER_114_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_114_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_114_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_114_1184 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1206 ();
 DECAPx4_ASAP7_75t_R FILLER_114_1213 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1243 ();
 FILLER_ASAP7_75t_R FILLER_114_1256 ();
 DECAPx6_ASAP7_75t_R FILLER_114_1264 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_1278 ();
 FILLER_ASAP7_75t_R FILLER_114_1284 ();
 FILLER_ASAP7_75t_R FILLER_114_1292 ();
 DECAPx1_ASAP7_75t_R FILLER_114_1303 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1307 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1316 ();
 FILLER_ASAP7_75t_R FILLER_114_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_114_1327 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1349 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_1355 ();
 DECAPx2_ASAP7_75t_R FILLER_114_1364 ();
 FILLER_ASAP7_75t_R FILLER_114_1375 ();
 DECAPx4_ASAP7_75t_R FILLER_115_2 ();
 FILLER_ASAP7_75t_R FILLER_115_12 ();
 FILLER_ASAP7_75t_R FILLER_115_20 ();
 DECAPx1_ASAP7_75t_R FILLER_115_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_29 ();
 DECAPx10_ASAP7_75t_R FILLER_115_33 ();
 DECAPx6_ASAP7_75t_R FILLER_115_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_69 ();
 DECAPx4_ASAP7_75t_R FILLER_115_76 ();
 FILLER_ASAP7_75t_R FILLER_115_86 ();
 DECAPx1_ASAP7_75t_R FILLER_115_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_118 ();
 FILLER_ASAP7_75t_R FILLER_115_125 ();
 DECAPx2_ASAP7_75t_R FILLER_115_130 ();
 FILLER_ASAP7_75t_R FILLER_115_136 ();
 DECAPx2_ASAP7_75t_R FILLER_115_144 ();
 DECAPx6_ASAP7_75t_R FILLER_115_153 ();
 FILLER_ASAP7_75t_R FILLER_115_167 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_175 ();
 DECAPx4_ASAP7_75t_R FILLER_115_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_210 ();
 DECAPx6_ASAP7_75t_R FILLER_115_217 ();
 DECAPx1_ASAP7_75t_R FILLER_115_231 ();
 DECAPx2_ASAP7_75t_R FILLER_115_245 ();
 DECAPx2_ASAP7_75t_R FILLER_115_257 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_263 ();
 DECAPx6_ASAP7_75t_R FILLER_115_272 ();
 FILLER_ASAP7_75t_R FILLER_115_312 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_317 ();
 FILLER_ASAP7_75t_R FILLER_115_328 ();
 DECAPx1_ASAP7_75t_R FILLER_115_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_340 ();
 FILLER_ASAP7_75t_R FILLER_115_347 ();
 DECAPx10_ASAP7_75t_R FILLER_115_375 ();
 FILLER_ASAP7_75t_R FILLER_115_397 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_407 ();
 DECAPx10_ASAP7_75t_R FILLER_115_418 ();
 FILLER_ASAP7_75t_R FILLER_115_447 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_455 ();
 FILLER_ASAP7_75t_R FILLER_115_468 ();
 DECAPx6_ASAP7_75t_R FILLER_115_482 ();
 DECAPx1_ASAP7_75t_R FILLER_115_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_500 ();
 FILLER_ASAP7_75t_R FILLER_115_504 ();
 DECAPx1_ASAP7_75t_R FILLER_115_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_516 ();
 DECAPx1_ASAP7_75t_R FILLER_115_523 ();
 FILLER_ASAP7_75t_R FILLER_115_534 ();
 DECAPx2_ASAP7_75t_R FILLER_115_542 ();
 DECAPx2_ASAP7_75t_R FILLER_115_554 ();
 FILLER_ASAP7_75t_R FILLER_115_566 ();
 DECAPx2_ASAP7_75t_R FILLER_115_576 ();
 FILLER_ASAP7_75t_R FILLER_115_590 ();
 FILLER_ASAP7_75t_R FILLER_115_598 ();
 DECAPx10_ASAP7_75t_R FILLER_115_606 ();
 DECAPx6_ASAP7_75t_R FILLER_115_628 ();
 DECAPx2_ASAP7_75t_R FILLER_115_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_648 ();
 FILLER_ASAP7_75t_R FILLER_115_657 ();
 DECAPx6_ASAP7_75t_R FILLER_115_665 ();
 DECAPx10_ASAP7_75t_R FILLER_115_685 ();
 DECAPx10_ASAP7_75t_R FILLER_115_707 ();
 DECAPx4_ASAP7_75t_R FILLER_115_729 ();
 FILLER_ASAP7_75t_R FILLER_115_739 ();
 DECAPx10_ASAP7_75t_R FILLER_115_744 ();
 DECAPx6_ASAP7_75t_R FILLER_115_766 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_780 ();
 DECAPx4_ASAP7_75t_R FILLER_115_789 ();
 FILLER_ASAP7_75t_R FILLER_115_807 ();
 FILLER_ASAP7_75t_R FILLER_115_816 ();
 FILLER_ASAP7_75t_R FILLER_115_821 ();
 DECAPx2_ASAP7_75t_R FILLER_115_829 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_835 ();
 FILLER_ASAP7_75t_R FILLER_115_841 ();
 FILLER_ASAP7_75t_R FILLER_115_852 ();
 DECAPx6_ASAP7_75t_R FILLER_115_862 ();
 FILLER_ASAP7_75t_R FILLER_115_879 ();
 FILLER_ASAP7_75t_R FILLER_115_890 ();
 DECAPx2_ASAP7_75t_R FILLER_115_898 ();
 DECAPx2_ASAP7_75t_R FILLER_115_916 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_922 ();
 DECAPx10_ASAP7_75t_R FILLER_115_927 ();
 DECAPx10_ASAP7_75t_R FILLER_115_949 ();
 DECAPx6_ASAP7_75t_R FILLER_115_971 ();
 DECAPx2_ASAP7_75t_R FILLER_115_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_991 ();
 DECAPx1_ASAP7_75t_R FILLER_115_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1004 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1035 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1054 ();
 FILLER_ASAP7_75t_R FILLER_115_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_115_1087 ();
 FILLER_ASAP7_75t_R FILLER_115_1101 ();
 FILLER_ASAP7_75t_R FILLER_115_1129 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_1139 ();
 FILLER_ASAP7_75t_R FILLER_115_1145 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1153 ();
 FILLER_ASAP7_75t_R FILLER_115_1159 ();
 FILLER_ASAP7_75t_R FILLER_115_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1198 ();
 FILLER_ASAP7_75t_R FILLER_115_1207 ();
 FILLER_ASAP7_75t_R FILLER_115_1218 ();
 DECAPx4_ASAP7_75t_R FILLER_115_1226 ();
 DECAPx2_ASAP7_75t_R FILLER_115_1244 ();
 FILLER_ASAP7_75t_R FILLER_115_1250 ();
 FILLER_ASAP7_75t_R FILLER_115_1260 ();
 FILLER_ASAP7_75t_R FILLER_115_1268 ();
 FILLER_ASAP7_75t_R FILLER_115_1273 ();
 FILLER_ASAP7_75t_R FILLER_115_1284 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_1292 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_1304 ();
 DECAPx6_ASAP7_75t_R FILLER_115_1310 ();
 DECAPx1_ASAP7_75t_R FILLER_115_1334 ();
 DECAPx1_ASAP7_75t_R FILLER_115_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_1348 ();
 FILLER_ASAP7_75t_R FILLER_115_1375 ();
 FILLER_ASAP7_75t_R FILLER_116_2 ();
 DECAPx10_ASAP7_75t_R FILLER_116_30 ();
 DECAPx2_ASAP7_75t_R FILLER_116_52 ();
 FILLER_ASAP7_75t_R FILLER_116_64 ();
 DECAPx2_ASAP7_75t_R FILLER_116_92 ();
 FILLER_ASAP7_75t_R FILLER_116_104 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_109 ();
 DECAPx10_ASAP7_75t_R FILLER_116_118 ();
 FILLER_ASAP7_75t_R FILLER_116_140 ();
 FILLER_ASAP7_75t_R FILLER_116_148 ();
 DECAPx1_ASAP7_75t_R FILLER_116_153 ();
 FILLER_ASAP7_75t_R FILLER_116_183 ();
 FILLER_ASAP7_75t_R FILLER_116_211 ();
 DECAPx4_ASAP7_75t_R FILLER_116_219 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_229 ();
 DECAPx1_ASAP7_75t_R FILLER_116_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_242 ();
 DECAPx6_ASAP7_75t_R FILLER_116_249 ();
 DECAPx2_ASAP7_75t_R FILLER_116_263 ();
 DECAPx6_ASAP7_75t_R FILLER_116_275 ();
 DECAPx1_ASAP7_75t_R FILLER_116_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_293 ();
 FILLER_ASAP7_75t_R FILLER_116_300 ();
 DECAPx2_ASAP7_75t_R FILLER_116_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_311 ();
 FILLER_ASAP7_75t_R FILLER_116_318 ();
 DECAPx4_ASAP7_75t_R FILLER_116_328 ();
 FILLER_ASAP7_75t_R FILLER_116_338 ();
 DECAPx2_ASAP7_75t_R FILLER_116_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_352 ();
 DECAPx1_ASAP7_75t_R FILLER_116_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_363 ();
 DECAPx2_ASAP7_75t_R FILLER_116_367 ();
 DECAPx4_ASAP7_75t_R FILLER_116_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_389 ();
 FILLER_ASAP7_75t_R FILLER_116_396 ();
 DECAPx2_ASAP7_75t_R FILLER_116_409 ();
 FILLER_ASAP7_75t_R FILLER_116_415 ();
 FILLER_ASAP7_75t_R FILLER_116_425 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_433 ();
 DECAPx6_ASAP7_75t_R FILLER_116_443 ();
 DECAPx1_ASAP7_75t_R FILLER_116_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_461 ();
 FILLER_ASAP7_75t_R FILLER_116_464 ();
 DECAPx2_ASAP7_75t_R FILLER_116_476 ();
 DECAPx10_ASAP7_75t_R FILLER_116_488 ();
 DECAPx2_ASAP7_75t_R FILLER_116_510 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_516 ();
 DECAPx2_ASAP7_75t_R FILLER_116_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_533 ();
 DECAPx6_ASAP7_75t_R FILLER_116_542 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_556 ();
 FILLER_ASAP7_75t_R FILLER_116_562 ();
 FILLER_ASAP7_75t_R FILLER_116_586 ();
 DECAPx2_ASAP7_75t_R FILLER_116_594 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_600 ();
 FILLER_ASAP7_75t_R FILLER_116_613 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_621 ();
 DECAPx10_ASAP7_75t_R FILLER_116_632 ();
 DECAPx10_ASAP7_75t_R FILLER_116_654 ();
 DECAPx10_ASAP7_75t_R FILLER_116_684 ();
 DECAPx1_ASAP7_75t_R FILLER_116_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_710 ();
 DECAPx2_ASAP7_75t_R FILLER_116_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_724 ();
 DECAPx1_ASAP7_75t_R FILLER_116_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_736 ();
 FILLER_ASAP7_75t_R FILLER_116_746 ();
 DECAPx2_ASAP7_75t_R FILLER_116_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_769 ();
 DECAPx10_ASAP7_75t_R FILLER_116_781 ();
 DECAPx10_ASAP7_75t_R FILLER_116_810 ();
 DECAPx6_ASAP7_75t_R FILLER_116_832 ();
 DECAPx1_ASAP7_75t_R FILLER_116_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_850 ();
 DECAPx4_ASAP7_75t_R FILLER_116_857 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_867 ();
 FILLER_ASAP7_75t_R FILLER_116_875 ();
 DECAPx10_ASAP7_75t_R FILLER_116_880 ();
 DECAPx2_ASAP7_75t_R FILLER_116_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_908 ();
 DECAPx6_ASAP7_75t_R FILLER_116_915 ();
 FILLER_ASAP7_75t_R FILLER_116_937 ();
 DECAPx2_ASAP7_75t_R FILLER_116_945 ();
 DECAPx10_ASAP7_75t_R FILLER_116_957 ();
 DECAPx4_ASAP7_75t_R FILLER_116_979 ();
 FILLER_ASAP7_75t_R FILLER_116_989 ();
 DECAPx1_ASAP7_75t_R FILLER_116_999 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1026 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_1036 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1047 ();
 FILLER_ASAP7_75t_R FILLER_116_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1071 ();
 FILLER_ASAP7_75t_R FILLER_116_1098 ();
 FILLER_ASAP7_75t_R FILLER_116_1106 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_1114 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_1120 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1129 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_1139 ();
 FILLER_ASAP7_75t_R FILLER_116_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1156 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1173 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1186 ();
 FILLER_ASAP7_75t_R FILLER_116_1197 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1202 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1218 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1228 ();
 FILLER_ASAP7_75t_R FILLER_116_1235 ();
 DECAPx2_ASAP7_75t_R FILLER_116_1246 ();
 DECAPx6_ASAP7_75t_R FILLER_116_1278 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1296 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1304 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1311 ();
 FILLER_ASAP7_75t_R FILLER_116_1321 ();
 DECAPx4_ASAP7_75t_R FILLER_116_1333 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1343 ();
 FILLER_ASAP7_75t_R FILLER_116_1350 ();
 DECAPx1_ASAP7_75t_R FILLER_116_1360 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_1364 ();
 FILLER_ASAP7_75t_R FILLER_116_1368 ();
 FILLER_ASAP7_75t_R FILLER_116_1375 ();
 FILLER_ASAP7_75t_R FILLER_117_2 ();
 FILLER_ASAP7_75t_R FILLER_117_10 ();
 FILLER_ASAP7_75t_R FILLER_117_18 ();
 DECAPx4_ASAP7_75t_R FILLER_117_23 ();
 DECAPx1_ASAP7_75t_R FILLER_117_36 ();
 DECAPx2_ASAP7_75t_R FILLER_117_48 ();
 FILLER_ASAP7_75t_R FILLER_117_54 ();
 DECAPx2_ASAP7_75t_R FILLER_117_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_70 ();
 DECAPx1_ASAP7_75t_R FILLER_117_77 ();
 DECAPx1_ASAP7_75t_R FILLER_117_84 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_94 ();
 DECAPx4_ASAP7_75t_R FILLER_117_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_113 ();
 FILLER_ASAP7_75t_R FILLER_117_120 ();
 DECAPx2_ASAP7_75t_R FILLER_117_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_161 ();
 DECAPx2_ASAP7_75t_R FILLER_117_170 ();
 DECAPx1_ASAP7_75t_R FILLER_117_179 ();
 FILLER_ASAP7_75t_R FILLER_117_189 ();
 FILLER_ASAP7_75t_R FILLER_117_197 ();
 DECAPx1_ASAP7_75t_R FILLER_117_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_206 ();
 FILLER_ASAP7_75t_R FILLER_117_213 ();
 FILLER_ASAP7_75t_R FILLER_117_221 ();
 DECAPx2_ASAP7_75t_R FILLER_117_229 ();
 DECAPx6_ASAP7_75t_R FILLER_117_241 ();
 DECAPx2_ASAP7_75t_R FILLER_117_255 ();
 DECAPx1_ASAP7_75t_R FILLER_117_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_271 ();
 DECAPx10_ASAP7_75t_R FILLER_117_278 ();
 DECAPx4_ASAP7_75t_R FILLER_117_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_316 ();
 DECAPx10_ASAP7_75t_R FILLER_117_323 ();
 DECAPx2_ASAP7_75t_R FILLER_117_345 ();
 FILLER_ASAP7_75t_R FILLER_117_351 ();
 DECAPx4_ASAP7_75t_R FILLER_117_359 ();
 FILLER_ASAP7_75t_R FILLER_117_372 ();
 FILLER_ASAP7_75t_R FILLER_117_382 ();
 DECAPx4_ASAP7_75t_R FILLER_117_399 ();
 FILLER_ASAP7_75t_R FILLER_117_409 ();
 FILLER_ASAP7_75t_R FILLER_117_417 ();
 DECAPx2_ASAP7_75t_R FILLER_117_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_431 ();
 FILLER_ASAP7_75t_R FILLER_117_458 ();
 DECAPx1_ASAP7_75t_R FILLER_117_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_467 ();
 DECAPx1_ASAP7_75t_R FILLER_117_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_475 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_482 ();
 DECAPx10_ASAP7_75t_R FILLER_117_493 ();
 DECAPx6_ASAP7_75t_R FILLER_117_515 ();
 DECAPx2_ASAP7_75t_R FILLER_117_529 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_543 ();
 DECAPx6_ASAP7_75t_R FILLER_117_549 ();
 DECAPx1_ASAP7_75t_R FILLER_117_563 ();
 DECAPx10_ASAP7_75t_R FILLER_117_574 ();
 DECAPx2_ASAP7_75t_R FILLER_117_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_602 ();
 DECAPx6_ASAP7_75t_R FILLER_117_609 ();
 DECAPx2_ASAP7_75t_R FILLER_117_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_645 ();
 FILLER_ASAP7_75t_R FILLER_117_652 ();
 DECAPx2_ASAP7_75t_R FILLER_117_662 ();
 FILLER_ASAP7_75t_R FILLER_117_674 ();
 DECAPx1_ASAP7_75t_R FILLER_117_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_688 ();
 FILLER_ASAP7_75t_R FILLER_117_695 ();
 DECAPx2_ASAP7_75t_R FILLER_117_703 ();
 FILLER_ASAP7_75t_R FILLER_117_717 ();
 FILLER_ASAP7_75t_R FILLER_117_727 ();
 DECAPx2_ASAP7_75t_R FILLER_117_738 ();
 FILLER_ASAP7_75t_R FILLER_117_750 ();
 FILLER_ASAP7_75t_R FILLER_117_763 ();
 FILLER_ASAP7_75t_R FILLER_117_776 ();
 DECAPx6_ASAP7_75t_R FILLER_117_789 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_803 ();
 FILLER_ASAP7_75t_R FILLER_117_815 ();
 FILLER_ASAP7_75t_R FILLER_117_825 ();
 DECAPx2_ASAP7_75t_R FILLER_117_830 ();
 DECAPx2_ASAP7_75t_R FILLER_117_842 ();
 FILLER_ASAP7_75t_R FILLER_117_848 ();
 FILLER_ASAP7_75t_R FILLER_117_859 ();
 FILLER_ASAP7_75t_R FILLER_117_870 ();
 DECAPx2_ASAP7_75t_R FILLER_117_880 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_886 ();
 DECAPx2_ASAP7_75t_R FILLER_117_901 ();
 DECAPx4_ASAP7_75t_R FILLER_117_913 ();
 FILLER_ASAP7_75t_R FILLER_117_923 ();
 FILLER_ASAP7_75t_R FILLER_117_927 ();
 FILLER_ASAP7_75t_R FILLER_117_955 ();
 FILLER_ASAP7_75t_R FILLER_117_967 ();
 FILLER_ASAP7_75t_R FILLER_117_974 ();
 DECAPx6_ASAP7_75t_R FILLER_117_983 ();
 DECAPx2_ASAP7_75t_R FILLER_117_1003 ();
 FILLER_ASAP7_75t_R FILLER_117_1009 ();
 DECAPx6_ASAP7_75t_R FILLER_117_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1033 ();
 FILLER_ASAP7_75t_R FILLER_117_1045 ();
 DECAPx2_ASAP7_75t_R FILLER_117_1053 ();
 FILLER_ASAP7_75t_R FILLER_117_1081 ();
 FILLER_ASAP7_75t_R FILLER_117_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_117_1135 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_1141 ();
 FILLER_ASAP7_75t_R FILLER_117_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_117_1155 ();
 FILLER_ASAP7_75t_R FILLER_117_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1170 ();
 FILLER_ASAP7_75t_R FILLER_117_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_117_1199 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_1209 ();
 FILLER_ASAP7_75t_R FILLER_117_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_117_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1233 ();
 FILLER_ASAP7_75t_R FILLER_117_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1242 ();
 FILLER_ASAP7_75t_R FILLER_117_1264 ();
 DECAPx6_ASAP7_75t_R FILLER_117_1269 ();
 DECAPx2_ASAP7_75t_R FILLER_117_1283 ();
 DECAPx4_ASAP7_75t_R FILLER_117_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_117_1313 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1335 ();
 FILLER_ASAP7_75t_R FILLER_117_1339 ();
 DECAPx1_ASAP7_75t_R FILLER_117_1350 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_1354 ();
 FILLER_ASAP7_75t_R FILLER_117_1361 ();
 FILLER_ASAP7_75t_R FILLER_117_1368 ();
 FILLER_ASAP7_75t_R FILLER_117_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_118_2 ();
 FILLER_ASAP7_75t_R FILLER_118_14 ();
 FILLER_ASAP7_75t_R FILLER_118_22 ();
 DECAPx2_ASAP7_75t_R FILLER_118_29 ();
 FILLER_ASAP7_75t_R FILLER_118_41 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_51 ();
 FILLER_ASAP7_75t_R FILLER_118_62 ();
 DECAPx6_ASAP7_75t_R FILLER_118_70 ();
 DECAPx1_ASAP7_75t_R FILLER_118_110 ();
 FILLER_ASAP7_75t_R FILLER_118_120 ();
 DECAPx2_ASAP7_75t_R FILLER_118_130 ();
 FILLER_ASAP7_75t_R FILLER_118_136 ();
 DECAPx2_ASAP7_75t_R FILLER_118_144 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_150 ();
 DECAPx10_ASAP7_75t_R FILLER_118_159 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_181 ();
 DECAPx1_ASAP7_75t_R FILLER_118_190 ();
 DECAPx6_ASAP7_75t_R FILLER_118_197 ();
 DECAPx1_ASAP7_75t_R FILLER_118_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_215 ();
 DECAPx2_ASAP7_75t_R FILLER_118_242 ();
 FILLER_ASAP7_75t_R FILLER_118_255 ();
 DECAPx2_ASAP7_75t_R FILLER_118_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_289 ();
 DECAPx6_ASAP7_75t_R FILLER_118_316 ();
 DECAPx2_ASAP7_75t_R FILLER_118_337 ();
 FILLER_ASAP7_75t_R FILLER_118_343 ();
 DECAPx4_ASAP7_75t_R FILLER_118_371 ();
 FILLER_ASAP7_75t_R FILLER_118_381 ();
 DECAPx10_ASAP7_75t_R FILLER_118_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_411 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_415 ();
 DECAPx6_ASAP7_75t_R FILLER_118_424 ();
 DECAPx1_ASAP7_75t_R FILLER_118_438 ();
 FILLER_ASAP7_75t_R FILLER_118_448 ();
 DECAPx2_ASAP7_75t_R FILLER_118_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_459 ();
 DECAPx1_ASAP7_75t_R FILLER_118_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_468 ();
 FILLER_ASAP7_75t_R FILLER_118_477 ();
 FILLER_ASAP7_75t_R FILLER_118_487 ();
 FILLER_ASAP7_75t_R FILLER_118_497 ();
 DECAPx4_ASAP7_75t_R FILLER_118_505 ();
 FILLER_ASAP7_75t_R FILLER_118_522 ();
 DECAPx2_ASAP7_75t_R FILLER_118_527 ();
 FILLER_ASAP7_75t_R FILLER_118_539 ();
 FILLER_ASAP7_75t_R FILLER_118_547 ();
 FILLER_ASAP7_75t_R FILLER_118_555 ();
 DECAPx1_ASAP7_75t_R FILLER_118_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_567 ();
 DECAPx2_ASAP7_75t_R FILLER_118_576 ();
 FILLER_ASAP7_75t_R FILLER_118_594 ();
 FILLER_ASAP7_75t_R FILLER_118_606 ();
 FILLER_ASAP7_75t_R FILLER_118_616 ();
 DECAPx2_ASAP7_75t_R FILLER_118_624 ();
 FILLER_ASAP7_75t_R FILLER_118_636 ();
 DECAPx1_ASAP7_75t_R FILLER_118_644 ();
 FILLER_ASAP7_75t_R FILLER_118_654 ();
 DECAPx2_ASAP7_75t_R FILLER_118_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_670 ();
 DECAPx1_ASAP7_75t_R FILLER_118_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_683 ();
 DECAPx2_ASAP7_75t_R FILLER_118_691 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_697 ();
 DECAPx2_ASAP7_75t_R FILLER_118_707 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_713 ();
 DECAPx2_ASAP7_75t_R FILLER_118_722 ();
 DECAPx10_ASAP7_75t_R FILLER_118_734 ();
 DECAPx2_ASAP7_75t_R FILLER_118_756 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_762 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_774 ();
 FILLER_ASAP7_75t_R FILLER_118_785 ();
 DECAPx4_ASAP7_75t_R FILLER_118_799 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_809 ();
 FILLER_ASAP7_75t_R FILLER_118_818 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_829 ();
 FILLER_ASAP7_75t_R FILLER_118_838 ();
 FILLER_ASAP7_75t_R FILLER_118_847 ();
 DECAPx1_ASAP7_75t_R FILLER_118_867 ();
 FILLER_ASAP7_75t_R FILLER_118_881 ();
 DECAPx2_ASAP7_75t_R FILLER_118_901 ();
 FILLER_ASAP7_75t_R FILLER_118_907 ();
 DECAPx4_ASAP7_75t_R FILLER_118_919 ();
 FILLER_ASAP7_75t_R FILLER_118_929 ();
 DECAPx2_ASAP7_75t_R FILLER_118_937 ();
 FILLER_ASAP7_75t_R FILLER_118_946 ();
 FILLER_ASAP7_75t_R FILLER_118_956 ();
 FILLER_ASAP7_75t_R FILLER_118_964 ();
 FILLER_ASAP7_75t_R FILLER_118_972 ();
 DECAPx2_ASAP7_75t_R FILLER_118_982 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_988 ();
 DECAPx4_ASAP7_75t_R FILLER_118_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1011 ();
 FILLER_ASAP7_75t_R FILLER_118_1018 ();
 DECAPx4_ASAP7_75t_R FILLER_118_1026 ();
 FILLER_ASAP7_75t_R FILLER_118_1036 ();
 DECAPx1_ASAP7_75t_R FILLER_118_1044 ();
 FILLER_ASAP7_75t_R FILLER_118_1054 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_1064 ();
 FILLER_ASAP7_75t_R FILLER_118_1074 ();
 FILLER_ASAP7_75t_R FILLER_118_1083 ();
 FILLER_ASAP7_75t_R FILLER_118_1091 ();
 FILLER_ASAP7_75t_R FILLER_118_1099 ();
 DECAPx6_ASAP7_75t_R FILLER_118_1104 ();
 FILLER_ASAP7_75t_R FILLER_118_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_118_1130 ();
 FILLER_ASAP7_75t_R FILLER_118_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_118_1154 ();
 DECAPx6_ASAP7_75t_R FILLER_118_1176 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1196 ();
 DECAPx4_ASAP7_75t_R FILLER_118_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1213 ();
 DECAPx6_ASAP7_75t_R FILLER_118_1220 ();
 DECAPx1_ASAP7_75t_R FILLER_118_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1238 ();
 DECAPx6_ASAP7_75t_R FILLER_118_1245 ();
 FILLER_ASAP7_75t_R FILLER_118_1259 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1271 ();
 DECAPx4_ASAP7_75t_R FILLER_118_1283 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_1293 ();
 FILLER_ASAP7_75t_R FILLER_118_1302 ();
 DECAPx1_ASAP7_75t_R FILLER_118_1330 ();
 FILLER_ASAP7_75t_R FILLER_118_1354 ();
 DECAPx2_ASAP7_75t_R FILLER_118_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_1369 ();
 FILLER_ASAP7_75t_R FILLER_118_1375 ();
 DECAPx1_ASAP7_75t_R FILLER_119_2 ();
 DECAPx1_ASAP7_75t_R FILLER_119_32 ();
 DECAPx4_ASAP7_75t_R FILLER_119_42 ();
 FILLER_ASAP7_75t_R FILLER_119_52 ();
 DECAPx10_ASAP7_75t_R FILLER_119_60 ();
 DECAPx6_ASAP7_75t_R FILLER_119_82 ();
 FILLER_ASAP7_75t_R FILLER_119_96 ();
 DECAPx6_ASAP7_75t_R FILLER_119_101 ();
 DECAPx2_ASAP7_75t_R FILLER_119_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_121 ();
 DECAPx2_ASAP7_75t_R FILLER_119_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_131 ();
 DECAPx4_ASAP7_75t_R FILLER_119_138 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_148 ();
 DECAPx1_ASAP7_75t_R FILLER_119_159 ();
 FILLER_ASAP7_75t_R FILLER_119_169 ();
 FILLER_ASAP7_75t_R FILLER_119_177 ();
 DECAPx4_ASAP7_75t_R FILLER_119_205 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_215 ();
 FILLER_ASAP7_75t_R FILLER_119_224 ();
 FILLER_ASAP7_75t_R FILLER_119_229 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_237 ();
 DECAPx4_ASAP7_75t_R FILLER_119_246 ();
 FILLER_ASAP7_75t_R FILLER_119_256 ();
 DECAPx2_ASAP7_75t_R FILLER_119_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_270 ();
 DECAPx1_ASAP7_75t_R FILLER_119_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_278 ();
 DECAPx4_ASAP7_75t_R FILLER_119_285 ();
 DECAPx1_ASAP7_75t_R FILLER_119_301 ();
 DECAPx1_ASAP7_75t_R FILLER_119_308 ();
 DECAPx2_ASAP7_75t_R FILLER_119_318 ();
 FILLER_ASAP7_75t_R FILLER_119_324 ();
 FILLER_ASAP7_75t_R FILLER_119_332 ();
 DECAPx2_ASAP7_75t_R FILLER_119_342 ();
 DECAPx2_ASAP7_75t_R FILLER_119_354 ();
 DECAPx2_ASAP7_75t_R FILLER_119_363 ();
 FILLER_ASAP7_75t_R FILLER_119_375 ();
 DECAPx2_ASAP7_75t_R FILLER_119_383 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_389 ();
 FILLER_ASAP7_75t_R FILLER_119_418 ();
 DECAPx6_ASAP7_75t_R FILLER_119_442 ();
 DECAPx2_ASAP7_75t_R FILLER_119_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_462 ();
 DECAPx6_ASAP7_75t_R FILLER_119_469 ();
 DECAPx1_ASAP7_75t_R FILLER_119_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_487 ();
 FILLER_ASAP7_75t_R FILLER_119_494 ();
 FILLER_ASAP7_75t_R FILLER_119_504 ();
 FILLER_ASAP7_75t_R FILLER_119_532 ();
 DECAPx2_ASAP7_75t_R FILLER_119_537 ();
 DECAPx2_ASAP7_75t_R FILLER_119_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_556 ();
 DECAPx6_ASAP7_75t_R FILLER_119_569 ();
 DECAPx6_ASAP7_75t_R FILLER_119_588 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_602 ();
 DECAPx1_ASAP7_75t_R FILLER_119_611 ();
 DECAPx1_ASAP7_75t_R FILLER_119_622 ();
 DECAPx2_ASAP7_75t_R FILLER_119_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_635 ();
 DECAPx6_ASAP7_75t_R FILLER_119_642 ();
 DECAPx1_ASAP7_75t_R FILLER_119_656 ();
 DECAPx6_ASAP7_75t_R FILLER_119_667 ();
 FILLER_ASAP7_75t_R FILLER_119_681 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_689 ();
 DECAPx2_ASAP7_75t_R FILLER_119_699 ();
 DECAPx10_ASAP7_75t_R FILLER_119_711 ();
 DECAPx1_ASAP7_75t_R FILLER_119_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_737 ();
 FILLER_ASAP7_75t_R FILLER_119_744 ();
 DECAPx10_ASAP7_75t_R FILLER_119_752 ();
 DECAPx6_ASAP7_75t_R FILLER_119_774 ();
 DECAPx2_ASAP7_75t_R FILLER_119_797 ();
 DECAPx2_ASAP7_75t_R FILLER_119_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_818 ();
 DECAPx2_ASAP7_75t_R FILLER_119_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_831 ();
 FILLER_ASAP7_75t_R FILLER_119_835 ();
 FILLER_ASAP7_75t_R FILLER_119_843 ();
 DECAPx1_ASAP7_75t_R FILLER_119_863 ();
 FILLER_ASAP7_75t_R FILLER_119_873 ();
 FILLER_ASAP7_75t_R FILLER_119_893 ();
 DECAPx2_ASAP7_75t_R FILLER_119_901 ();
 DECAPx4_ASAP7_75t_R FILLER_119_913 ();
 FILLER_ASAP7_75t_R FILLER_119_923 ();
 FILLER_ASAP7_75t_R FILLER_119_927 ();
 FILLER_ASAP7_75t_R FILLER_119_935 ();
 DECAPx10_ASAP7_75t_R FILLER_119_943 ();
 DECAPx2_ASAP7_75t_R FILLER_119_965 ();
 FILLER_ASAP7_75t_R FILLER_119_977 ();
 DECAPx1_ASAP7_75t_R FILLER_119_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_989 ();
 FILLER_ASAP7_75t_R FILLER_119_996 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1033 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_1039 ();
 FILLER_ASAP7_75t_R FILLER_119_1049 ();
 FILLER_ASAP7_75t_R FILLER_119_1061 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1081 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1097 ();
 FILLER_ASAP7_75t_R FILLER_119_1107 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1135 ();
 FILLER_ASAP7_75t_R FILLER_119_1142 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_1154 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_1160 ();
 FILLER_ASAP7_75t_R FILLER_119_1171 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1194 ();
 DECAPx6_ASAP7_75t_R FILLER_119_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1220 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1227 ();
 FILLER_ASAP7_75t_R FILLER_119_1237 ();
 FILLER_ASAP7_75t_R FILLER_119_1265 ();
 FILLER_ASAP7_75t_R FILLER_119_1277 ();
 FILLER_ASAP7_75t_R FILLER_119_1289 ();
 DECAPx2_ASAP7_75t_R FILLER_119_1301 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1313 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_1317 ();
 DECAPx4_ASAP7_75t_R FILLER_119_1321 ();
 FILLER_ASAP7_75t_R FILLER_119_1337 ();
 DECAPx1_ASAP7_75t_R FILLER_119_1345 ();
 FILLER_ASAP7_75t_R FILLER_119_1375 ();
 DECAPx1_ASAP7_75t_R FILLER_120_2 ();
 DECAPx4_ASAP7_75t_R FILLER_120_32 ();
 FILLER_ASAP7_75t_R FILLER_120_42 ();
 FILLER_ASAP7_75t_R FILLER_120_50 ();
 DECAPx6_ASAP7_75t_R FILLER_120_55 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_120_69 ();
 FILLER_ASAP7_75t_R FILLER_120_78 ();
 DECAPx6_ASAP7_75t_R FILLER_120_86 ();
 FILLER_ASAP7_75t_R FILLER_120_100 ();
 FILLER_ASAP7_75t_R FILLER_120_108 ();
 DECAPx6_ASAP7_75t_R FILLER_120_116 ();
 FILLER_ASAP7_75t_R FILLER_120_130 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_120_138 ();
 FILLER_ASAP7_75t_R FILLER_120_147 ();
 DECAPx1_ASAP7_75t_R FILLER_120_155 ();
 DECAPx2_ASAP7_75t_R FILLER_120_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_191 ();
 FILLER_ASAP7_75t_R FILLER_120_198 ();
 DECAPx2_ASAP7_75t_R FILLER_120_226 ();
 FILLER_ASAP7_75t_R FILLER_120_232 ();
 DECAPx10_ASAP7_75t_R FILLER_120_240 ();
 DECAPx2_ASAP7_75t_R FILLER_120_262 ();
 FILLER_ASAP7_75t_R FILLER_120_274 ();
 FILLER_ASAP7_75t_R FILLER_120_302 ();
 FILLER_ASAP7_75t_R FILLER_120_330 ();
 DECAPx10_ASAP7_75t_R FILLER_120_338 ();
 DECAPx1_ASAP7_75t_R FILLER_120_360 ();
 DECAPx2_ASAP7_75t_R FILLER_120_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_376 ();
 DECAPx4_ASAP7_75t_R FILLER_120_380 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_120_390 ();
 FILLER_ASAP7_75t_R FILLER_120_399 ();
 FILLER_ASAP7_75t_R FILLER_120_407 ();
 FILLER_ASAP7_75t_R FILLER_120_412 ();
 FILLER_ASAP7_75t_R FILLER_120_440 ();
 DECAPx2_ASAP7_75t_R FILLER_120_448 ();
 FILLER_ASAP7_75t_R FILLER_120_460 ();
 FILLER_ASAP7_75t_R FILLER_120_464 ();
 DECAPx10_ASAP7_75t_R FILLER_120_472 ();
 DECAPx10_ASAP7_75t_R FILLER_120_494 ();
 FILLER_ASAP7_75t_R FILLER_120_516 ();
 DECAPx10_ASAP7_75t_R FILLER_120_524 ();
 DECAPx6_ASAP7_75t_R FILLER_120_546 ();
 DECAPx2_ASAP7_75t_R FILLER_120_563 ();
 DECAPx2_ASAP7_75t_R FILLER_120_581 ();
 FILLER_ASAP7_75t_R FILLER_120_587 ();
 DECAPx6_ASAP7_75t_R FILLER_120_596 ();
 DECAPx2_ASAP7_75t_R FILLER_120_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_616 ();
 DECAPx4_ASAP7_75t_R FILLER_120_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_635 ();
 DECAPx2_ASAP7_75t_R FILLER_120_646 ();
 DECAPx4_ASAP7_75t_R FILLER_120_659 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_120_669 ();
 DECAPx2_ASAP7_75t_R FILLER_120_679 ();
 DECAPx1_ASAP7_75t_R FILLER_120_696 ();
 DECAPx6_ASAP7_75t_R FILLER_120_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_720 ();
 DECAPx4_ASAP7_75t_R FILLER_120_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_737 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_120_745 ();
 DECAPx4_ASAP7_75t_R FILLER_120_755 ();
 FILLER_ASAP7_75t_R FILLER_120_765 ();
 DECAPx1_ASAP7_75t_R FILLER_120_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_777 ();
 DECAPx10_ASAP7_75t_R FILLER_120_790 ();
 DECAPx10_ASAP7_75t_R FILLER_120_812 ();
 DECAPx10_ASAP7_75t_R FILLER_120_834 ();
 DECAPx6_ASAP7_75t_R FILLER_120_856 ();
 FILLER_ASAP7_75t_R FILLER_120_870 ();
 DECAPx2_ASAP7_75t_R FILLER_120_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_884 ();
 DECAPx10_ASAP7_75t_R FILLER_120_892 ();
 DECAPx2_ASAP7_75t_R FILLER_120_914 ();
 FILLER_ASAP7_75t_R FILLER_120_926 ();
 DECAPx6_ASAP7_75t_R FILLER_120_938 ();
 FILLER_ASAP7_75t_R FILLER_120_958 ();
 DECAPx10_ASAP7_75t_R FILLER_120_963 ();
 DECAPx10_ASAP7_75t_R FILLER_120_985 ();
 FILLER_ASAP7_75t_R FILLER_120_1035 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_120_1063 ();
 FILLER_ASAP7_75t_R FILLER_120_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_120_1110 ();
 FILLER_ASAP7_75t_R FILLER_120_1119 ();
 FILLER_ASAP7_75t_R FILLER_120_1129 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_120_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_120_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_1240 ();
 FILLER_ASAP7_75t_R FILLER_120_1249 ();
 FILLER_ASAP7_75t_R FILLER_120_1257 ();
 DECAPx4_ASAP7_75t_R FILLER_120_1262 ();
 FILLER_ASAP7_75t_R FILLER_120_1272 ();
 FILLER_ASAP7_75t_R FILLER_120_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_120_1302 ();
 DECAPx4_ASAP7_75t_R FILLER_120_1324 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_120_1334 ();
 DECAPx4_ASAP7_75t_R FILLER_120_1340 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_120_1350 ();
 FILLER_ASAP7_75t_R FILLER_120_1361 ();
 FILLER_ASAP7_75t_R FILLER_120_1369 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_120_1374 ();
 DECAPx1_ASAP7_75t_R FILLER_121_2 ();
 FILLER_ASAP7_75t_R FILLER_121_12 ();
 DECAPx4_ASAP7_75t_R FILLER_121_20 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_56 ();
 FILLER_ASAP7_75t_R FILLER_121_65 ();
 FILLER_ASAP7_75t_R FILLER_121_93 ();
 DECAPx6_ASAP7_75t_R FILLER_121_98 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_112 ();
 DECAPx6_ASAP7_75t_R FILLER_121_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_135 ();
 FILLER_ASAP7_75t_R FILLER_121_146 ();
 FILLER_ASAP7_75t_R FILLER_121_154 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_159 ();
 DECAPx1_ASAP7_75t_R FILLER_121_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_172 ();
 DECAPx10_ASAP7_75t_R FILLER_121_176 ();
 DECAPx1_ASAP7_75t_R FILLER_121_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_202 ();
 DECAPx1_ASAP7_75t_R FILLER_121_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_213 ();
 DECAPx10_ASAP7_75t_R FILLER_121_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_239 ();
 DECAPx1_ASAP7_75t_R FILLER_121_246 ();
 FILLER_ASAP7_75t_R FILLER_121_264 ();
 DECAPx1_ASAP7_75t_R FILLER_121_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_276 ();
 DECAPx2_ASAP7_75t_R FILLER_121_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_289 ();
 DECAPx6_ASAP7_75t_R FILLER_121_293 ();
 DECAPx1_ASAP7_75t_R FILLER_121_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_317 ();
 DECAPx4_ASAP7_75t_R FILLER_121_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_331 ();
 DECAPx6_ASAP7_75t_R FILLER_121_335 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_349 ();
 DECAPx10_ASAP7_75t_R FILLER_121_378 ();
 DECAPx6_ASAP7_75t_R FILLER_121_400 ();
 DECAPx2_ASAP7_75t_R FILLER_121_414 ();
 FILLER_ASAP7_75t_R FILLER_121_426 ();
 FILLER_ASAP7_75t_R FILLER_121_431 ();
 DECAPx1_ASAP7_75t_R FILLER_121_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_463 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_472 ();
 DECAPx2_ASAP7_75t_R FILLER_121_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_488 ();
 DECAPx6_ASAP7_75t_R FILLER_121_495 ();
 DECAPx4_ASAP7_75t_R FILLER_121_516 ();
 FILLER_ASAP7_75t_R FILLER_121_526 ();
 DECAPx4_ASAP7_75t_R FILLER_121_534 ();
 DECAPx4_ASAP7_75t_R FILLER_121_550 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_560 ();
 FILLER_ASAP7_75t_R FILLER_121_573 ();
 DECAPx6_ASAP7_75t_R FILLER_121_585 ();
 DECAPx1_ASAP7_75t_R FILLER_121_599 ();
 FILLER_ASAP7_75t_R FILLER_121_609 ();
 DECAPx6_ASAP7_75t_R FILLER_121_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_631 ();
 DECAPx4_ASAP7_75t_R FILLER_121_638 ();
 DECAPx4_ASAP7_75t_R FILLER_121_662 ();
 FILLER_ASAP7_75t_R FILLER_121_678 ();
 DECAPx4_ASAP7_75t_R FILLER_121_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_696 ();
 DECAPx6_ASAP7_75t_R FILLER_121_703 ();
 DECAPx2_ASAP7_75t_R FILLER_121_717 ();
 DECAPx2_ASAP7_75t_R FILLER_121_729 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_735 ();
 DECAPx2_ASAP7_75t_R FILLER_121_748 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_754 ();
 FILLER_ASAP7_75t_R FILLER_121_760 ();
 FILLER_ASAP7_75t_R FILLER_121_771 ();
 DECAPx10_ASAP7_75t_R FILLER_121_781 ();
 DECAPx6_ASAP7_75t_R FILLER_121_811 ();
 DECAPx2_ASAP7_75t_R FILLER_121_835 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_841 ();
 DECAPx2_ASAP7_75t_R FILLER_121_854 ();
 FILLER_ASAP7_75t_R FILLER_121_863 ();
 FILLER_ASAP7_75t_R FILLER_121_874 ();
 DECAPx1_ASAP7_75t_R FILLER_121_882 ();
 DECAPx2_ASAP7_75t_R FILLER_121_896 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_902 ();
 DECAPx4_ASAP7_75t_R FILLER_121_915 ();
 DECAPx6_ASAP7_75t_R FILLER_121_927 ();
 DECAPx1_ASAP7_75t_R FILLER_121_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_945 ();
 FILLER_ASAP7_75t_R FILLER_121_955 ();
 DECAPx6_ASAP7_75t_R FILLER_121_965 ();
 DECAPx2_ASAP7_75t_R FILLER_121_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_985 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_992 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1000 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_1006 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1016 ();
 FILLER_ASAP7_75t_R FILLER_121_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1043 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1058 ();
 DECAPx6_ASAP7_75t_R FILLER_121_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_121_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1098 ();
 DECAPx4_ASAP7_75t_R FILLER_121_1102 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1145 ();
 DECAPx4_ASAP7_75t_R FILLER_121_1167 ();
 FILLER_ASAP7_75t_R FILLER_121_1177 ();
 FILLER_ASAP7_75t_R FILLER_121_1185 ();
 FILLER_ASAP7_75t_R FILLER_121_1193 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_121_1270 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1292 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_1298 ();
 DECAPx4_ASAP7_75t_R FILLER_121_1311 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_1321 ();
 DECAPx6_ASAP7_75t_R FILLER_121_1325 ();
 DECAPx2_ASAP7_75t_R FILLER_121_1339 ();
 FILLER_ASAP7_75t_R FILLER_121_1350 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_1358 ();
 FILLER_ASAP7_75t_R FILLER_121_1366 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_1374 ();
 FILLER_ASAP7_75t_R FILLER_122_2 ();
 DECAPx4_ASAP7_75t_R FILLER_122_10 ();
 DECAPx6_ASAP7_75t_R FILLER_122_23 ();
 FILLER_ASAP7_75t_R FILLER_122_43 ();
 DECAPx2_ASAP7_75t_R FILLER_122_48 ();
 FILLER_ASAP7_75t_R FILLER_122_54 ();
 FILLER_ASAP7_75t_R FILLER_122_82 ();
 DECAPx4_ASAP7_75t_R FILLER_122_87 ();
 FILLER_ASAP7_75t_R FILLER_122_97 ();
 FILLER_ASAP7_75t_R FILLER_122_107 ();
 FILLER_ASAP7_75t_R FILLER_122_117 ();
 DECAPx10_ASAP7_75t_R FILLER_122_127 ();
 DECAPx10_ASAP7_75t_R FILLER_122_149 ();
 DECAPx4_ASAP7_75t_R FILLER_122_171 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_181 ();
 FILLER_ASAP7_75t_R FILLER_122_190 ();
 DECAPx4_ASAP7_75t_R FILLER_122_195 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_205 ();
 DECAPx1_ASAP7_75t_R FILLER_122_214 ();
 FILLER_ASAP7_75t_R FILLER_122_221 ();
 DECAPx2_ASAP7_75t_R FILLER_122_229 ();
 FILLER_ASAP7_75t_R FILLER_122_235 ();
 FILLER_ASAP7_75t_R FILLER_122_243 ();
 FILLER_ASAP7_75t_R FILLER_122_251 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_259 ();
 DECAPx10_ASAP7_75t_R FILLER_122_268 ();
 DECAPx10_ASAP7_75t_R FILLER_122_290 ();
 DECAPx1_ASAP7_75t_R FILLER_122_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_316 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_323 ();
 DECAPx4_ASAP7_75t_R FILLER_122_332 ();
 FILLER_ASAP7_75t_R FILLER_122_342 ();
 DECAPx2_ASAP7_75t_R FILLER_122_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_356 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_363 ();
 DECAPx4_ASAP7_75t_R FILLER_122_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_379 ();
 DECAPx2_ASAP7_75t_R FILLER_122_388 ();
 FILLER_ASAP7_75t_R FILLER_122_394 ();
 FILLER_ASAP7_75t_R FILLER_122_402 ();
 DECAPx10_ASAP7_75t_R FILLER_122_407 ();
 DECAPx2_ASAP7_75t_R FILLER_122_429 ();
 FILLER_ASAP7_75t_R FILLER_122_435 ();
 DECAPx1_ASAP7_75t_R FILLER_122_444 ();
 DECAPx2_ASAP7_75t_R FILLER_122_451 ();
 FILLER_ASAP7_75t_R FILLER_122_460 ();
 FILLER_ASAP7_75t_R FILLER_122_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_473 ();
 FILLER_ASAP7_75t_R FILLER_122_482 ();
 FILLER_ASAP7_75t_R FILLER_122_492 ();
 FILLER_ASAP7_75t_R FILLER_122_501 ();
 FILLER_ASAP7_75t_R FILLER_122_529 ();
 DECAPx1_ASAP7_75t_R FILLER_122_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_541 ();
 FILLER_ASAP7_75t_R FILLER_122_552 ();
 DECAPx4_ASAP7_75t_R FILLER_122_560 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_570 ();
 DECAPx6_ASAP7_75t_R FILLER_122_579 ();
 FILLER_ASAP7_75t_R FILLER_122_599 ();
 FILLER_ASAP7_75t_R FILLER_122_609 ();
 FILLER_ASAP7_75t_R FILLER_122_619 ();
 FILLER_ASAP7_75t_R FILLER_122_627 ();
 FILLER_ASAP7_75t_R FILLER_122_635 ();
 DECAPx6_ASAP7_75t_R FILLER_122_657 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_671 ();
 DECAPx6_ASAP7_75t_R FILLER_122_680 ();
 FILLER_ASAP7_75t_R FILLER_122_694 ();
 DECAPx1_ASAP7_75t_R FILLER_122_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_708 ();
 FILLER_ASAP7_75t_R FILLER_122_717 ();
 FILLER_ASAP7_75t_R FILLER_122_727 ();
 DECAPx4_ASAP7_75t_R FILLER_122_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_745 ();
 DECAPx6_ASAP7_75t_R FILLER_122_754 ();
 FILLER_ASAP7_75t_R FILLER_122_774 ();
 DECAPx2_ASAP7_75t_R FILLER_122_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_785 ();
 FILLER_ASAP7_75t_R FILLER_122_789 ();
 FILLER_ASAP7_75t_R FILLER_122_800 ();
 FILLER_ASAP7_75t_R FILLER_122_811 ();
 DECAPx1_ASAP7_75t_R FILLER_122_819 ();
 FILLER_ASAP7_75t_R FILLER_122_833 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_842 ();
 DECAPx1_ASAP7_75t_R FILLER_122_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_861 ();
 FILLER_ASAP7_75t_R FILLER_122_866 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_874 ();
 FILLER_ASAP7_75t_R FILLER_122_887 ();
 FILLER_ASAP7_75t_R FILLER_122_915 ();
 FILLER_ASAP7_75t_R FILLER_122_929 ();
 DECAPx6_ASAP7_75t_R FILLER_122_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_948 ();
 FILLER_ASAP7_75t_R FILLER_122_952 ();
 FILLER_ASAP7_75t_R FILLER_122_963 ();
 FILLER_ASAP7_75t_R FILLER_122_975 ();
 DECAPx1_ASAP7_75t_R FILLER_122_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_987 ();
 DECAPx2_ASAP7_75t_R FILLER_122_998 ();
 FILLER_ASAP7_75t_R FILLER_122_1004 ();
 DECAPx6_ASAP7_75t_R FILLER_122_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1054 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1099 ();
 DECAPx1_ASAP7_75t_R FILLER_122_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_122_1128 ();
 FILLER_ASAP7_75t_R FILLER_122_1138 ();
 DECAPx4_ASAP7_75t_R FILLER_122_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_122_1169 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_1191 ();
 DECAPx4_ASAP7_75t_R FILLER_122_1204 ();
 FILLER_ASAP7_75t_R FILLER_122_1214 ();
 DECAPx6_ASAP7_75t_R FILLER_122_1224 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_1238 ();
 DECAPx1_ASAP7_75t_R FILLER_122_1247 ();
 FILLER_ASAP7_75t_R FILLER_122_1259 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1269 ();
 FILLER_ASAP7_75t_R FILLER_122_1275 ();
 DECAPx4_ASAP7_75t_R FILLER_122_1283 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_1293 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_1304 ();
 FILLER_ASAP7_75t_R FILLER_122_1333 ();
 DECAPx2_ASAP7_75t_R FILLER_122_1345 ();
 FILLER_ASAP7_75t_R FILLER_122_1359 ();
 FILLER_ASAP7_75t_R FILLER_122_1369 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_1374 ();
 FILLER_ASAP7_75t_R FILLER_123_2 ();
 DECAPx10_ASAP7_75t_R FILLER_123_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_31 ();
 DECAPx10_ASAP7_75t_R FILLER_123_38 ();
 DECAPx1_ASAP7_75t_R FILLER_123_60 ();
 FILLER_ASAP7_75t_R FILLER_123_70 ();
 DECAPx10_ASAP7_75t_R FILLER_123_75 ();
 DECAPx2_ASAP7_75t_R FILLER_123_103 ();
 FILLER_ASAP7_75t_R FILLER_123_109 ();
 FILLER_ASAP7_75t_R FILLER_123_119 ();
 DECAPx10_ASAP7_75t_R FILLER_123_127 ();
 DECAPx2_ASAP7_75t_R FILLER_123_149 ();
 FILLER_ASAP7_75t_R FILLER_123_155 ();
 DECAPx2_ASAP7_75t_R FILLER_123_163 ();
 FILLER_ASAP7_75t_R FILLER_123_169 ();
 DECAPx2_ASAP7_75t_R FILLER_123_197 ();
 FILLER_ASAP7_75t_R FILLER_123_229 ();
 DECAPx10_ASAP7_75t_R FILLER_123_237 ();
 DECAPx2_ASAP7_75t_R FILLER_123_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_265 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_292 ();
 FILLER_ASAP7_75t_R FILLER_123_301 ();
 DECAPx1_ASAP7_75t_R FILLER_123_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_310 ();
 FILLER_ASAP7_75t_R FILLER_123_337 ();
 DECAPx1_ASAP7_75t_R FILLER_123_365 ();
 FILLER_ASAP7_75t_R FILLER_123_372 ();
 FILLER_ASAP7_75t_R FILLER_123_380 ();
 DECAPx2_ASAP7_75t_R FILLER_123_392 ();
 FILLER_ASAP7_75t_R FILLER_123_404 ();
 DECAPx10_ASAP7_75t_R FILLER_123_414 ();
 DECAPx2_ASAP7_75t_R FILLER_123_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_442 ();
 DECAPx10_ASAP7_75t_R FILLER_123_446 ();
 DECAPx6_ASAP7_75t_R FILLER_123_468 ();
 FILLER_ASAP7_75t_R FILLER_123_482 ();
 DECAPx2_ASAP7_75t_R FILLER_123_490 ();
 FILLER_ASAP7_75t_R FILLER_123_496 ();
 DECAPx2_ASAP7_75t_R FILLER_123_505 ();
 DECAPx1_ASAP7_75t_R FILLER_123_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_521 ();
 FILLER_ASAP7_75t_R FILLER_123_525 ();
 DECAPx4_ASAP7_75t_R FILLER_123_535 ();
 FILLER_ASAP7_75t_R FILLER_123_545 ();
 DECAPx2_ASAP7_75t_R FILLER_123_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_560 ();
 DECAPx4_ASAP7_75t_R FILLER_123_569 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_579 ();
 DECAPx1_ASAP7_75t_R FILLER_123_588 ();
 DECAPx2_ASAP7_75t_R FILLER_123_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_610 ();
 DECAPx10_ASAP7_75t_R FILLER_123_617 ();
 DECAPx2_ASAP7_75t_R FILLER_123_639 ();
 FILLER_ASAP7_75t_R FILLER_123_645 ();
 FILLER_ASAP7_75t_R FILLER_123_653 ();
 DECAPx2_ASAP7_75t_R FILLER_123_662 ();
 FILLER_ASAP7_75t_R FILLER_123_668 ();
 FILLER_ASAP7_75t_R FILLER_123_678 ();
 DECAPx1_ASAP7_75t_R FILLER_123_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_692 ();
 FILLER_ASAP7_75t_R FILLER_123_701 ();
 DECAPx1_ASAP7_75t_R FILLER_123_709 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_720 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_731 ();
 DECAPx4_ASAP7_75t_R FILLER_123_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_750 ();
 DECAPx10_ASAP7_75t_R FILLER_123_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_780 ();
 FILLER_ASAP7_75t_R FILLER_123_787 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_795 ();
 FILLER_ASAP7_75t_R FILLER_123_804 ();
 DECAPx1_ASAP7_75t_R FILLER_123_809 ();
 FILLER_ASAP7_75t_R FILLER_123_823 ();
 DECAPx6_ASAP7_75t_R FILLER_123_832 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_846 ();
 DECAPx6_ASAP7_75t_R FILLER_123_852 ();
 FILLER_ASAP7_75t_R FILLER_123_866 ();
 DECAPx6_ASAP7_75t_R FILLER_123_876 ();
 DECAPx1_ASAP7_75t_R FILLER_123_890 ();
 FILLER_ASAP7_75t_R FILLER_123_900 ();
 FILLER_ASAP7_75t_R FILLER_123_908 ();
 DECAPx4_ASAP7_75t_R FILLER_123_913 ();
 FILLER_ASAP7_75t_R FILLER_123_923 ();
 FILLER_ASAP7_75t_R FILLER_123_927 ();
 DECAPx1_ASAP7_75t_R FILLER_123_932 ();
 DECAPx6_ASAP7_75t_R FILLER_123_942 ();
 DECAPx1_ASAP7_75t_R FILLER_123_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_960 ();
 FILLER_ASAP7_75t_R FILLER_123_967 ();
 DECAPx1_ASAP7_75t_R FILLER_123_972 ();
 DECAPx2_ASAP7_75t_R FILLER_123_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_985 ();
 DECAPx6_ASAP7_75t_R FILLER_123_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_123_1017 ();
 FILLER_ASAP7_75t_R FILLER_123_1027 ();
 FILLER_ASAP7_75t_R FILLER_123_1039 ();
 DECAPx4_ASAP7_75t_R FILLER_123_1047 ();
 DECAPx4_ASAP7_75t_R FILLER_123_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1113 ();
 FILLER_ASAP7_75t_R FILLER_123_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_123_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1148 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_1154 ();
 DECAPx1_ASAP7_75t_R FILLER_123_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1171 ();
 FILLER_ASAP7_75t_R FILLER_123_1175 ();
 FILLER_ASAP7_75t_R FILLER_123_1186 ();
 FILLER_ASAP7_75t_R FILLER_123_1194 ();
 FILLER_ASAP7_75t_R FILLER_123_1199 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1207 ();
 DECAPx1_ASAP7_75t_R FILLER_123_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_1243 ();
 FILLER_ASAP7_75t_R FILLER_123_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_123_1278 ();
 FILLER_ASAP7_75t_R FILLER_123_1292 ();
 FILLER_ASAP7_75t_R FILLER_123_1300 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_1308 ();
 DECAPx2_ASAP7_75t_R FILLER_123_1319 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_1325 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_1338 ();
 FILLER_ASAP7_75t_R FILLER_123_1347 ();
 FILLER_ASAP7_75t_R FILLER_123_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_124_2 ();
 DECAPx2_ASAP7_75t_R FILLER_124_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_22 ();
 DECAPx10_ASAP7_75t_R FILLER_124_49 ();
 DECAPx6_ASAP7_75t_R FILLER_124_71 ();
 DECAPx1_ASAP7_75t_R FILLER_124_85 ();
 DECAPx4_ASAP7_75t_R FILLER_124_95 ();
 FILLER_ASAP7_75t_R FILLER_124_105 ();
 DECAPx4_ASAP7_75t_R FILLER_124_113 ();
 FILLER_ASAP7_75t_R FILLER_124_126 ();
 DECAPx1_ASAP7_75t_R FILLER_124_134 ();
 DECAPx2_ASAP7_75t_R FILLER_124_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_147 ();
 DECAPx1_ASAP7_75t_R FILLER_124_174 ();
 DECAPx1_ASAP7_75t_R FILLER_124_184 ();
 FILLER_ASAP7_75t_R FILLER_124_194 ();
 DECAPx1_ASAP7_75t_R FILLER_124_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_203 ();
 DECAPx4_ASAP7_75t_R FILLER_124_210 ();
 FILLER_ASAP7_75t_R FILLER_124_220 ();
 DECAPx1_ASAP7_75t_R FILLER_124_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_252 ();
 FILLER_ASAP7_75t_R FILLER_124_259 ();
 DECAPx1_ASAP7_75t_R FILLER_124_267 ();
 DECAPx2_ASAP7_75t_R FILLER_124_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_283 ();
 DECAPx6_ASAP7_75t_R FILLER_124_310 ();
 FILLER_ASAP7_75t_R FILLER_124_324 ();
 DECAPx4_ASAP7_75t_R FILLER_124_329 ();
 FILLER_ASAP7_75t_R FILLER_124_339 ();
 DECAPx2_ASAP7_75t_R FILLER_124_347 ();
 DECAPx6_ASAP7_75t_R FILLER_124_356 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_370 ();
 FILLER_ASAP7_75t_R FILLER_124_379 ();
 DECAPx6_ASAP7_75t_R FILLER_124_387 ();
 DECAPx1_ASAP7_75t_R FILLER_124_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_405 ();
 FILLER_ASAP7_75t_R FILLER_124_412 ();
 DECAPx2_ASAP7_75t_R FILLER_124_420 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_426 ();
 FILLER_ASAP7_75t_R FILLER_124_455 ();
 FILLER_ASAP7_75t_R FILLER_124_460 ();
 DECAPx6_ASAP7_75t_R FILLER_124_464 ();
 FILLER_ASAP7_75t_R FILLER_124_478 ();
 DECAPx10_ASAP7_75t_R FILLER_124_487 ();
 DECAPx2_ASAP7_75t_R FILLER_124_509 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_515 ();
 DECAPx2_ASAP7_75t_R FILLER_124_521 ();
 FILLER_ASAP7_75t_R FILLER_124_527 ();
 DECAPx2_ASAP7_75t_R FILLER_124_536 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_542 ();
 FILLER_ASAP7_75t_R FILLER_124_552 ();
 FILLER_ASAP7_75t_R FILLER_124_560 ();
 DECAPx1_ASAP7_75t_R FILLER_124_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_578 ();
 DECAPx10_ASAP7_75t_R FILLER_124_586 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_608 ();
 DECAPx4_ASAP7_75t_R FILLER_124_618 ();
 FILLER_ASAP7_75t_R FILLER_124_638 ();
 DECAPx2_ASAP7_75t_R FILLER_124_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_652 ();
 DECAPx10_ASAP7_75t_R FILLER_124_659 ();
 DECAPx2_ASAP7_75t_R FILLER_124_681 ();
 FILLER_ASAP7_75t_R FILLER_124_687 ();
 DECAPx2_ASAP7_75t_R FILLER_124_697 ();
 DECAPx4_ASAP7_75t_R FILLER_124_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_719 ();
 DECAPx1_ASAP7_75t_R FILLER_124_728 ();
 FILLER_ASAP7_75t_R FILLER_124_750 ();
 DECAPx1_ASAP7_75t_R FILLER_124_759 ();
 DECAPx1_ASAP7_75t_R FILLER_124_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_774 ();
 DECAPx10_ASAP7_75t_R FILLER_124_781 ();
 DECAPx10_ASAP7_75t_R FILLER_124_803 ();
 DECAPx6_ASAP7_75t_R FILLER_124_825 ();
 FILLER_ASAP7_75t_R FILLER_124_839 ();
 DECAPx1_ASAP7_75t_R FILLER_124_844 ();
 DECAPx10_ASAP7_75t_R FILLER_124_851 ();
 DECAPx4_ASAP7_75t_R FILLER_124_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_883 ();
 DECAPx2_ASAP7_75t_R FILLER_124_890 ();
 FILLER_ASAP7_75t_R FILLER_124_896 ();
 DECAPx6_ASAP7_75t_R FILLER_124_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_920 ();
 FILLER_ASAP7_75t_R FILLER_124_931 ();
 DECAPx10_ASAP7_75t_R FILLER_124_959 ();
 DECAPx10_ASAP7_75t_R FILLER_124_981 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_1003 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1022 ();
 FILLER_ASAP7_75t_R FILLER_124_1029 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1037 ();
 FILLER_ASAP7_75t_R FILLER_124_1047 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1052 ();
 FILLER_ASAP7_75t_R FILLER_124_1062 ();
 FILLER_ASAP7_75t_R FILLER_124_1072 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_1077 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_1083 ();
 FILLER_ASAP7_75t_R FILLER_124_1094 ();
 FILLER_ASAP7_75t_R FILLER_124_1122 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1133 ();
 FILLER_ASAP7_75t_R FILLER_124_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1191 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_1197 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1207 ();
 FILLER_ASAP7_75t_R FILLER_124_1223 ();
 FILLER_ASAP7_75t_R FILLER_124_1231 ();
 DECAPx6_ASAP7_75t_R FILLER_124_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1250 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_1263 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1274 ();
 FILLER_ASAP7_75t_R FILLER_124_1290 ();
 DECAPx2_ASAP7_75t_R FILLER_124_1301 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_1307 ();
 DECAPx4_ASAP7_75t_R FILLER_124_1336 ();
 DECAPx6_ASAP7_75t_R FILLER_124_1352 ();
 DECAPx1_ASAP7_75t_R FILLER_124_1366 ();
 FILLER_ASAP7_75t_R FILLER_124_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_125_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_24 ();
 DECAPx1_ASAP7_75t_R FILLER_125_33 ();
 DECAPx2_ASAP7_75t_R FILLER_125_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_46 ();
 DECAPx1_ASAP7_75t_R FILLER_125_53 ();
 FILLER_ASAP7_75t_R FILLER_125_63 ();
 FILLER_ASAP7_75t_R FILLER_125_71 ();
 DECAPx1_ASAP7_75t_R FILLER_125_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_80 ();
 DECAPx2_ASAP7_75t_R FILLER_125_107 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_113 ();
 FILLER_ASAP7_75t_R FILLER_125_122 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_150 ();
 DECAPx1_ASAP7_75t_R FILLER_125_159 ();
 DECAPx10_ASAP7_75t_R FILLER_125_166 ();
 DECAPx2_ASAP7_75t_R FILLER_125_194 ();
 FILLER_ASAP7_75t_R FILLER_125_200 ();
 DECAPx6_ASAP7_75t_R FILLER_125_208 ();
 DECAPx1_ASAP7_75t_R FILLER_125_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_226 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_233 ();
 DECAPx2_ASAP7_75t_R FILLER_125_239 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_245 ();
 DECAPx1_ASAP7_75t_R FILLER_125_274 ();
 DECAPx1_ASAP7_75t_R FILLER_125_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_288 ();
 DECAPx1_ASAP7_75t_R FILLER_125_295 ();
 FILLER_ASAP7_75t_R FILLER_125_302 ();
 DECAPx2_ASAP7_75t_R FILLER_125_310 ();
 FILLER_ASAP7_75t_R FILLER_125_316 ();
 DECAPx1_ASAP7_75t_R FILLER_125_324 ();
 DECAPx10_ASAP7_75t_R FILLER_125_331 ();
 DECAPx1_ASAP7_75t_R FILLER_125_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_357 ();
 FILLER_ASAP7_75t_R FILLER_125_364 ();
 DECAPx4_ASAP7_75t_R FILLER_125_369 ();
 FILLER_ASAP7_75t_R FILLER_125_379 ();
 DECAPx2_ASAP7_75t_R FILLER_125_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_413 ();
 DECAPx4_ASAP7_75t_R FILLER_125_420 ();
 FILLER_ASAP7_75t_R FILLER_125_430 ();
 FILLER_ASAP7_75t_R FILLER_125_439 ();
 DECAPx2_ASAP7_75t_R FILLER_125_447 ();
 FILLER_ASAP7_75t_R FILLER_125_463 ();
 DECAPx6_ASAP7_75t_R FILLER_125_475 ();
 DECAPx1_ASAP7_75t_R FILLER_125_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_493 ();
 DECAPx4_ASAP7_75t_R FILLER_125_501 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_519 ();
 DECAPx6_ASAP7_75t_R FILLER_125_528 ();
 DECAPx1_ASAP7_75t_R FILLER_125_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_546 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_555 ();
 DECAPx4_ASAP7_75t_R FILLER_125_564 ();
 FILLER_ASAP7_75t_R FILLER_125_574 ();
 DECAPx2_ASAP7_75t_R FILLER_125_584 ();
 FILLER_ASAP7_75t_R FILLER_125_590 ();
 FILLER_ASAP7_75t_R FILLER_125_600 ();
 DECAPx6_ASAP7_75t_R FILLER_125_608 ();
 FILLER_ASAP7_75t_R FILLER_125_622 ();
 FILLER_ASAP7_75t_R FILLER_125_630 ();
 FILLER_ASAP7_75t_R FILLER_125_638 ();
 FILLER_ASAP7_75t_R FILLER_125_660 ();
 DECAPx10_ASAP7_75t_R FILLER_125_668 ();
 DECAPx10_ASAP7_75t_R FILLER_125_690 ();
 DECAPx4_ASAP7_75t_R FILLER_125_712 ();
 FILLER_ASAP7_75t_R FILLER_125_722 ();
 DECAPx10_ASAP7_75t_R FILLER_125_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_764 ();
 DECAPx10_ASAP7_75t_R FILLER_125_777 ();
 DECAPx2_ASAP7_75t_R FILLER_125_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_805 ();
 DECAPx4_ASAP7_75t_R FILLER_125_812 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_822 ();
 DECAPx1_ASAP7_75t_R FILLER_125_835 ();
 FILLER_ASAP7_75t_R FILLER_125_848 ();
 DECAPx4_ASAP7_75t_R FILLER_125_856 ();
 DECAPx2_ASAP7_75t_R FILLER_125_869 ();
 FILLER_ASAP7_75t_R FILLER_125_875 ();
 FILLER_ASAP7_75t_R FILLER_125_883 ();
 DECAPx2_ASAP7_75t_R FILLER_125_895 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_901 ();
 DECAPx4_ASAP7_75t_R FILLER_125_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_922 ();
 FILLER_ASAP7_75t_R FILLER_125_927 ();
 FILLER_ASAP7_75t_R FILLER_125_936 ();
 FILLER_ASAP7_75t_R FILLER_125_944 ();
 FILLER_ASAP7_75t_R FILLER_125_949 ();
 FILLER_ASAP7_75t_R FILLER_125_958 ();
 DECAPx4_ASAP7_75t_R FILLER_125_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_976 ();
 FILLER_ASAP7_75t_R FILLER_125_980 ();
 DECAPx4_ASAP7_75t_R FILLER_125_990 ();
 FILLER_ASAP7_75t_R FILLER_125_1000 ();
 FILLER_ASAP7_75t_R FILLER_125_1008 ();
 DECAPx1_ASAP7_75t_R FILLER_125_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1020 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_1047 ();
 FILLER_ASAP7_75t_R FILLER_125_1058 ();
 DECAPx6_ASAP7_75t_R FILLER_125_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_125_1077 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_1090 ();
 FILLER_ASAP7_75t_R FILLER_125_1099 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1111 ();
 DECAPx4_ASAP7_75t_R FILLER_125_1123 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_1133 ();
 DECAPx4_ASAP7_75t_R FILLER_125_1142 ();
 FILLER_ASAP7_75t_R FILLER_125_1152 ();
 DECAPx6_ASAP7_75t_R FILLER_125_1157 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_1171 ();
 FILLER_ASAP7_75t_R FILLER_125_1180 ();
 FILLER_ASAP7_75t_R FILLER_125_1192 ();
 DECAPx4_ASAP7_75t_R FILLER_125_1202 ();
 DECAPx4_ASAP7_75t_R FILLER_125_1215 ();
 FILLER_ASAP7_75t_R FILLER_125_1225 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1237 ();
 DECAPx6_ASAP7_75t_R FILLER_125_1246 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1269 ();
 FILLER_ASAP7_75t_R FILLER_125_1275 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1283 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_1289 ();
 DECAPx4_ASAP7_75t_R FILLER_125_1295 ();
 FILLER_ASAP7_75t_R FILLER_125_1305 ();
 FILLER_ASAP7_75t_R FILLER_125_1313 ();
 DECAPx1_ASAP7_75t_R FILLER_125_1321 ();
 DECAPx4_ASAP7_75t_R FILLER_125_1328 ();
 FILLER_ASAP7_75t_R FILLER_125_1338 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_1349 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1358 ();
 FILLER_ASAP7_75t_R FILLER_125_1364 ();
 DECAPx2_ASAP7_75t_R FILLER_125_1369 ();
 FILLER_ASAP7_75t_R FILLER_125_1375 ();
 FILLER_ASAP7_75t_R FILLER_126_2 ();
 DECAPx4_ASAP7_75t_R FILLER_126_10 ();
 FILLER_ASAP7_75t_R FILLER_126_20 ();
 DECAPx4_ASAP7_75t_R FILLER_126_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_38 ();
 DECAPx1_ASAP7_75t_R FILLER_126_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_69 ();
 DECAPx2_ASAP7_75t_R FILLER_126_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_84 ();
 DECAPx1_ASAP7_75t_R FILLER_126_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_95 ();
 DECAPx6_ASAP7_75t_R FILLER_126_99 ();
 FILLER_ASAP7_75t_R FILLER_126_113 ();
 DECAPx4_ASAP7_75t_R FILLER_126_121 ();
 FILLER_ASAP7_75t_R FILLER_126_131 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_155 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_164 ();
 DECAPx4_ASAP7_75t_R FILLER_126_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_183 ();
 DECAPx1_ASAP7_75t_R FILLER_126_192 ();
 FILLER_ASAP7_75t_R FILLER_126_222 ();
 DECAPx4_ASAP7_75t_R FILLER_126_250 ();
 FILLER_ASAP7_75t_R FILLER_126_260 ();
 DECAPx6_ASAP7_75t_R FILLER_126_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_279 ();
 DECAPx10_ASAP7_75t_R FILLER_126_283 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_311 ();
 FILLER_ASAP7_75t_R FILLER_126_340 ();
 FILLER_ASAP7_75t_R FILLER_126_348 ();
 DECAPx4_ASAP7_75t_R FILLER_126_376 ();
 FILLER_ASAP7_75t_R FILLER_126_392 ();
 FILLER_ASAP7_75t_R FILLER_126_400 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_428 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_438 ();
 DECAPx1_ASAP7_75t_R FILLER_126_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_448 ();
 FILLER_ASAP7_75t_R FILLER_126_452 ();
 FILLER_ASAP7_75t_R FILLER_126_460 ();
 DECAPx1_ASAP7_75t_R FILLER_126_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_468 ();
 DECAPx2_ASAP7_75t_R FILLER_126_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_487 ();
 FILLER_ASAP7_75t_R FILLER_126_514 ();
 FILLER_ASAP7_75t_R FILLER_126_522 ();
 FILLER_ASAP7_75t_R FILLER_126_532 ();
 FILLER_ASAP7_75t_R FILLER_126_541 ();
 DECAPx4_ASAP7_75t_R FILLER_126_549 ();
 DECAPx6_ASAP7_75t_R FILLER_126_565 ();
 DECAPx1_ASAP7_75t_R FILLER_126_579 ();
 DECAPx1_ASAP7_75t_R FILLER_126_589 ();
 FILLER_ASAP7_75t_R FILLER_126_601 ();
 DECAPx4_ASAP7_75t_R FILLER_126_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_621 ();
 DECAPx4_ASAP7_75t_R FILLER_126_628 ();
 DECAPx2_ASAP7_75t_R FILLER_126_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_650 ();
 FILLER_ASAP7_75t_R FILLER_126_657 ();
 DECAPx2_ASAP7_75t_R FILLER_126_667 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_673 ();
 FILLER_ASAP7_75t_R FILLER_126_683 ();
 DECAPx1_ASAP7_75t_R FILLER_126_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_695 ();
 FILLER_ASAP7_75t_R FILLER_126_702 ();
 FILLER_ASAP7_75t_R FILLER_126_710 ();
 DECAPx2_ASAP7_75t_R FILLER_126_718 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_724 ();
 FILLER_ASAP7_75t_R FILLER_126_735 ();
 FILLER_ASAP7_75t_R FILLER_126_743 ();
 DECAPx4_ASAP7_75t_R FILLER_126_751 ();
 DECAPx2_ASAP7_75t_R FILLER_126_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_773 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_784 ();
 FILLER_ASAP7_75t_R FILLER_126_799 ();
 FILLER_ASAP7_75t_R FILLER_126_813 ();
 FILLER_ASAP7_75t_R FILLER_126_823 ();
 FILLER_ASAP7_75t_R FILLER_126_831 ();
 DECAPx2_ASAP7_75t_R FILLER_126_839 ();
 DECAPx2_ASAP7_75t_R FILLER_126_853 ();
 FILLER_ASAP7_75t_R FILLER_126_859 ();
 FILLER_ASAP7_75t_R FILLER_126_870 ();
 DECAPx2_ASAP7_75t_R FILLER_126_878 ();
 DECAPx2_ASAP7_75t_R FILLER_126_896 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_902 ();
 FILLER_ASAP7_75t_R FILLER_126_925 ();
 DECAPx4_ASAP7_75t_R FILLER_126_935 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_945 ();
 FILLER_ASAP7_75t_R FILLER_126_952 ();
 DECAPx2_ASAP7_75t_R FILLER_126_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_966 ();
 FILLER_ASAP7_75t_R FILLER_126_970 ();
 FILLER_ASAP7_75t_R FILLER_126_981 ();
 FILLER_ASAP7_75t_R FILLER_126_992 ();
 FILLER_ASAP7_75t_R FILLER_126_1000 ();
 DECAPx4_ASAP7_75t_R FILLER_126_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1016 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1055 ();
 FILLER_ASAP7_75t_R FILLER_126_1068 ();
 DECAPx4_ASAP7_75t_R FILLER_126_1073 ();
 FILLER_ASAP7_75t_R FILLER_126_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1154 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1176 ();
 FILLER_ASAP7_75t_R FILLER_126_1206 ();
 FILLER_ASAP7_75t_R FILLER_126_1211 ();
 FILLER_ASAP7_75t_R FILLER_126_1222 ();
 DECAPx4_ASAP7_75t_R FILLER_126_1227 ();
 FILLER_ASAP7_75t_R FILLER_126_1243 ();
 FILLER_ASAP7_75t_R FILLER_126_1254 ();
 DECAPx4_ASAP7_75t_R FILLER_126_1259 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_1269 ();
 FILLER_ASAP7_75t_R FILLER_126_1278 ();
 FILLER_ASAP7_75t_R FILLER_126_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_126_1297 ();
 DECAPx6_ASAP7_75t_R FILLER_126_1319 ();
 DECAPx1_ASAP7_75t_R FILLER_126_1333 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_1337 ();
 FILLER_ASAP7_75t_R FILLER_126_1347 ();
 FILLER_ASAP7_75t_R FILLER_126_1375 ();
 DECAPx1_ASAP7_75t_R FILLER_127_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_6 ();
 FILLER_ASAP7_75t_R FILLER_127_33 ();
 DECAPx2_ASAP7_75t_R FILLER_127_38 ();
 DECAPx1_ASAP7_75t_R FILLER_127_50 ();
 DECAPx6_ASAP7_75t_R FILLER_127_57 ();
 DECAPx1_ASAP7_75t_R FILLER_127_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_75 ();
 FILLER_ASAP7_75t_R FILLER_127_82 ();
 DECAPx4_ASAP7_75t_R FILLER_127_90 ();
 DECAPx4_ASAP7_75t_R FILLER_127_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_136 ();
 DECAPx1_ASAP7_75t_R FILLER_127_163 ();
 FILLER_ASAP7_75t_R FILLER_127_175 ();
 DECAPx1_ASAP7_75t_R FILLER_127_183 ();
 DECAPx2_ASAP7_75t_R FILLER_127_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_201 ();
 DECAPx1_ASAP7_75t_R FILLER_127_208 ();
 FILLER_ASAP7_75t_R FILLER_127_215 ();
 DECAPx10_ASAP7_75t_R FILLER_127_255 ();
 DECAPx2_ASAP7_75t_R FILLER_127_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_283 ();
 DECAPx4_ASAP7_75t_R FILLER_127_290 ();
 DECAPx2_ASAP7_75t_R FILLER_127_308 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_314 ();
 DECAPx2_ASAP7_75t_R FILLER_127_323 ();
 FILLER_ASAP7_75t_R FILLER_127_329 ();
 FILLER_ASAP7_75t_R FILLER_127_357 ();
 DECAPx2_ASAP7_75t_R FILLER_127_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_371 ();
 DECAPx6_ASAP7_75t_R FILLER_127_378 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_392 ();
 DECAPx4_ASAP7_75t_R FILLER_127_398 ();
 FILLER_ASAP7_75t_R FILLER_127_408 ();
 FILLER_ASAP7_75t_R FILLER_127_416 ();
 DECAPx1_ASAP7_75t_R FILLER_127_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_425 ();
 DECAPx1_ASAP7_75t_R FILLER_127_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_456 ();
 DECAPx1_ASAP7_75t_R FILLER_127_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_467 ();
 DECAPx6_ASAP7_75t_R FILLER_127_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_488 ();
 DECAPx1_ASAP7_75t_R FILLER_127_496 ();
 FILLER_ASAP7_75t_R FILLER_127_506 ();
 DECAPx10_ASAP7_75t_R FILLER_127_511 ();
 DECAPx10_ASAP7_75t_R FILLER_127_533 ();
 FILLER_ASAP7_75t_R FILLER_127_555 ();
 FILLER_ASAP7_75t_R FILLER_127_563 ();
 DECAPx10_ASAP7_75t_R FILLER_127_571 ();
 DECAPx2_ASAP7_75t_R FILLER_127_593 ();
 FILLER_ASAP7_75t_R FILLER_127_599 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_607 ();
 DECAPx2_ASAP7_75t_R FILLER_127_613 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_619 ();
 DECAPx6_ASAP7_75t_R FILLER_127_628 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_642 ();
 DECAPx4_ASAP7_75t_R FILLER_127_653 ();
 FILLER_ASAP7_75t_R FILLER_127_670 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_684 ();
 DECAPx4_ASAP7_75t_R FILLER_127_694 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_712 ();
 DECAPx4_ASAP7_75t_R FILLER_127_722 ();
 DECAPx2_ASAP7_75t_R FILLER_127_739 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_745 ();
 FILLER_ASAP7_75t_R FILLER_127_756 ();
 DECAPx4_ASAP7_75t_R FILLER_127_764 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_774 ();
 DECAPx4_ASAP7_75t_R FILLER_127_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_793 ();
 DECAPx4_ASAP7_75t_R FILLER_127_797 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_807 ();
 DECAPx6_ASAP7_75t_R FILLER_127_820 ();
 DECAPx2_ASAP7_75t_R FILLER_127_834 ();
 FILLER_ASAP7_75t_R FILLER_127_844 ();
 DECAPx6_ASAP7_75t_R FILLER_127_852 ();
 DECAPx2_ASAP7_75t_R FILLER_127_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_880 ();
 DECAPx6_ASAP7_75t_R FILLER_127_887 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_901 ();
 DECAPx4_ASAP7_75t_R FILLER_127_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_922 ();
 DECAPx1_ASAP7_75t_R FILLER_127_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_931 ();
 DECAPx6_ASAP7_75t_R FILLER_127_938 ();
 FILLER_ASAP7_75t_R FILLER_127_952 ();
 DECAPx2_ASAP7_75t_R FILLER_127_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_966 ();
 FILLER_ASAP7_75t_R FILLER_127_989 ();
 DECAPx2_ASAP7_75t_R FILLER_127_997 ();
 FILLER_ASAP7_75t_R FILLER_127_1003 ();
 DECAPx6_ASAP7_75t_R FILLER_127_1011 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1036 ();
 FILLER_ASAP7_75t_R FILLER_127_1052 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_1060 ();
 DECAPx6_ASAP7_75t_R FILLER_127_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1092 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1114 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_1120 ();
 FILLER_ASAP7_75t_R FILLER_127_1131 ();
 DECAPx4_ASAP7_75t_R FILLER_127_1139 ();
 FILLER_ASAP7_75t_R FILLER_127_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_127_1157 ();
 DECAPx4_ASAP7_75t_R FILLER_127_1173 ();
 FILLER_ASAP7_75t_R FILLER_127_1190 ();
 DECAPx4_ASAP7_75t_R FILLER_127_1202 ();
 FILLER_ASAP7_75t_R FILLER_127_1212 ();
 DECAPx4_ASAP7_75t_R FILLER_127_1220 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_1230 ();
 DECAPx6_ASAP7_75t_R FILLER_127_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1259 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1281 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1290 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_1302 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_127_1329 ();
 DECAPx1_ASAP7_75t_R FILLER_127_1351 ();
 DECAPx2_ASAP7_75t_R FILLER_127_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_1369 ();
 FILLER_ASAP7_75t_R FILLER_127_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_128_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_16 ();
 FILLER_ASAP7_75t_R FILLER_128_23 ();
 DECAPx10_ASAP7_75t_R FILLER_128_28 ();
 DECAPx1_ASAP7_75t_R FILLER_128_50 ();
 FILLER_ASAP7_75t_R FILLER_128_60 ();
 FILLER_ASAP7_75t_R FILLER_128_68 ();
 FILLER_ASAP7_75t_R FILLER_128_78 ();
 DECAPx10_ASAP7_75t_R FILLER_128_86 ();
 FILLER_ASAP7_75t_R FILLER_128_114 ();
 DECAPx6_ASAP7_75t_R FILLER_128_119 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_133 ();
 FILLER_ASAP7_75t_R FILLER_128_142 ();
 FILLER_ASAP7_75t_R FILLER_128_150 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_155 ();
 FILLER_ASAP7_75t_R FILLER_128_164 ();
 DECAPx1_ASAP7_75t_R FILLER_128_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_173 ();
 DECAPx10_ASAP7_75t_R FILLER_128_180 ();
 DECAPx10_ASAP7_75t_R FILLER_128_202 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_224 ();
 FILLER_ASAP7_75t_R FILLER_128_233 ();
 FILLER_ASAP7_75t_R FILLER_128_253 ();
 DECAPx2_ASAP7_75t_R FILLER_128_258 ();
 FILLER_ASAP7_75t_R FILLER_128_264 ();
 DECAPx1_ASAP7_75t_R FILLER_128_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_276 ();
 FILLER_ASAP7_75t_R FILLER_128_283 ();
 DECAPx2_ASAP7_75t_R FILLER_128_293 ();
 FILLER_ASAP7_75t_R FILLER_128_307 ();
 DECAPx2_ASAP7_75t_R FILLER_128_331 ();
 FILLER_ASAP7_75t_R FILLER_128_337 ();
 FILLER_ASAP7_75t_R FILLER_128_345 ();
 DECAPx6_ASAP7_75t_R FILLER_128_350 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_364 ();
 DECAPx10_ASAP7_75t_R FILLER_128_393 ();
 DECAPx10_ASAP7_75t_R FILLER_128_415 ();
 FILLER_ASAP7_75t_R FILLER_128_437 ();
 DECAPx6_ASAP7_75t_R FILLER_128_445 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_459 ();
 DECAPx4_ASAP7_75t_R FILLER_128_464 ();
 DECAPx10_ASAP7_75t_R FILLER_128_482 ();
 DECAPx6_ASAP7_75t_R FILLER_128_504 ();
 DECAPx1_ASAP7_75t_R FILLER_128_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_522 ();
 DECAPx1_ASAP7_75t_R FILLER_128_529 ();
 DECAPx1_ASAP7_75t_R FILLER_128_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_540 ();
 DECAPx4_ASAP7_75t_R FILLER_128_548 ();
 FILLER_ASAP7_75t_R FILLER_128_565 ();
 DECAPx2_ASAP7_75t_R FILLER_128_577 ();
 DECAPx2_ASAP7_75t_R FILLER_128_589 ();
 DECAPx4_ASAP7_75t_R FILLER_128_601 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_611 ();
 FILLER_ASAP7_75t_R FILLER_128_620 ();
 DECAPx6_ASAP7_75t_R FILLER_128_632 ();
 DECAPx1_ASAP7_75t_R FILLER_128_646 ();
 DECAPx10_ASAP7_75t_R FILLER_128_656 ();
 DECAPx10_ASAP7_75t_R FILLER_128_678 ();
 FILLER_ASAP7_75t_R FILLER_128_716 ();
 DECAPx1_ASAP7_75t_R FILLER_128_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_730 ();
 DECAPx1_ASAP7_75t_R FILLER_128_737 ();
 DECAPx2_ASAP7_75t_R FILLER_128_751 ();
 FILLER_ASAP7_75t_R FILLER_128_765 ();
 DECAPx6_ASAP7_75t_R FILLER_128_773 ();
 DECAPx6_ASAP7_75t_R FILLER_128_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_808 ();
 DECAPx2_ASAP7_75t_R FILLER_128_819 ();
 FILLER_ASAP7_75t_R FILLER_128_825 ();
 DECAPx4_ASAP7_75t_R FILLER_128_833 ();
 DECAPx6_ASAP7_75t_R FILLER_128_852 ();
 FILLER_ASAP7_75t_R FILLER_128_866 ();
 DECAPx10_ASAP7_75t_R FILLER_128_874 ();
 DECAPx2_ASAP7_75t_R FILLER_128_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_902 ();
 DECAPx2_ASAP7_75t_R FILLER_128_910 ();
 DECAPx4_ASAP7_75t_R FILLER_128_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_929 ();
 FILLER_ASAP7_75t_R FILLER_128_950 ();
 DECAPx2_ASAP7_75t_R FILLER_128_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_984 ();
 DECAPx2_ASAP7_75t_R FILLER_128_993 ();
 FILLER_ASAP7_75t_R FILLER_128_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_128_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_128_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1053 ();
 FILLER_ASAP7_75t_R FILLER_128_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1079 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1090 ();
 FILLER_ASAP7_75t_R FILLER_128_1106 ();
 FILLER_ASAP7_75t_R FILLER_128_1134 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1145 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1178 ();
 DECAPx6_ASAP7_75t_R FILLER_128_1187 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1205 ();
 FILLER_ASAP7_75t_R FILLER_128_1212 ();
 DECAPx6_ASAP7_75t_R FILLER_128_1224 ();
 DECAPx2_ASAP7_75t_R FILLER_128_1238 ();
 FILLER_ASAP7_75t_R FILLER_128_1250 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1266 ();
 DECAPx6_ASAP7_75t_R FILLER_128_1270 ();
 FILLER_ASAP7_75t_R FILLER_128_1287 ();
 DECAPx1_ASAP7_75t_R FILLER_128_1298 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_1302 ();
 FILLER_ASAP7_75t_R FILLER_128_1329 ();
 FILLER_ASAP7_75t_R FILLER_128_1351 ();
 FILLER_ASAP7_75t_R FILLER_128_1361 ();
 FILLER_ASAP7_75t_R FILLER_128_1366 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_1374 ();
 FILLER_ASAP7_75t_R FILLER_129_2 ();
 DECAPx6_ASAP7_75t_R FILLER_129_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_24 ();
 FILLER_ASAP7_75t_R FILLER_129_31 ();
 DECAPx2_ASAP7_75t_R FILLER_129_39 ();
 FILLER_ASAP7_75t_R FILLER_129_45 ();
 FILLER_ASAP7_75t_R FILLER_129_53 ();
 DECAPx10_ASAP7_75t_R FILLER_129_65 ();
 FILLER_ASAP7_75t_R FILLER_129_87 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_97 ();
 DECAPx4_ASAP7_75t_R FILLER_129_106 ();
 FILLER_ASAP7_75t_R FILLER_129_122 ();
 DECAPx10_ASAP7_75t_R FILLER_129_130 ();
 DECAPx6_ASAP7_75t_R FILLER_129_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_166 ();
 FILLER_ASAP7_75t_R FILLER_129_173 ();
 DECAPx2_ASAP7_75t_R FILLER_129_181 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_187 ();
 FILLER_ASAP7_75t_R FILLER_129_196 ();
 DECAPx2_ASAP7_75t_R FILLER_129_204 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_210 ();
 DECAPx1_ASAP7_75t_R FILLER_129_219 ();
 DECAPx2_ASAP7_75t_R FILLER_129_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_232 ();
 FILLER_ASAP7_75t_R FILLER_129_236 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_264 ();
 FILLER_ASAP7_75t_R FILLER_129_275 ();
 FILLER_ASAP7_75t_R FILLER_129_283 ();
 FILLER_ASAP7_75t_R FILLER_129_307 ();
 DECAPx4_ASAP7_75t_R FILLER_129_315 ();
 FILLER_ASAP7_75t_R FILLER_129_331 ();
 DECAPx6_ASAP7_75t_R FILLER_129_336 ();
 DECAPx2_ASAP7_75t_R FILLER_129_350 ();
 DECAPx6_ASAP7_75t_R FILLER_129_362 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_376 ();
 DECAPx2_ASAP7_75t_R FILLER_129_385 ();
 DECAPx1_ASAP7_75t_R FILLER_129_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_398 ();
 FILLER_ASAP7_75t_R FILLER_129_405 ();
 DECAPx1_ASAP7_75t_R FILLER_129_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_437 ();
 DECAPx4_ASAP7_75t_R FILLER_129_444 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_460 ();
 DECAPx1_ASAP7_75t_R FILLER_129_469 ();
 DECAPx6_ASAP7_75t_R FILLER_129_481 ();
 DECAPx6_ASAP7_75t_R FILLER_129_501 ();
 DECAPx1_ASAP7_75t_R FILLER_129_515 ();
 FILLER_ASAP7_75t_R FILLER_129_525 ();
 FILLER_ASAP7_75t_R FILLER_129_533 ();
 DECAPx2_ASAP7_75t_R FILLER_129_543 ();
 FILLER_ASAP7_75t_R FILLER_129_549 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_558 ();
 FILLER_ASAP7_75t_R FILLER_129_573 ();
 FILLER_ASAP7_75t_R FILLER_129_581 ();
 DECAPx2_ASAP7_75t_R FILLER_129_593 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_605 ();
 DECAPx2_ASAP7_75t_R FILLER_129_614 ();
 FILLER_ASAP7_75t_R FILLER_129_620 ();
 DECAPx2_ASAP7_75t_R FILLER_129_632 ();
 DECAPx1_ASAP7_75t_R FILLER_129_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_648 ();
 DECAPx2_ASAP7_75t_R FILLER_129_665 ();
 DECAPx4_ASAP7_75t_R FILLER_129_677 ();
 FILLER_ASAP7_75t_R FILLER_129_687 ();
 DECAPx6_ASAP7_75t_R FILLER_129_696 ();
 DECAPx1_ASAP7_75t_R FILLER_129_710 ();
 DECAPx2_ASAP7_75t_R FILLER_129_721 ();
 FILLER_ASAP7_75t_R FILLER_129_727 ();
 DECAPx6_ASAP7_75t_R FILLER_129_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_749 ();
 DECAPx4_ASAP7_75t_R FILLER_129_757 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_767 ();
 DECAPx6_ASAP7_75t_R FILLER_129_780 ();
 DECAPx2_ASAP7_75t_R FILLER_129_800 ();
 FILLER_ASAP7_75t_R FILLER_129_806 ();
 DECAPx2_ASAP7_75t_R FILLER_129_813 ();
 DECAPx4_ASAP7_75t_R FILLER_129_845 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_855 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_861 ();
 FILLER_ASAP7_75t_R FILLER_129_867 ();
 DECAPx2_ASAP7_75t_R FILLER_129_878 ();
 FILLER_ASAP7_75t_R FILLER_129_884 ();
 DECAPx1_ASAP7_75t_R FILLER_129_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_896 ();
 DECAPx1_ASAP7_75t_R FILLER_129_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_904 ();
 DECAPx2_ASAP7_75t_R FILLER_129_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_917 ();
 FILLER_ASAP7_75t_R FILLER_129_923 ();
 DECAPx2_ASAP7_75t_R FILLER_129_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_933 ();
 DECAPx10_ASAP7_75t_R FILLER_129_941 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_963 ();
 FILLER_ASAP7_75t_R FILLER_129_969 ();
 DECAPx4_ASAP7_75t_R FILLER_129_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_984 ();
 FILLER_ASAP7_75t_R FILLER_129_995 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1006 ();
 FILLER_ASAP7_75t_R FILLER_129_1018 ();
 DECAPx6_ASAP7_75t_R FILLER_129_1030 ();
 DECAPx4_ASAP7_75t_R FILLER_129_1052 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_1062 ();
 DECAPx4_ASAP7_75t_R FILLER_129_1068 ();
 FILLER_ASAP7_75t_R FILLER_129_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1114 ();
 FILLER_ASAP7_75t_R FILLER_129_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1137 ();
 FILLER_ASAP7_75t_R FILLER_129_1147 ();
 FILLER_ASAP7_75t_R FILLER_129_1157 ();
 FILLER_ASAP7_75t_R FILLER_129_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1178 ();
 DECAPx4_ASAP7_75t_R FILLER_129_1205 ();
 DECAPx4_ASAP7_75t_R FILLER_129_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1251 ();
 FILLER_ASAP7_75t_R FILLER_129_1278 ();
 FILLER_ASAP7_75t_R FILLER_129_1290 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1298 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_1304 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1313 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1317 ();
 DECAPx2_ASAP7_75t_R FILLER_129_1321 ();
 FILLER_ASAP7_75t_R FILLER_129_1327 ();
 FILLER_ASAP7_75t_R FILLER_129_1336 ();
 DECAPx1_ASAP7_75t_R FILLER_129_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_1348 ();
 FILLER_ASAP7_75t_R FILLER_129_1375 ();
 FILLER_ASAP7_75t_R FILLER_130_2 ();
 DECAPx4_ASAP7_75t_R FILLER_130_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_19 ();
 DECAPx2_ASAP7_75t_R FILLER_130_46 ();
 DECAPx4_ASAP7_75t_R FILLER_130_58 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_68 ();
 DECAPx2_ASAP7_75t_R FILLER_130_77 ();
 FILLER_ASAP7_75t_R FILLER_130_83 ();
 FILLER_ASAP7_75t_R FILLER_130_91 ();
 DECAPx1_ASAP7_75t_R FILLER_130_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_123 ();
 FILLER_ASAP7_75t_R FILLER_130_132 ();
 FILLER_ASAP7_75t_R FILLER_130_142 ();
 DECAPx2_ASAP7_75t_R FILLER_130_150 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_156 ();
 DECAPx2_ASAP7_75t_R FILLER_130_169 ();
 FILLER_ASAP7_75t_R FILLER_130_175 ();
 DECAPx2_ASAP7_75t_R FILLER_130_184 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_190 ();
 DECAPx2_ASAP7_75t_R FILLER_130_201 ();
 FILLER_ASAP7_75t_R FILLER_130_207 ();
 DECAPx1_ASAP7_75t_R FILLER_130_235 ();
 FILLER_ASAP7_75t_R FILLER_130_245 ();
 FILLER_ASAP7_75t_R FILLER_130_253 ();
 DECAPx1_ASAP7_75t_R FILLER_130_258 ();
 FILLER_ASAP7_75t_R FILLER_130_265 ();
 DECAPx2_ASAP7_75t_R FILLER_130_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_281 ();
 FILLER_ASAP7_75t_R FILLER_130_290 ();
 DECAPx2_ASAP7_75t_R FILLER_130_298 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_311 ();
 DECAPx2_ASAP7_75t_R FILLER_130_340 ();
 FILLER_ASAP7_75t_R FILLER_130_346 ();
 DECAPx2_ASAP7_75t_R FILLER_130_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_380 ();
 DECAPx4_ASAP7_75t_R FILLER_130_384 ();
 FILLER_ASAP7_75t_R FILLER_130_394 ();
 FILLER_ASAP7_75t_R FILLER_130_404 ();
 FILLER_ASAP7_75t_R FILLER_130_412 ();
 DECAPx2_ASAP7_75t_R FILLER_130_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_426 ();
 DECAPx2_ASAP7_75t_R FILLER_130_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_459 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_464 ();
 FILLER_ASAP7_75t_R FILLER_130_473 ();
 FILLER_ASAP7_75t_R FILLER_130_483 ();
 FILLER_ASAP7_75t_R FILLER_130_492 ();
 FILLER_ASAP7_75t_R FILLER_130_502 ();
 DECAPx1_ASAP7_75t_R FILLER_130_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_514 ();
 DECAPx10_ASAP7_75t_R FILLER_130_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_547 ();
 DECAPx10_ASAP7_75t_R FILLER_130_560 ();
 DECAPx4_ASAP7_75t_R FILLER_130_582 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_592 ();
 FILLER_ASAP7_75t_R FILLER_130_610 ();
 DECAPx4_ASAP7_75t_R FILLER_130_622 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_632 ();
 FILLER_ASAP7_75t_R FILLER_130_643 ();
 DECAPx2_ASAP7_75t_R FILLER_130_652 ();
 DECAPx2_ASAP7_75t_R FILLER_130_664 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_670 ();
 DECAPx2_ASAP7_75t_R FILLER_130_680 ();
 DECAPx10_ASAP7_75t_R FILLER_130_696 ();
 DECAPx2_ASAP7_75t_R FILLER_130_718 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_724 ();
 DECAPx10_ASAP7_75t_R FILLER_130_733 ();
 DECAPx1_ASAP7_75t_R FILLER_130_755 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_767 ();
 FILLER_ASAP7_75t_R FILLER_130_777 ();
 FILLER_ASAP7_75t_R FILLER_130_786 ();
 DECAPx1_ASAP7_75t_R FILLER_130_794 ();
 DECAPx6_ASAP7_75t_R FILLER_130_806 ();
 DECAPx1_ASAP7_75t_R FILLER_130_820 ();
 FILLER_ASAP7_75t_R FILLER_130_830 ();
 FILLER_ASAP7_75t_R FILLER_130_835 ();
 DECAPx6_ASAP7_75t_R FILLER_130_840 ();
 FILLER_ASAP7_75t_R FILLER_130_854 ();
 DECAPx6_ASAP7_75t_R FILLER_130_866 ();
 FILLER_ASAP7_75t_R FILLER_130_880 ();
 DECAPx1_ASAP7_75t_R FILLER_130_908 ();
 FILLER_ASAP7_75t_R FILLER_130_926 ();
 DECAPx2_ASAP7_75t_R FILLER_130_934 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_940 ();
 FILLER_ASAP7_75t_R FILLER_130_949 ();
 DECAPx10_ASAP7_75t_R FILLER_130_977 ();
 DECAPx6_ASAP7_75t_R FILLER_130_999 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1024 ();
 FILLER_ASAP7_75t_R FILLER_130_1054 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_1059 ();
 FILLER_ASAP7_75t_R FILLER_130_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1078 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_1084 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1095 ();
 FILLER_ASAP7_75t_R FILLER_130_1101 ();
 DECAPx6_ASAP7_75t_R FILLER_130_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1120 ();
 FILLER_ASAP7_75t_R FILLER_130_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1138 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_1144 ();
 DECAPx6_ASAP7_75t_R FILLER_130_1153 ();
 FILLER_ASAP7_75t_R FILLER_130_1170 ();
 FILLER_ASAP7_75t_R FILLER_130_1181 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1192 ();
 FILLER_ASAP7_75t_R FILLER_130_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1205 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1228 ();
 DECAPx6_ASAP7_75t_R FILLER_130_1232 ();
 DECAPx2_ASAP7_75t_R FILLER_130_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_130_1261 ();
 DECAPx4_ASAP7_75t_R FILLER_130_1283 ();
 DECAPx6_ASAP7_75t_R FILLER_130_1299 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_1313 ();
 FILLER_ASAP7_75t_R FILLER_130_1326 ();
 FILLER_ASAP7_75t_R FILLER_130_1331 ();
 DECAPx1_ASAP7_75t_R FILLER_130_1342 ();
 FILLER_ASAP7_75t_R FILLER_130_1354 ();
 FILLER_ASAP7_75t_R FILLER_130_1361 ();
 FILLER_ASAP7_75t_R FILLER_130_1368 ();
 FILLER_ASAP7_75t_R FILLER_130_1375 ();
 FILLER_ASAP7_75t_R FILLER_131_2 ();
 DECAPx4_ASAP7_75t_R FILLER_131_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_19 ();
 DECAPx1_ASAP7_75t_R FILLER_131_26 ();
 FILLER_ASAP7_75t_R FILLER_131_33 ();
 DECAPx4_ASAP7_75t_R FILLER_131_38 ();
 FILLER_ASAP7_75t_R FILLER_131_48 ();
 FILLER_ASAP7_75t_R FILLER_131_56 ();
 DECAPx2_ASAP7_75t_R FILLER_131_64 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_70 ();
 DECAPx4_ASAP7_75t_R FILLER_131_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_89 ();
 FILLER_ASAP7_75t_R FILLER_131_96 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_104 ();
 FILLER_ASAP7_75t_R FILLER_131_114 ();
 FILLER_ASAP7_75t_R FILLER_131_123 ();
 FILLER_ASAP7_75t_R FILLER_131_131 ();
 DECAPx6_ASAP7_75t_R FILLER_131_139 ();
 DECAPx1_ASAP7_75t_R FILLER_131_153 ();
 DECAPx2_ASAP7_75t_R FILLER_131_171 ();
 FILLER_ASAP7_75t_R FILLER_131_177 ();
 DECAPx2_ASAP7_75t_R FILLER_131_185 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_191 ();
 FILLER_ASAP7_75t_R FILLER_131_202 ();
 FILLER_ASAP7_75t_R FILLER_131_210 ();
 DECAPx10_ASAP7_75t_R FILLER_131_218 ();
 FILLER_ASAP7_75t_R FILLER_131_240 ();
 DECAPx10_ASAP7_75t_R FILLER_131_248 ();
 DECAPx1_ASAP7_75t_R FILLER_131_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_274 ();
 DECAPx4_ASAP7_75t_R FILLER_131_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_291 ();
 DECAPx1_ASAP7_75t_R FILLER_131_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_302 ();
 DECAPx4_ASAP7_75t_R FILLER_131_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_319 ();
 DECAPx2_ASAP7_75t_R FILLER_131_326 ();
 FILLER_ASAP7_75t_R FILLER_131_340 ();
 DECAPx2_ASAP7_75t_R FILLER_131_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_351 ();
 DECAPx1_ASAP7_75t_R FILLER_131_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_362 ();
 DECAPx4_ASAP7_75t_R FILLER_131_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_376 ();
 DECAPx6_ASAP7_75t_R FILLER_131_383 ();
 FILLER_ASAP7_75t_R FILLER_131_397 ();
 DECAPx1_ASAP7_75t_R FILLER_131_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_411 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_418 ();
 DECAPx2_ASAP7_75t_R FILLER_131_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_430 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_438 ();
 DECAPx2_ASAP7_75t_R FILLER_131_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_450 ();
 FILLER_ASAP7_75t_R FILLER_131_454 ();
 FILLER_ASAP7_75t_R FILLER_131_464 ();
 DECAPx1_ASAP7_75t_R FILLER_131_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_476 ();
 DECAPx1_ASAP7_75t_R FILLER_131_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_488 ();
 FILLER_ASAP7_75t_R FILLER_131_495 ();
 DECAPx1_ASAP7_75t_R FILLER_131_503 ();
 DECAPx2_ASAP7_75t_R FILLER_131_514 ();
 DECAPx10_ASAP7_75t_R FILLER_131_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_548 ();
 DECAPx10_ASAP7_75t_R FILLER_131_552 ();
 DECAPx4_ASAP7_75t_R FILLER_131_574 ();
 DECAPx4_ASAP7_75t_R FILLER_131_590 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_600 ();
 DECAPx10_ASAP7_75t_R FILLER_131_618 ();
 DECAPx6_ASAP7_75t_R FILLER_131_640 ();
 DECAPx2_ASAP7_75t_R FILLER_131_654 ();
 DECAPx1_ASAP7_75t_R FILLER_131_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_672 ();
 DECAPx4_ASAP7_75t_R FILLER_131_679 ();
 FILLER_ASAP7_75t_R FILLER_131_696 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_701 ();
 DECAPx1_ASAP7_75t_R FILLER_131_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_716 ();
 DECAPx6_ASAP7_75t_R FILLER_131_725 ();
 DECAPx2_ASAP7_75t_R FILLER_131_739 ();
 FILLER_ASAP7_75t_R FILLER_131_752 ();
 DECAPx4_ASAP7_75t_R FILLER_131_760 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_770 ();
 DECAPx10_ASAP7_75t_R FILLER_131_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_801 ();
 DECAPx6_ASAP7_75t_R FILLER_131_811 ();
 DECAPx1_ASAP7_75t_R FILLER_131_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_829 ();
 DECAPx1_ASAP7_75t_R FILLER_131_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_843 ();
 DECAPx4_ASAP7_75t_R FILLER_131_858 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_868 ();
 DECAPx4_ASAP7_75t_R FILLER_131_878 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_888 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_897 ();
 DECAPx4_ASAP7_75t_R FILLER_131_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_924 ();
 FILLER_ASAP7_75t_R FILLER_131_927 ();
 FILLER_ASAP7_75t_R FILLER_131_936 ();
 FILLER_ASAP7_75t_R FILLER_131_944 ();
 FILLER_ASAP7_75t_R FILLER_131_952 ();
 FILLER_ASAP7_75t_R FILLER_131_960 ();
 DECAPx1_ASAP7_75t_R FILLER_131_968 ();
 DECAPx2_ASAP7_75t_R FILLER_131_975 ();
 FILLER_ASAP7_75t_R FILLER_131_981 ();
 DECAPx4_ASAP7_75t_R FILLER_131_987 ();
 FILLER_ASAP7_75t_R FILLER_131_997 ();
 FILLER_ASAP7_75t_R FILLER_131_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1010 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_1016 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1057 ();
 DECAPx4_ASAP7_75t_R FILLER_131_1067 ();
 FILLER_ASAP7_75t_R FILLER_131_1077 ();
 DECAPx4_ASAP7_75t_R FILLER_131_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1095 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_1102 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1128 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1132 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_1146 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1155 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_131_1181 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_131_1220 ();
 FILLER_ASAP7_75t_R FILLER_131_1226 ();
 DECAPx4_ASAP7_75t_R FILLER_131_1238 ();
 FILLER_ASAP7_75t_R FILLER_131_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_131_1259 ();
 DECAPx6_ASAP7_75t_R FILLER_131_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_131_1305 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_1327 ();
 FILLER_ASAP7_75t_R FILLER_131_1331 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1336 ();
 DECAPx1_ASAP7_75t_R FILLER_131_1349 ();
 FILLER_ASAP7_75t_R FILLER_131_1359 ();
 FILLER_ASAP7_75t_R FILLER_131_1367 ();
 FILLER_ASAP7_75t_R FILLER_131_1375 ();
 DECAPx4_ASAP7_75t_R FILLER_132_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_12 ();
 DECAPx4_ASAP7_75t_R FILLER_132_41 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_51 ();
 DECAPx1_ASAP7_75t_R FILLER_132_62 ();
 FILLER_ASAP7_75t_R FILLER_132_74 ();
 DECAPx2_ASAP7_75t_R FILLER_132_84 ();
 FILLER_ASAP7_75t_R FILLER_132_96 ();
 FILLER_ASAP7_75t_R FILLER_132_105 ();
 FILLER_ASAP7_75t_R FILLER_132_114 ();
 DECAPx1_ASAP7_75t_R FILLER_132_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_123 ();
 DECAPx6_ASAP7_75t_R FILLER_132_131 ();
 FILLER_ASAP7_75t_R FILLER_132_145 ();
 DECAPx10_ASAP7_75t_R FILLER_132_167 ();
 DECAPx10_ASAP7_75t_R FILLER_132_189 ();
 DECAPx2_ASAP7_75t_R FILLER_132_211 ();
 FILLER_ASAP7_75t_R FILLER_132_217 ();
 DECAPx2_ASAP7_75t_R FILLER_132_225 ();
 FILLER_ASAP7_75t_R FILLER_132_257 ();
 DECAPx10_ASAP7_75t_R FILLER_132_262 ();
 DECAPx1_ASAP7_75t_R FILLER_132_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_288 ();
 DECAPx6_ASAP7_75t_R FILLER_132_315 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_329 ();
 FILLER_ASAP7_75t_R FILLER_132_340 ();
 DECAPx2_ASAP7_75t_R FILLER_132_348 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_354 ();
 DECAPx1_ASAP7_75t_R FILLER_132_363 ();
 FILLER_ASAP7_75t_R FILLER_132_370 ();
 DECAPx10_ASAP7_75t_R FILLER_132_398 ();
 DECAPx10_ASAP7_75t_R FILLER_132_420 ();
 DECAPx6_ASAP7_75t_R FILLER_132_442 ();
 DECAPx2_ASAP7_75t_R FILLER_132_456 ();
 FILLER_ASAP7_75t_R FILLER_132_464 ();
 DECAPx10_ASAP7_75t_R FILLER_132_474 ();
 DECAPx4_ASAP7_75t_R FILLER_132_496 ();
 FILLER_ASAP7_75t_R FILLER_132_506 ();
 DECAPx2_ASAP7_75t_R FILLER_132_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_520 ();
 FILLER_ASAP7_75t_R FILLER_132_533 ();
 FILLER_ASAP7_75t_R FILLER_132_561 ();
 DECAPx2_ASAP7_75t_R FILLER_132_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_572 ();
 FILLER_ASAP7_75t_R FILLER_132_583 ();
 DECAPx1_ASAP7_75t_R FILLER_132_591 ();
 DECAPx2_ASAP7_75t_R FILLER_132_603 ();
 FILLER_ASAP7_75t_R FILLER_132_609 ();
 DECAPx4_ASAP7_75t_R FILLER_132_617 ();
 FILLER_ASAP7_75t_R FILLER_132_627 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_635 ();
 DECAPx1_ASAP7_75t_R FILLER_132_646 ();
 DECAPx4_ASAP7_75t_R FILLER_132_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_670 ();
 FILLER_ASAP7_75t_R FILLER_132_683 ();
 DECAPx2_ASAP7_75t_R FILLER_132_697 ();
 FILLER_ASAP7_75t_R FILLER_132_711 ();
 DECAPx2_ASAP7_75t_R FILLER_132_723 ();
 DECAPx6_ASAP7_75t_R FILLER_132_737 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_751 ();
 FILLER_ASAP7_75t_R FILLER_132_761 ();
 DECAPx6_ASAP7_75t_R FILLER_132_769 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_783 ();
 DECAPx4_ASAP7_75t_R FILLER_132_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_806 ();
 DECAPx6_ASAP7_75t_R FILLER_132_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_832 ();
 DECAPx4_ASAP7_75t_R FILLER_132_839 ();
 DECAPx4_ASAP7_75t_R FILLER_132_855 ();
 FILLER_ASAP7_75t_R FILLER_132_877 ();
 DECAPx10_ASAP7_75t_R FILLER_132_887 ();
 DECAPx2_ASAP7_75t_R FILLER_132_909 ();
 FILLER_ASAP7_75t_R FILLER_132_915 ();
 FILLER_ASAP7_75t_R FILLER_132_925 ();
 DECAPx4_ASAP7_75t_R FILLER_132_937 ();
 FILLER_ASAP7_75t_R FILLER_132_947 ();
 FILLER_ASAP7_75t_R FILLER_132_955 ();
 FILLER_ASAP7_75t_R FILLER_132_983 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_993 ();
 FILLER_ASAP7_75t_R FILLER_132_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1015 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_1031 ();
 DECAPx6_ASAP7_75t_R FILLER_132_1040 ();
 DECAPx1_ASAP7_75t_R FILLER_132_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1058 ();
 DECAPx6_ASAP7_75t_R FILLER_132_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1076 ();
 DECAPx6_ASAP7_75t_R FILLER_132_1087 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_1101 ();
 FILLER_ASAP7_75t_R FILLER_132_1113 ();
 FILLER_ASAP7_75t_R FILLER_132_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_132_1131 ();
 DECAPx1_ASAP7_75t_R FILLER_132_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_132_1158 ();
 FILLER_ASAP7_75t_R FILLER_132_1180 ();
 DECAPx4_ASAP7_75t_R FILLER_132_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1202 ();
 DECAPx6_ASAP7_75t_R FILLER_132_1223 ();
 DECAPx1_ASAP7_75t_R FILLER_132_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1241 ();
 DECAPx6_ASAP7_75t_R FILLER_132_1245 ();
 DECAPx2_ASAP7_75t_R FILLER_132_1259 ();
 DECAPx1_ASAP7_75t_R FILLER_132_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1295 ();
 DECAPx4_ASAP7_75t_R FILLER_132_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1332 ();
 DECAPx1_ASAP7_75t_R FILLER_132_1353 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_1357 ();
 DECAPx1_ASAP7_75t_R FILLER_132_1366 ();
 FILLER_ASAP7_75t_R FILLER_132_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_133_2 ();
 FILLER_ASAP7_75t_R FILLER_133_16 ();
 DECAPx6_ASAP7_75t_R FILLER_133_24 ();
 DECAPx2_ASAP7_75t_R FILLER_133_38 ();
 DECAPx2_ASAP7_75t_R FILLER_133_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_53 ();
 DECAPx10_ASAP7_75t_R FILLER_133_57 ();
 DECAPx4_ASAP7_75t_R FILLER_133_79 ();
 FILLER_ASAP7_75t_R FILLER_133_115 ();
 DECAPx1_ASAP7_75t_R FILLER_133_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_127 ();
 DECAPx4_ASAP7_75t_R FILLER_133_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_147 ();
 DECAPx6_ASAP7_75t_R FILLER_133_156 ();
 DECAPx1_ASAP7_75t_R FILLER_133_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_174 ();
 DECAPx6_ASAP7_75t_R FILLER_133_183 ();
 FILLER_ASAP7_75t_R FILLER_133_203 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_133_208 ();
 FILLER_ASAP7_75t_R FILLER_133_237 ();
 DECAPx2_ASAP7_75t_R FILLER_133_245 ();
 FILLER_ASAP7_75t_R FILLER_133_257 ();
 DECAPx1_ASAP7_75t_R FILLER_133_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_269 ();
 FILLER_ASAP7_75t_R FILLER_133_278 ();
 DECAPx2_ASAP7_75t_R FILLER_133_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_293 ();
 FILLER_ASAP7_75t_R FILLER_133_297 ();
 DECAPx2_ASAP7_75t_R FILLER_133_305 ();
 DECAPx6_ASAP7_75t_R FILLER_133_317 ();
 DECAPx1_ASAP7_75t_R FILLER_133_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_335 ();
 DECAPx4_ASAP7_75t_R FILLER_133_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_352 ();
 DECAPx1_ASAP7_75t_R FILLER_133_379 ();
 FILLER_ASAP7_75t_R FILLER_133_389 ();
 DECAPx10_ASAP7_75t_R FILLER_133_394 ();
 DECAPx6_ASAP7_75t_R FILLER_133_416 ();
 FILLER_ASAP7_75t_R FILLER_133_430 ();
 FILLER_ASAP7_75t_R FILLER_133_439 ();
 FILLER_ASAP7_75t_R FILLER_133_447 ();
 DECAPx4_ASAP7_75t_R FILLER_133_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_462 ();
 DECAPx4_ASAP7_75t_R FILLER_133_466 ();
 FILLER_ASAP7_75t_R FILLER_133_476 ();
 DECAPx10_ASAP7_75t_R FILLER_133_485 ();
 DECAPx1_ASAP7_75t_R FILLER_133_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_511 ();
 DECAPx1_ASAP7_75t_R FILLER_133_522 ();
 FILLER_ASAP7_75t_R FILLER_133_532 ();
 DECAPx6_ASAP7_75t_R FILLER_133_541 ();
 DECAPx1_ASAP7_75t_R FILLER_133_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_559 ();
 DECAPx4_ASAP7_75t_R FILLER_133_568 ();
 DECAPx10_ASAP7_75t_R FILLER_133_588 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_133_610 ();
 DECAPx2_ASAP7_75t_R FILLER_133_619 ();
 FILLER_ASAP7_75t_R FILLER_133_631 ();
 DECAPx4_ASAP7_75t_R FILLER_133_639 ();
 FILLER_ASAP7_75t_R FILLER_133_649 ();
 DECAPx10_ASAP7_75t_R FILLER_133_661 ();
 DECAPx4_ASAP7_75t_R FILLER_133_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_693 ();
 DECAPx2_ASAP7_75t_R FILLER_133_700 ();
 FILLER_ASAP7_75t_R FILLER_133_706 ();
 DECAPx2_ASAP7_75t_R FILLER_133_714 ();
 FILLER_ASAP7_75t_R FILLER_133_720 ();
 DECAPx2_ASAP7_75t_R FILLER_133_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_736 ();
 FILLER_ASAP7_75t_R FILLER_133_743 ();
 DECAPx1_ASAP7_75t_R FILLER_133_751 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_133_761 ();
 FILLER_ASAP7_75t_R FILLER_133_770 ();
 DECAPx4_ASAP7_75t_R FILLER_133_782 ();
 FILLER_ASAP7_75t_R FILLER_133_792 ();
 DECAPx1_ASAP7_75t_R FILLER_133_800 ();
 FILLER_ASAP7_75t_R FILLER_133_818 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_133_830 ();
 DECAPx10_ASAP7_75t_R FILLER_133_841 ();
 DECAPx2_ASAP7_75t_R FILLER_133_863 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_133_869 ();
 DECAPx4_ASAP7_75t_R FILLER_133_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_886 ();
 DECAPx10_ASAP7_75t_R FILLER_133_893 ();
 DECAPx4_ASAP7_75t_R FILLER_133_915 ();
 DECAPx4_ASAP7_75t_R FILLER_133_927 ();
 DECAPx10_ASAP7_75t_R FILLER_133_943 ();
 DECAPx10_ASAP7_75t_R FILLER_133_965 ();
 DECAPx4_ASAP7_75t_R FILLER_133_987 ();
 FILLER_ASAP7_75t_R FILLER_133_997 ();
 FILLER_ASAP7_75t_R FILLER_133_1008 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1016 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_133_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1035 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1049 ();
 DECAPx4_ASAP7_75t_R FILLER_133_1061 ();
 FILLER_ASAP7_75t_R FILLER_133_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1103 ();
 FILLER_ASAP7_75t_R FILLER_133_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1135 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_133_1141 ();
 FILLER_ASAP7_75t_R FILLER_133_1170 ();
 FILLER_ASAP7_75t_R FILLER_133_1178 ();
 FILLER_ASAP7_75t_R FILLER_133_1206 ();
 FILLER_ASAP7_75t_R FILLER_133_1211 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1223 ();
 FILLER_ASAP7_75t_R FILLER_133_1253 ();
 DECAPx2_ASAP7_75t_R FILLER_133_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1267 ();
 FILLER_ASAP7_75t_R FILLER_133_1278 ();
 DECAPx1_ASAP7_75t_R FILLER_133_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_1292 ();
 FILLER_ASAP7_75t_R FILLER_133_1301 ();
 FILLER_ASAP7_75t_R FILLER_133_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_133_1314 ();
 DECAPx4_ASAP7_75t_R FILLER_133_1336 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_133_1346 ();
 FILLER_ASAP7_75t_R FILLER_133_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_134_2 ();
 DECAPx2_ASAP7_75t_R FILLER_134_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_22 ();
 DECAPx1_ASAP7_75t_R FILLER_134_29 ();
 DECAPx2_ASAP7_75t_R FILLER_134_39 ();
 FILLER_ASAP7_75t_R FILLER_134_45 ();
 FILLER_ASAP7_75t_R FILLER_134_73 ();
 DECAPx2_ASAP7_75t_R FILLER_134_81 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_87 ();
 FILLER_ASAP7_75t_R FILLER_134_100 ();
 FILLER_ASAP7_75t_R FILLER_134_105 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_114 ();
 FILLER_ASAP7_75t_R FILLER_134_123 ();
 DECAPx4_ASAP7_75t_R FILLER_134_131 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_141 ();
 DECAPx2_ASAP7_75t_R FILLER_134_153 ();
 FILLER_ASAP7_75t_R FILLER_134_165 ();
 FILLER_ASAP7_75t_R FILLER_134_173 ();
 DECAPx2_ASAP7_75t_R FILLER_134_181 ();
 FILLER_ASAP7_75t_R FILLER_134_213 ();
 DECAPx1_ASAP7_75t_R FILLER_134_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_225 ();
 DECAPx4_ASAP7_75t_R FILLER_134_229 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_239 ();
 FILLER_ASAP7_75t_R FILLER_134_245 ();
 FILLER_ASAP7_75t_R FILLER_134_273 ();
 DECAPx10_ASAP7_75t_R FILLER_134_281 ();
 FILLER_ASAP7_75t_R FILLER_134_303 ();
 FILLER_ASAP7_75t_R FILLER_134_311 ();
 DECAPx2_ASAP7_75t_R FILLER_134_321 ();
 FILLER_ASAP7_75t_R FILLER_134_327 ();
 DECAPx6_ASAP7_75t_R FILLER_134_335 ();
 FILLER_ASAP7_75t_R FILLER_134_355 ();
 DECAPx10_ASAP7_75t_R FILLER_134_363 ();
 DECAPx2_ASAP7_75t_R FILLER_134_385 ();
 FILLER_ASAP7_75t_R FILLER_134_394 ();
 FILLER_ASAP7_75t_R FILLER_134_404 ();
 FILLER_ASAP7_75t_R FILLER_134_413 ();
 DECAPx1_ASAP7_75t_R FILLER_134_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_425 ();
 FILLER_ASAP7_75t_R FILLER_134_452 ();
 DECAPx1_ASAP7_75t_R FILLER_134_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_461 ();
 FILLER_ASAP7_75t_R FILLER_134_464 ();
 DECAPx2_ASAP7_75t_R FILLER_134_472 ();
 FILLER_ASAP7_75t_R FILLER_134_478 ();
 DECAPx6_ASAP7_75t_R FILLER_134_486 ();
 FILLER_ASAP7_75t_R FILLER_134_500 ();
 DECAPx1_ASAP7_75t_R FILLER_134_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_512 ();
 DECAPx1_ASAP7_75t_R FILLER_134_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_527 ();
 DECAPx4_ASAP7_75t_R FILLER_134_534 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_544 ();
 DECAPx1_ASAP7_75t_R FILLER_134_550 ();
 FILLER_ASAP7_75t_R FILLER_134_560 ();
 DECAPx2_ASAP7_75t_R FILLER_134_570 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_576 ();
 DECAPx10_ASAP7_75t_R FILLER_134_585 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_607 ();
 DECAPx2_ASAP7_75t_R FILLER_134_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_622 ();
 FILLER_ASAP7_75t_R FILLER_134_629 ();
 DECAPx1_ASAP7_75t_R FILLER_134_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_643 ();
 DECAPx4_ASAP7_75t_R FILLER_134_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_661 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_669 ();
 FILLER_ASAP7_75t_R FILLER_134_679 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_687 ();
 DECAPx4_ASAP7_75t_R FILLER_134_702 ();
 FILLER_ASAP7_75t_R FILLER_134_712 ();
 DECAPx10_ASAP7_75t_R FILLER_134_720 ();
 DECAPx4_ASAP7_75t_R FILLER_134_742 ();
 FILLER_ASAP7_75t_R FILLER_134_752 ();
 DECAPx6_ASAP7_75t_R FILLER_134_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_775 ();
 DECAPx2_ASAP7_75t_R FILLER_134_787 ();
 FILLER_ASAP7_75t_R FILLER_134_793 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_802 ();
 FILLER_ASAP7_75t_R FILLER_134_808 ();
 DECAPx6_ASAP7_75t_R FILLER_134_813 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_827 ();
 FILLER_ASAP7_75t_R FILLER_134_839 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_844 ();
 DECAPx6_ASAP7_75t_R FILLER_134_859 ();
 DECAPx1_ASAP7_75t_R FILLER_134_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_877 ();
 DECAPx1_ASAP7_75t_R FILLER_134_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_885 ();
 FILLER_ASAP7_75t_R FILLER_134_892 ();
 DECAPx2_ASAP7_75t_R FILLER_134_904 ();
 FILLER_ASAP7_75t_R FILLER_134_916 ();
 DECAPx4_ASAP7_75t_R FILLER_134_921 ();
 FILLER_ASAP7_75t_R FILLER_134_931 ();
 FILLER_ASAP7_75t_R FILLER_134_940 ();
 DECAPx2_ASAP7_75t_R FILLER_134_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_955 ();
 DECAPx4_ASAP7_75t_R FILLER_134_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_974 ();
 DECAPx6_ASAP7_75t_R FILLER_134_981 ();
 FILLER_ASAP7_75t_R FILLER_134_995 ();
 DECAPx6_ASAP7_75t_R FILLER_134_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1014 ();
 FILLER_ASAP7_75t_R FILLER_134_1023 ();
 DECAPx6_ASAP7_75t_R FILLER_134_1028 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1048 ();
 FILLER_ASAP7_75t_R FILLER_134_1055 ();
 DECAPx6_ASAP7_75t_R FILLER_134_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1079 ();
 FILLER_ASAP7_75t_R FILLER_134_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1093 ();
 FILLER_ASAP7_75t_R FILLER_134_1103 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_134_1127 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1139 ();
 FILLER_ASAP7_75t_R FILLER_134_1149 ();
 FILLER_ASAP7_75t_R FILLER_134_1159 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1164 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_1174 ();
 FILLER_ASAP7_75t_R FILLER_134_1183 ();
 FILLER_ASAP7_75t_R FILLER_134_1193 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1198 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_1208 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1217 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_1223 ();
 FILLER_ASAP7_75t_R FILLER_134_1234 ();
 FILLER_ASAP7_75t_R FILLER_134_1244 ();
 FILLER_ASAP7_75t_R FILLER_134_1249 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1260 ();
 FILLER_ASAP7_75t_R FILLER_134_1272 ();
 FILLER_ASAP7_75t_R FILLER_134_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_134_1307 ();
 FILLER_ASAP7_75t_R FILLER_134_1335 ();
 DECAPx4_ASAP7_75t_R FILLER_134_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_1353 ();
 FILLER_ASAP7_75t_R FILLER_134_1364 ();
 DECAPx2_ASAP7_75t_R FILLER_134_1369 ();
 FILLER_ASAP7_75t_R FILLER_134_1375 ();
 FILLER_ASAP7_75t_R FILLER_135_2 ();
 DECAPx2_ASAP7_75t_R FILLER_135_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_16 ();
 DECAPx2_ASAP7_75t_R FILLER_135_43 ();
 FILLER_ASAP7_75t_R FILLER_135_49 ();
 DECAPx4_ASAP7_75t_R FILLER_135_57 ();
 FILLER_ASAP7_75t_R FILLER_135_67 ();
 DECAPx6_ASAP7_75t_R FILLER_135_95 ();
 FILLER_ASAP7_75t_R FILLER_135_109 ();
 DECAPx6_ASAP7_75t_R FILLER_135_117 ();
 FILLER_ASAP7_75t_R FILLER_135_138 ();
 DECAPx6_ASAP7_75t_R FILLER_135_148 ();
 DECAPx2_ASAP7_75t_R FILLER_135_168 ();
 FILLER_ASAP7_75t_R FILLER_135_174 ();
 DECAPx6_ASAP7_75t_R FILLER_135_179 ();
 FILLER_ASAP7_75t_R FILLER_135_199 ();
 DECAPx6_ASAP7_75t_R FILLER_135_204 ();
 DECAPx2_ASAP7_75t_R FILLER_135_218 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_230 ();
 DECAPx10_ASAP7_75t_R FILLER_135_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_261 ();
 DECAPx1_ASAP7_75t_R FILLER_135_265 ();
 DECAPx6_ASAP7_75t_R FILLER_135_275 ();
 DECAPx1_ASAP7_75t_R FILLER_135_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_293 ();
 DECAPx4_ASAP7_75t_R FILLER_135_300 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_310 ();
 DECAPx1_ASAP7_75t_R FILLER_135_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_325 ();
 FILLER_ASAP7_75t_R FILLER_135_337 ();
 DECAPx2_ASAP7_75t_R FILLER_135_346 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_352 ();
 DECAPx4_ASAP7_75t_R FILLER_135_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_371 ();
 DECAPx6_ASAP7_75t_R FILLER_135_378 ();
 DECAPx2_ASAP7_75t_R FILLER_135_392 ();
 FILLER_ASAP7_75t_R FILLER_135_420 ();
 DECAPx6_ASAP7_75t_R FILLER_135_428 ();
 DECAPx2_ASAP7_75t_R FILLER_135_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_470 ();
 DECAPx2_ASAP7_75t_R FILLER_135_480 ();
 FILLER_ASAP7_75t_R FILLER_135_492 ();
 FILLER_ASAP7_75t_R FILLER_135_503 ();
 DECAPx2_ASAP7_75t_R FILLER_135_512 ();
 FILLER_ASAP7_75t_R FILLER_135_518 ();
 DECAPx1_ASAP7_75t_R FILLER_135_532 ();
 FILLER_ASAP7_75t_R FILLER_135_542 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_550 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_561 ();
 DECAPx6_ASAP7_75t_R FILLER_135_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_584 ();
 FILLER_ASAP7_75t_R FILLER_135_589 ();
 DECAPx4_ASAP7_75t_R FILLER_135_601 ();
 DECAPx6_ASAP7_75t_R FILLER_135_619 ();
 FILLER_ASAP7_75t_R FILLER_135_633 ();
 FILLER_ASAP7_75t_R FILLER_135_641 ();
 DECAPx10_ASAP7_75t_R FILLER_135_650 ();
 DECAPx1_ASAP7_75t_R FILLER_135_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_688 ();
 DECAPx10_ASAP7_75t_R FILLER_135_697 ();
 FILLER_ASAP7_75t_R FILLER_135_719 ();
 DECAPx4_ASAP7_75t_R FILLER_135_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_739 ();
 FILLER_ASAP7_75t_R FILLER_135_747 ();
 FILLER_ASAP7_75t_R FILLER_135_755 ();
 DECAPx4_ASAP7_75t_R FILLER_135_765 ();
 DECAPx6_ASAP7_75t_R FILLER_135_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_805 ();
 DECAPx4_ASAP7_75t_R FILLER_135_815 ();
 FILLER_ASAP7_75t_R FILLER_135_825 ();
 FILLER_ASAP7_75t_R FILLER_135_836 ();
 DECAPx2_ASAP7_75t_R FILLER_135_844 ();
 FILLER_ASAP7_75t_R FILLER_135_850 ();
 DECAPx4_ASAP7_75t_R FILLER_135_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_870 ();
 DECAPx4_ASAP7_75t_R FILLER_135_879 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_889 ();
 DECAPx2_ASAP7_75t_R FILLER_135_898 ();
 FILLER_ASAP7_75t_R FILLER_135_913 ();
 FILLER_ASAP7_75t_R FILLER_135_923 ();
 FILLER_ASAP7_75t_R FILLER_135_927 ();
 DECAPx6_ASAP7_75t_R FILLER_135_935 ();
 DECAPx2_ASAP7_75t_R FILLER_135_963 ();
 FILLER_ASAP7_75t_R FILLER_135_969 ();
 FILLER_ASAP7_75t_R FILLER_135_980 ();
 DECAPx2_ASAP7_75t_R FILLER_135_990 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_996 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_135_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1053 ();
 DECAPx6_ASAP7_75t_R FILLER_135_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1107 ();
 DECAPx6_ASAP7_75t_R FILLER_135_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_135_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1200 ();
 DECAPx2_ASAP7_75t_R FILLER_135_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1228 ();
 FILLER_ASAP7_75t_R FILLER_135_1235 ();
 DECAPx2_ASAP7_75t_R FILLER_135_1243 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_135_1255 ();
 DECAPx6_ASAP7_75t_R FILLER_135_1285 ();
 DECAPx1_ASAP7_75t_R FILLER_135_1299 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1303 ();
 FILLER_ASAP7_75t_R FILLER_135_1310 ();
 DECAPx4_ASAP7_75t_R FILLER_135_1318 ();
 FILLER_ASAP7_75t_R FILLER_135_1328 ();
 DECAPx6_ASAP7_75t_R FILLER_135_1336 ();
 DECAPx2_ASAP7_75t_R FILLER_135_1350 ();
 DECAPx6_ASAP7_75t_R FILLER_135_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_1376 ();
 FILLER_ASAP7_75t_R FILLER_136_2 ();
 DECAPx6_ASAP7_75t_R FILLER_136_10 ();
 DECAPx2_ASAP7_75t_R FILLER_136_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_30 ();
 DECAPx6_ASAP7_75t_R FILLER_136_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_48 ();
 DECAPx2_ASAP7_75t_R FILLER_136_55 ();
 DECAPx2_ASAP7_75t_R FILLER_136_64 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_70 ();
 DECAPx1_ASAP7_75t_R FILLER_136_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_83 ();
 DECAPx10_ASAP7_75t_R FILLER_136_87 ();
 DECAPx4_ASAP7_75t_R FILLER_136_109 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_119 ();
 DECAPx4_ASAP7_75t_R FILLER_136_128 ();
 FILLER_ASAP7_75t_R FILLER_136_146 ();
 DECAPx1_ASAP7_75t_R FILLER_136_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_158 ();
 DECAPx10_ASAP7_75t_R FILLER_136_185 ();
 DECAPx2_ASAP7_75t_R FILLER_136_207 ();
 FILLER_ASAP7_75t_R FILLER_136_213 ();
 DECAPx1_ASAP7_75t_R FILLER_136_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_225 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_232 ();
 DECAPx10_ASAP7_75t_R FILLER_136_243 ();
 DECAPx6_ASAP7_75t_R FILLER_136_265 ();
 DECAPx1_ASAP7_75t_R FILLER_136_279 ();
 FILLER_ASAP7_75t_R FILLER_136_309 ();
 DECAPx10_ASAP7_75t_R FILLER_136_314 ();
 DECAPx6_ASAP7_75t_R FILLER_136_336 ();
 FILLER_ASAP7_75t_R FILLER_136_350 ();
 FILLER_ASAP7_75t_R FILLER_136_362 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_370 ();
 FILLER_ASAP7_75t_R FILLER_136_381 ();
 DECAPx2_ASAP7_75t_R FILLER_136_386 ();
 FILLER_ASAP7_75t_R FILLER_136_392 ();
 FILLER_ASAP7_75t_R FILLER_136_402 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_410 ();
 FILLER_ASAP7_75t_R FILLER_136_439 ();
 DECAPx1_ASAP7_75t_R FILLER_136_447 ();
 DECAPx2_ASAP7_75t_R FILLER_136_454 ();
 FILLER_ASAP7_75t_R FILLER_136_460 ();
 FILLER_ASAP7_75t_R FILLER_136_464 ();
 DECAPx10_ASAP7_75t_R FILLER_136_472 ();
 DECAPx1_ASAP7_75t_R FILLER_136_494 ();
 DECAPx10_ASAP7_75t_R FILLER_136_504 ();
 DECAPx1_ASAP7_75t_R FILLER_136_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_530 ();
 DECAPx2_ASAP7_75t_R FILLER_136_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_547 ();
 DECAPx4_ASAP7_75t_R FILLER_136_554 ();
 FILLER_ASAP7_75t_R FILLER_136_572 ();
 DECAPx1_ASAP7_75t_R FILLER_136_580 ();
 FILLER_ASAP7_75t_R FILLER_136_590 ();
 DECAPx2_ASAP7_75t_R FILLER_136_600 ();
 FILLER_ASAP7_75t_R FILLER_136_606 ();
 DECAPx10_ASAP7_75t_R FILLER_136_616 ();
 DECAPx2_ASAP7_75t_R FILLER_136_638 ();
 FILLER_ASAP7_75t_R FILLER_136_644 ();
 DECAPx1_ASAP7_75t_R FILLER_136_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_666 ();
 DECAPx6_ASAP7_75t_R FILLER_136_673 ();
 DECAPx2_ASAP7_75t_R FILLER_136_687 ();
 DECAPx2_ASAP7_75t_R FILLER_136_701 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_707 ();
 DECAPx2_ASAP7_75t_R FILLER_136_716 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_722 ();
 DECAPx2_ASAP7_75t_R FILLER_136_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_739 ();
 DECAPx2_ASAP7_75t_R FILLER_136_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_753 ();
 FILLER_ASAP7_75t_R FILLER_136_765 ();
 DECAPx6_ASAP7_75t_R FILLER_136_775 ();
 DECAPx1_ASAP7_75t_R FILLER_136_789 ();
 DECAPx1_ASAP7_75t_R FILLER_136_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_803 ();
 DECAPx1_ASAP7_75t_R FILLER_136_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_815 ();
 DECAPx6_ASAP7_75t_R FILLER_136_823 ();
 DECAPx1_ASAP7_75t_R FILLER_136_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_841 ();
 FILLER_ASAP7_75t_R FILLER_136_848 ();
 FILLER_ASAP7_75t_R FILLER_136_860 ();
 DECAPx10_ASAP7_75t_R FILLER_136_876 ();
 DECAPx2_ASAP7_75t_R FILLER_136_898 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_904 ();
 DECAPx2_ASAP7_75t_R FILLER_136_910 ();
 DECAPx1_ASAP7_75t_R FILLER_136_925 ();
 DECAPx2_ASAP7_75t_R FILLER_136_935 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_941 ();
 DECAPx2_ASAP7_75t_R FILLER_136_951 ();
 DECAPx1_ASAP7_75t_R FILLER_136_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_968 ();
 DECAPx1_ASAP7_75t_R FILLER_136_972 ();
 DECAPx4_ASAP7_75t_R FILLER_136_979 ();
 FILLER_ASAP7_75t_R FILLER_136_989 ();
 DECAPx1_ASAP7_75t_R FILLER_136_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_998 ();
 FILLER_ASAP7_75t_R FILLER_136_1005 ();
 FILLER_ASAP7_75t_R FILLER_136_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1021 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_1027 ();
 FILLER_ASAP7_75t_R FILLER_136_1037 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1065 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_1075 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1087 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_1103 ();
 FILLER_ASAP7_75t_R FILLER_136_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1120 ();
 FILLER_ASAP7_75t_R FILLER_136_1126 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1146 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1153 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_1166 ();
 DECAPx4_ASAP7_75t_R FILLER_136_1177 ();
 FILLER_ASAP7_75t_R FILLER_136_1213 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1223 ();
 DECAPx6_ASAP7_75t_R FILLER_136_1232 ();
 FILLER_ASAP7_75t_R FILLER_136_1246 ();
 DECAPx6_ASAP7_75t_R FILLER_136_1256 ();
 DECAPx1_ASAP7_75t_R FILLER_136_1296 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_1300 ();
 FILLER_ASAP7_75t_R FILLER_136_1309 ();
 FILLER_ASAP7_75t_R FILLER_136_1337 ();
 DECAPx2_ASAP7_75t_R FILLER_136_1349 ();
 FILLER_ASAP7_75t_R FILLER_136_1355 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_1367 ();
 FILLER_ASAP7_75t_R FILLER_136_1375 ();
 FILLER_ASAP7_75t_R FILLER_137_2 ();
 DECAPx2_ASAP7_75t_R FILLER_137_10 ();
 FILLER_ASAP7_75t_R FILLER_137_16 ();
 DECAPx6_ASAP7_75t_R FILLER_137_24 ();
 DECAPx1_ASAP7_75t_R FILLER_137_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_42 ();
 DECAPx10_ASAP7_75t_R FILLER_137_49 ();
 DECAPx1_ASAP7_75t_R FILLER_137_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_75 ();
 FILLER_ASAP7_75t_R FILLER_137_102 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_110 ();
 FILLER_ASAP7_75t_R FILLER_137_119 ();
 FILLER_ASAP7_75t_R FILLER_137_129 ();
 DECAPx10_ASAP7_75t_R FILLER_137_137 ();
 FILLER_ASAP7_75t_R FILLER_137_159 ();
 DECAPx2_ASAP7_75t_R FILLER_137_167 ();
 DECAPx2_ASAP7_75t_R FILLER_137_176 ();
 FILLER_ASAP7_75t_R FILLER_137_188 ();
 DECAPx2_ASAP7_75t_R FILLER_137_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_202 ();
 DECAPx1_ASAP7_75t_R FILLER_137_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_233 ();
 DECAPx6_ASAP7_75t_R FILLER_137_244 ();
 DECAPx2_ASAP7_75t_R FILLER_137_264 ();
 FILLER_ASAP7_75t_R FILLER_137_270 ();
 DECAPx1_ASAP7_75t_R FILLER_137_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_279 ();
 FILLER_ASAP7_75t_R FILLER_137_288 ();
 FILLER_ASAP7_75t_R FILLER_137_296 ();
 DECAPx10_ASAP7_75t_R FILLER_137_301 ();
 DECAPx4_ASAP7_75t_R FILLER_137_323 ();
 FILLER_ASAP7_75t_R FILLER_137_333 ();
 DECAPx2_ASAP7_75t_R FILLER_137_346 ();
 DECAPx4_ASAP7_75t_R FILLER_137_358 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_368 ();
 FILLER_ASAP7_75t_R FILLER_137_377 ();
 DECAPx4_ASAP7_75t_R FILLER_137_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_395 ();
 FILLER_ASAP7_75t_R FILLER_137_402 ();
 DECAPx2_ASAP7_75t_R FILLER_137_410 ();
 DECAPx2_ASAP7_75t_R FILLER_137_422 ();
 FILLER_ASAP7_75t_R FILLER_137_431 ();
 FILLER_ASAP7_75t_R FILLER_137_440 ();
 DECAPx1_ASAP7_75t_R FILLER_137_445 ();
 FILLER_ASAP7_75t_R FILLER_137_455 ();
 FILLER_ASAP7_75t_R FILLER_137_465 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_474 ();
 FILLER_ASAP7_75t_R FILLER_137_483 ();
 DECAPx1_ASAP7_75t_R FILLER_137_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_501 ();
 DECAPx4_ASAP7_75t_R FILLER_137_508 ();
 FILLER_ASAP7_75t_R FILLER_137_518 ();
 DECAPx10_ASAP7_75t_R FILLER_137_526 ();
 DECAPx10_ASAP7_75t_R FILLER_137_548 ();
 DECAPx6_ASAP7_75t_R FILLER_137_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_584 ();
 DECAPx4_ASAP7_75t_R FILLER_137_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_605 ();
 DECAPx1_ASAP7_75t_R FILLER_137_612 ();
 DECAPx2_ASAP7_75t_R FILLER_137_623 ();
 FILLER_ASAP7_75t_R FILLER_137_635 ();
 DECAPx6_ASAP7_75t_R FILLER_137_644 ();
 FILLER_ASAP7_75t_R FILLER_137_658 ();
 FILLER_ASAP7_75t_R FILLER_137_666 ();
 DECAPx6_ASAP7_75t_R FILLER_137_679 ();
 FILLER_ASAP7_75t_R FILLER_137_693 ();
 DECAPx2_ASAP7_75t_R FILLER_137_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_709 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_716 ();
 FILLER_ASAP7_75t_R FILLER_137_725 ();
 FILLER_ASAP7_75t_R FILLER_137_733 ();
 DECAPx10_ASAP7_75t_R FILLER_137_741 ();
 DECAPx4_ASAP7_75t_R FILLER_137_763 ();
 FILLER_ASAP7_75t_R FILLER_137_773 ();
 DECAPx4_ASAP7_75t_R FILLER_137_781 ();
 FILLER_ASAP7_75t_R FILLER_137_799 ();
 FILLER_ASAP7_75t_R FILLER_137_810 ();
 FILLER_ASAP7_75t_R FILLER_137_819 ();
 FILLER_ASAP7_75t_R FILLER_137_828 ();
 DECAPx10_ASAP7_75t_R FILLER_137_835 ();
 DECAPx2_ASAP7_75t_R FILLER_137_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_863 ();
 DECAPx6_ASAP7_75t_R FILLER_137_875 ();
 DECAPx10_ASAP7_75t_R FILLER_137_897 ();
 DECAPx2_ASAP7_75t_R FILLER_137_919 ();
 DECAPx2_ASAP7_75t_R FILLER_137_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_933 ();
 DECAPx10_ASAP7_75t_R FILLER_137_944 ();
 DECAPx2_ASAP7_75t_R FILLER_137_966 ();
 FILLER_ASAP7_75t_R FILLER_137_972 ();
 FILLER_ASAP7_75t_R FILLER_137_983 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_991 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1019 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1026 ();
 FILLER_ASAP7_75t_R FILLER_137_1040 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1052 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_137_1065 ();
 FILLER_ASAP7_75t_R FILLER_137_1087 ();
 FILLER_ASAP7_75t_R FILLER_137_1092 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1103 ();
 FILLER_ASAP7_75t_R FILLER_137_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1122 ();
 FILLER_ASAP7_75t_R FILLER_137_1128 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1138 ();
 FILLER_ASAP7_75t_R FILLER_137_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1156 ();
 FILLER_ASAP7_75t_R FILLER_137_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1197 ();
 FILLER_ASAP7_75t_R FILLER_137_1215 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1227 ();
 FILLER_ASAP7_75t_R FILLER_137_1237 ();
 FILLER_ASAP7_75t_R FILLER_137_1242 ();
 DECAPx1_ASAP7_75t_R FILLER_137_1270 ();
 FILLER_ASAP7_75t_R FILLER_137_1284 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1289 ();
 FILLER_ASAP7_75t_R FILLER_137_1299 ();
 FILLER_ASAP7_75t_R FILLER_137_1304 ();
 FILLER_ASAP7_75t_R FILLER_137_1312 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1317 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_1323 ();
 DECAPx4_ASAP7_75t_R FILLER_137_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_1339 ();
 DECAPx2_ASAP7_75t_R FILLER_137_1343 ();
 FILLER_ASAP7_75t_R FILLER_137_1375 ();
 DECAPx1_ASAP7_75t_R FILLER_138_2 ();
 FILLER_ASAP7_75t_R FILLER_138_32 ();
 FILLER_ASAP7_75t_R FILLER_138_60 ();
 DECAPx2_ASAP7_75t_R FILLER_138_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_76 ();
 FILLER_ASAP7_75t_R FILLER_138_83 ();
 DECAPx1_ASAP7_75t_R FILLER_138_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_95 ();
 FILLER_ASAP7_75t_R FILLER_138_122 ();
 DECAPx4_ASAP7_75t_R FILLER_138_127 ();
 FILLER_ASAP7_75t_R FILLER_138_137 ();
 DECAPx6_ASAP7_75t_R FILLER_138_145 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_138_165 ();
 DECAPx4_ASAP7_75t_R FILLER_138_171 ();
 DECAPx1_ASAP7_75t_R FILLER_138_207 ();
 FILLER_ASAP7_75t_R FILLER_138_217 ();
 DECAPx2_ASAP7_75t_R FILLER_138_222 ();
 FILLER_ASAP7_75t_R FILLER_138_228 ();
 DECAPx2_ASAP7_75t_R FILLER_138_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_239 ();
 FILLER_ASAP7_75t_R FILLER_138_246 ();
 FILLER_ASAP7_75t_R FILLER_138_274 ();
 FILLER_ASAP7_75t_R FILLER_138_286 ();
 DECAPx4_ASAP7_75t_R FILLER_138_294 ();
 FILLER_ASAP7_75t_R FILLER_138_304 ();
 DECAPx4_ASAP7_75t_R FILLER_138_312 ();
 FILLER_ASAP7_75t_R FILLER_138_330 ();
 FILLER_ASAP7_75t_R FILLER_138_340 ();
 DECAPx2_ASAP7_75t_R FILLER_138_348 ();
 DECAPx4_ASAP7_75t_R FILLER_138_360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_138_370 ();
 DECAPx6_ASAP7_75t_R FILLER_138_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_393 ();
 FILLER_ASAP7_75t_R FILLER_138_400 ();
 DECAPx2_ASAP7_75t_R FILLER_138_420 ();
 FILLER_ASAP7_75t_R FILLER_138_426 ();
 DECAPx2_ASAP7_75t_R FILLER_138_454 ();
 FILLER_ASAP7_75t_R FILLER_138_460 ();
 FILLER_ASAP7_75t_R FILLER_138_464 ();
 DECAPx2_ASAP7_75t_R FILLER_138_473 ();
 DECAPx6_ASAP7_75t_R FILLER_138_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_501 ();
 FILLER_ASAP7_75t_R FILLER_138_509 ();
 FILLER_ASAP7_75t_R FILLER_138_518 ();
 FILLER_ASAP7_75t_R FILLER_138_528 ();
 DECAPx1_ASAP7_75t_R FILLER_138_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_540 ();
 FILLER_ASAP7_75t_R FILLER_138_547 ();
 DECAPx2_ASAP7_75t_R FILLER_138_556 ();
 FILLER_ASAP7_75t_R FILLER_138_562 ();
 FILLER_ASAP7_75t_R FILLER_138_571 ();
 DECAPx6_ASAP7_75t_R FILLER_138_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_593 ();
 DECAPx2_ASAP7_75t_R FILLER_138_600 ();
 FILLER_ASAP7_75t_R FILLER_138_606 ();
 DECAPx1_ASAP7_75t_R FILLER_138_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_620 ();
 DECAPx10_ASAP7_75t_R FILLER_138_627 ();
 DECAPx6_ASAP7_75t_R FILLER_138_649 ();
 DECAPx2_ASAP7_75t_R FILLER_138_663 ();
 DECAPx4_ASAP7_75t_R FILLER_138_675 ();
 DECAPx6_ASAP7_75t_R FILLER_138_693 ();
 FILLER_ASAP7_75t_R FILLER_138_707 ();
 DECAPx10_ASAP7_75t_R FILLER_138_716 ();
 DECAPx10_ASAP7_75t_R FILLER_138_738 ();
 DECAPx2_ASAP7_75t_R FILLER_138_760 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_138_766 ();
 DECAPx10_ASAP7_75t_R FILLER_138_776 ();
 DECAPx6_ASAP7_75t_R FILLER_138_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_812 ();
 DECAPx4_ASAP7_75t_R FILLER_138_819 ();
 FILLER_ASAP7_75t_R FILLER_138_829 ();
 DECAPx2_ASAP7_75t_R FILLER_138_836 ();
 FILLER_ASAP7_75t_R FILLER_138_842 ();
 DECAPx6_ASAP7_75t_R FILLER_138_852 ();
 DECAPx2_ASAP7_75t_R FILLER_138_875 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_138_881 ();
 FILLER_ASAP7_75t_R FILLER_138_890 ();
 FILLER_ASAP7_75t_R FILLER_138_895 ();
 DECAPx4_ASAP7_75t_R FILLER_138_900 ();
 FILLER_ASAP7_75t_R FILLER_138_910 ();
 DECAPx6_ASAP7_75t_R FILLER_138_918 ();
 DECAPx2_ASAP7_75t_R FILLER_138_938 ();
 FILLER_ASAP7_75t_R FILLER_138_944 ();
 FILLER_ASAP7_75t_R FILLER_138_954 ();
 DECAPx6_ASAP7_75t_R FILLER_138_964 ();
 FILLER_ASAP7_75t_R FILLER_138_978 ();
 DECAPx10_ASAP7_75t_R FILLER_138_990 ();
 DECAPx4_ASAP7_75t_R FILLER_138_1012 ();
 DECAPx4_ASAP7_75t_R FILLER_138_1048 ();
 FILLER_ASAP7_75t_R FILLER_138_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1096 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_138_1102 ();
 FILLER_ASAP7_75t_R FILLER_138_1131 ();
 FILLER_ASAP7_75t_R FILLER_138_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1167 ();
 DECAPx1_ASAP7_75t_R FILLER_138_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_138_1189 ();
 FILLER_ASAP7_75t_R FILLER_138_1199 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_138_1216 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_138_1238 ();
 FILLER_ASAP7_75t_R FILLER_138_1247 ();
 FILLER_ASAP7_75t_R FILLER_138_1257 ();
 DECAPx4_ASAP7_75t_R FILLER_138_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_1272 ();
 FILLER_ASAP7_75t_R FILLER_138_1279 ();
 DECAPx4_ASAP7_75t_R FILLER_138_1287 ();
 DECAPx4_ASAP7_75t_R FILLER_138_1303 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_138_1313 ();
 FILLER_ASAP7_75t_R FILLER_138_1325 ();
 FILLER_ASAP7_75t_R FILLER_138_1333 ();
 FILLER_ASAP7_75t_R FILLER_138_1342 ();
 DECAPx2_ASAP7_75t_R FILLER_138_1353 ();
 FILLER_ASAP7_75t_R FILLER_138_1359 ();
 FILLER_ASAP7_75t_R FILLER_138_1369 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_138_1374 ();
 FILLER_ASAP7_75t_R FILLER_139_2 ();
 DECAPx1_ASAP7_75t_R FILLER_139_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_13 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_20 ();
 DECAPx2_ASAP7_75t_R FILLER_139_26 ();
 FILLER_ASAP7_75t_R FILLER_139_35 ();
 DECAPx1_ASAP7_75t_R FILLER_139_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_47 ();
 DECAPx1_ASAP7_75t_R FILLER_139_51 ();
 FILLER_ASAP7_75t_R FILLER_139_61 ();
 DECAPx6_ASAP7_75t_R FILLER_139_71 ();
 DECAPx2_ASAP7_75t_R FILLER_139_85 ();
 DECAPx4_ASAP7_75t_R FILLER_139_94 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_104 ();
 FILLER_ASAP7_75t_R FILLER_139_113 ();
 DECAPx2_ASAP7_75t_R FILLER_139_118 ();
 FILLER_ASAP7_75t_R FILLER_139_124 ();
 FILLER_ASAP7_75t_R FILLER_139_152 ();
 DECAPx6_ASAP7_75t_R FILLER_139_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_194 ();
 DECAPx10_ASAP7_75t_R FILLER_139_198 ();
 DECAPx10_ASAP7_75t_R FILLER_139_220 ();
 DECAPx4_ASAP7_75t_R FILLER_139_242 ();
 FILLER_ASAP7_75t_R FILLER_139_252 ();
 FILLER_ASAP7_75t_R FILLER_139_260 ();
 DECAPx6_ASAP7_75t_R FILLER_139_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_279 ();
 FILLER_ASAP7_75t_R FILLER_139_295 ();
 FILLER_ASAP7_75t_R FILLER_139_323 ();
 DECAPx6_ASAP7_75t_R FILLER_139_331 ();
 DECAPx2_ASAP7_75t_R FILLER_139_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_351 ();
 DECAPx4_ASAP7_75t_R FILLER_139_358 ();
 FILLER_ASAP7_75t_R FILLER_139_371 ();
 DECAPx6_ASAP7_75t_R FILLER_139_381 ();
 DECAPx1_ASAP7_75t_R FILLER_139_421 ();
 DECAPx10_ASAP7_75t_R FILLER_139_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_453 ();
 DECAPx2_ASAP7_75t_R FILLER_139_460 ();
 FILLER_ASAP7_75t_R FILLER_139_472 ();
 FILLER_ASAP7_75t_R FILLER_139_481 ();
 FILLER_ASAP7_75t_R FILLER_139_489 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_497 ();
 FILLER_ASAP7_75t_R FILLER_139_503 ();
 DECAPx2_ASAP7_75t_R FILLER_139_513 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_519 ();
 FILLER_ASAP7_75t_R FILLER_139_528 ();
 FILLER_ASAP7_75t_R FILLER_139_537 ();
 FILLER_ASAP7_75t_R FILLER_139_549 ();
 DECAPx2_ASAP7_75t_R FILLER_139_559 ();
 FILLER_ASAP7_75t_R FILLER_139_565 ();
 FILLER_ASAP7_75t_R FILLER_139_575 ();
 DECAPx1_ASAP7_75t_R FILLER_139_583 ();
 DECAPx2_ASAP7_75t_R FILLER_139_601 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_607 ();
 FILLER_ASAP7_75t_R FILLER_139_618 ();
 DECAPx6_ASAP7_75t_R FILLER_139_630 ();
 FILLER_ASAP7_75t_R FILLER_139_652 ();
 DECAPx6_ASAP7_75t_R FILLER_139_661 ();
 DECAPx1_ASAP7_75t_R FILLER_139_675 ();
 DECAPx2_ASAP7_75t_R FILLER_139_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_691 ();
 DECAPx4_ASAP7_75t_R FILLER_139_698 ();
 DECAPx4_ASAP7_75t_R FILLER_139_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_724 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_740 ();
 FILLER_ASAP7_75t_R FILLER_139_750 ();
 FILLER_ASAP7_75t_R FILLER_139_758 ();
 DECAPx6_ASAP7_75t_R FILLER_139_766 ();
 DECAPx2_ASAP7_75t_R FILLER_139_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_786 ();
 FILLER_ASAP7_75t_R FILLER_139_796 ();
 DECAPx6_ASAP7_75t_R FILLER_139_805 ();
 FILLER_ASAP7_75t_R FILLER_139_819 ();
 DECAPx4_ASAP7_75t_R FILLER_139_828 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_838 ();
 FILLER_ASAP7_75t_R FILLER_139_844 ();
 DECAPx6_ASAP7_75t_R FILLER_139_854 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_868 ();
 DECAPx4_ASAP7_75t_R FILLER_139_877 ();
 DECAPx2_ASAP7_75t_R FILLER_139_901 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_907 ();
 DECAPx2_ASAP7_75t_R FILLER_139_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_924 ();
 FILLER_ASAP7_75t_R FILLER_139_927 ();
 DECAPx10_ASAP7_75t_R FILLER_139_933 ();
 DECAPx6_ASAP7_75t_R FILLER_139_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_969 ();
 DECAPx10_ASAP7_75t_R FILLER_139_977 ();
 DECAPx2_ASAP7_75t_R FILLER_139_999 ();
 FILLER_ASAP7_75t_R FILLER_139_1005 ();
 DECAPx4_ASAP7_75t_R FILLER_139_1010 ();
 FILLER_ASAP7_75t_R FILLER_139_1020 ();
 FILLER_ASAP7_75t_R FILLER_139_1028 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_1036 ();
 FILLER_ASAP7_75t_R FILLER_139_1045 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_1057 ();
 FILLER_ASAP7_75t_R FILLER_139_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1094 ();
 DECAPx1_ASAP7_75t_R FILLER_139_1116 ();
 DECAPx4_ASAP7_75t_R FILLER_139_1123 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_1133 ();
 FILLER_ASAP7_75t_R FILLER_139_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1147 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_1153 ();
 FILLER_ASAP7_75t_R FILLER_139_1162 ();
 FILLER_ASAP7_75t_R FILLER_139_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1200 ();
 FILLER_ASAP7_75t_R FILLER_139_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_139_1228 ();
 DECAPx6_ASAP7_75t_R FILLER_139_1250 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_1264 ();
 DECAPx6_ASAP7_75t_R FILLER_139_1276 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1290 ();
 FILLER_ASAP7_75t_R FILLER_139_1294 ();
 FILLER_ASAP7_75t_R FILLER_139_1305 ();
 DECAPx6_ASAP7_75t_R FILLER_139_1310 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_1324 ();
 DECAPx1_ASAP7_75t_R FILLER_139_1337 ();
 DECAPx4_ASAP7_75t_R FILLER_139_1344 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_1354 ();
 DECAPx2_ASAP7_75t_R FILLER_139_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_1369 ();
 FILLER_ASAP7_75t_R FILLER_139_1375 ();
 FILLER_ASAP7_75t_R FILLER_140_2 ();
 DECAPx6_ASAP7_75t_R FILLER_140_10 ();
 DECAPx2_ASAP7_75t_R FILLER_140_24 ();
 DECAPx10_ASAP7_75t_R FILLER_140_33 ();
 DECAPx1_ASAP7_75t_R FILLER_140_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_59 ();
 DECAPx10_ASAP7_75t_R FILLER_140_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_88 ();
 DECAPx10_ASAP7_75t_R FILLER_140_95 ();
 DECAPx6_ASAP7_75t_R FILLER_140_117 ();
 DECAPx1_ASAP7_75t_R FILLER_140_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_135 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_142 ();
 DECAPx2_ASAP7_75t_R FILLER_140_148 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_154 ();
 DECAPx4_ASAP7_75t_R FILLER_140_163 ();
 FILLER_ASAP7_75t_R FILLER_140_173 ();
 DECAPx4_ASAP7_75t_R FILLER_140_181 ();
 FILLER_ASAP7_75t_R FILLER_140_197 ();
 DECAPx6_ASAP7_75t_R FILLER_140_202 ();
 DECAPx2_ASAP7_75t_R FILLER_140_222 ();
 FILLER_ASAP7_75t_R FILLER_140_228 ();
 FILLER_ASAP7_75t_R FILLER_140_236 ();
 DECAPx4_ASAP7_75t_R FILLER_140_244 ();
 DECAPx2_ASAP7_75t_R FILLER_140_260 ();
 FILLER_ASAP7_75t_R FILLER_140_266 ();
 FILLER_ASAP7_75t_R FILLER_140_275 ();
 FILLER_ASAP7_75t_R FILLER_140_285 ();
 DECAPx2_ASAP7_75t_R FILLER_140_294 ();
 FILLER_ASAP7_75t_R FILLER_140_300 ();
 DECAPx1_ASAP7_75t_R FILLER_140_308 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_315 ();
 FILLER_ASAP7_75t_R FILLER_140_324 ();
 DECAPx4_ASAP7_75t_R FILLER_140_334 ();
 FILLER_ASAP7_75t_R FILLER_140_344 ();
 DECAPx6_ASAP7_75t_R FILLER_140_372 ();
 DECAPx2_ASAP7_75t_R FILLER_140_386 ();
 DECAPx1_ASAP7_75t_R FILLER_140_398 ();
 FILLER_ASAP7_75t_R FILLER_140_408 ();
 FILLER_ASAP7_75t_R FILLER_140_413 ();
 DECAPx6_ASAP7_75t_R FILLER_140_441 ();
 DECAPx2_ASAP7_75t_R FILLER_140_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_461 ();
 FILLER_ASAP7_75t_R FILLER_140_464 ();
 FILLER_ASAP7_75t_R FILLER_140_472 ();
 FILLER_ASAP7_75t_R FILLER_140_481 ();
 DECAPx2_ASAP7_75t_R FILLER_140_490 ();
 FILLER_ASAP7_75t_R FILLER_140_503 ();
 DECAPx6_ASAP7_75t_R FILLER_140_511 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_525 ();
 DECAPx10_ASAP7_75t_R FILLER_140_535 ();
 DECAPx4_ASAP7_75t_R FILLER_140_557 ();
 DECAPx6_ASAP7_75t_R FILLER_140_573 ();
 DECAPx1_ASAP7_75t_R FILLER_140_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_591 ();
 DECAPx6_ASAP7_75t_R FILLER_140_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_616 ();
 DECAPx2_ASAP7_75t_R FILLER_140_624 ();
 FILLER_ASAP7_75t_R FILLER_140_638 ();
 DECAPx2_ASAP7_75t_R FILLER_140_646 ();
 DECAPx2_ASAP7_75t_R FILLER_140_659 ();
 DECAPx6_ASAP7_75t_R FILLER_140_673 ();
 FILLER_ASAP7_75t_R FILLER_140_697 ();
 FILLER_ASAP7_75t_R FILLER_140_707 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_715 ();
 FILLER_ASAP7_75t_R FILLER_140_733 ();
 FILLER_ASAP7_75t_R FILLER_140_741 ();
 DECAPx4_ASAP7_75t_R FILLER_140_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_759 ();
 FILLER_ASAP7_75t_R FILLER_140_768 ();
 DECAPx1_ASAP7_75t_R FILLER_140_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_780 ();
 FILLER_ASAP7_75t_R FILLER_140_795 ();
 FILLER_ASAP7_75t_R FILLER_140_800 ();
 FILLER_ASAP7_75t_R FILLER_140_813 ();
 FILLER_ASAP7_75t_R FILLER_140_821 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_833 ();
 FILLER_ASAP7_75t_R FILLER_140_850 ();
 DECAPx2_ASAP7_75t_R FILLER_140_861 ();
 DECAPx2_ASAP7_75t_R FILLER_140_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_879 ();
 DECAPx1_ASAP7_75t_R FILLER_140_886 ();
 DECAPx4_ASAP7_75t_R FILLER_140_901 ();
 FILLER_ASAP7_75t_R FILLER_140_920 ();
 FILLER_ASAP7_75t_R FILLER_140_930 ();
 DECAPx2_ASAP7_75t_R FILLER_140_939 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_945 ();
 DECAPx1_ASAP7_75t_R FILLER_140_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_961 ();
 FILLER_ASAP7_75t_R FILLER_140_966 ();
 FILLER_ASAP7_75t_R FILLER_140_978 ();
 DECAPx1_ASAP7_75t_R FILLER_140_983 ();
 DECAPx1_ASAP7_75t_R FILLER_140_994 ();
 FILLER_ASAP7_75t_R FILLER_140_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1016 ();
 FILLER_ASAP7_75t_R FILLER_140_1022 ();
 DECAPx4_ASAP7_75t_R FILLER_140_1034 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1050 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_1072 ();
 DECAPx6_ASAP7_75t_R FILLER_140_1078 ();
 FILLER_ASAP7_75t_R FILLER_140_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_140_1097 ();
 DECAPx6_ASAP7_75t_R FILLER_140_1119 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1142 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1166 ();
 FILLER_ASAP7_75t_R FILLER_140_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1191 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1195 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_1201 ();
 FILLER_ASAP7_75t_R FILLER_140_1207 ();
 FILLER_ASAP7_75t_R FILLER_140_1218 ();
 FILLER_ASAP7_75t_R FILLER_140_1228 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1254 ();
 DECAPx2_ASAP7_75t_R FILLER_140_1263 ();
 DECAPx6_ASAP7_75t_R FILLER_140_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1286 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1293 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1297 ();
 FILLER_ASAP7_75t_R FILLER_140_1306 ();
 DECAPx6_ASAP7_75t_R FILLER_140_1334 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1348 ();
 DECAPx1_ASAP7_75t_R FILLER_140_1360 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_1364 ();
 FILLER_ASAP7_75t_R FILLER_140_1368 ();
 FILLER_ASAP7_75t_R FILLER_140_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_141_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_8 ();
 DECAPx2_ASAP7_75t_R FILLER_141_17 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_49 ();
 DECAPx6_ASAP7_75t_R FILLER_141_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_72 ();
 DECAPx2_ASAP7_75t_R FILLER_141_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_85 ();
 FILLER_ASAP7_75t_R FILLER_141_112 ();
 DECAPx2_ASAP7_75t_R FILLER_141_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_126 ();
 DECAPx6_ASAP7_75t_R FILLER_141_135 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_149 ();
 DECAPx2_ASAP7_75t_R FILLER_141_158 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_164 ();
 DECAPx1_ASAP7_75t_R FILLER_141_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_197 ();
 DECAPx1_ASAP7_75t_R FILLER_141_204 ();
 DECAPx2_ASAP7_75t_R FILLER_141_234 ();
 DECAPx2_ASAP7_75t_R FILLER_141_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_254 ();
 FILLER_ASAP7_75t_R FILLER_141_262 ();
 FILLER_ASAP7_75t_R FILLER_141_271 ();
 DECAPx6_ASAP7_75t_R FILLER_141_295 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_309 ();
 FILLER_ASAP7_75t_R FILLER_141_319 ();
 DECAPx2_ASAP7_75t_R FILLER_141_324 ();
 FILLER_ASAP7_75t_R FILLER_141_330 ();
 DECAPx4_ASAP7_75t_R FILLER_141_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_348 ();
 DECAPx2_ASAP7_75t_R FILLER_141_355 ();
 DECAPx6_ASAP7_75t_R FILLER_141_364 ();
 DECAPx2_ASAP7_75t_R FILLER_141_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_384 ();
 FILLER_ASAP7_75t_R FILLER_141_411 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_416 ();
 DECAPx1_ASAP7_75t_R FILLER_141_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_429 ();
 DECAPx6_ASAP7_75t_R FILLER_141_433 ();
 FILLER_ASAP7_75t_R FILLER_141_447 ();
 FILLER_ASAP7_75t_R FILLER_141_457 ();
 DECAPx2_ASAP7_75t_R FILLER_141_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_473 ();
 FILLER_ASAP7_75t_R FILLER_141_481 ();
 DECAPx2_ASAP7_75t_R FILLER_141_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_496 ();
 DECAPx10_ASAP7_75t_R FILLER_141_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_545 ();
 FILLER_ASAP7_75t_R FILLER_141_552 ();
 DECAPx4_ASAP7_75t_R FILLER_141_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_567 ();
 DECAPx4_ASAP7_75t_R FILLER_141_574 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_584 ();
 DECAPx6_ASAP7_75t_R FILLER_141_594 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_608 ();
 DECAPx4_ASAP7_75t_R FILLER_141_617 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_627 ();
 DECAPx2_ASAP7_75t_R FILLER_141_636 ();
 DECAPx4_ASAP7_75t_R FILLER_141_648 ();
 FILLER_ASAP7_75t_R FILLER_141_658 ();
 FILLER_ASAP7_75t_R FILLER_141_668 ();
 DECAPx10_ASAP7_75t_R FILLER_141_682 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_704 ();
 DECAPx10_ASAP7_75t_R FILLER_141_713 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_735 ();
 FILLER_ASAP7_75t_R FILLER_141_746 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_754 ();
 DECAPx1_ASAP7_75t_R FILLER_141_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_767 ();
 DECAPx2_ASAP7_75t_R FILLER_141_771 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_777 ();
 FILLER_ASAP7_75t_R FILLER_141_788 ();
 DECAPx10_ASAP7_75t_R FILLER_141_793 ();
 DECAPx6_ASAP7_75t_R FILLER_141_815 ();
 DECAPx2_ASAP7_75t_R FILLER_141_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_835 ();
 FILLER_ASAP7_75t_R FILLER_141_847 ();
 DECAPx2_ASAP7_75t_R FILLER_141_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_858 ();
 FILLER_ASAP7_75t_R FILLER_141_866 ();
 FILLER_ASAP7_75t_R FILLER_141_874 ();
 DECAPx2_ASAP7_75t_R FILLER_141_882 ();
 FILLER_ASAP7_75t_R FILLER_141_888 ();
 FILLER_ASAP7_75t_R FILLER_141_899 ();
 DECAPx6_ASAP7_75t_R FILLER_141_908 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_922 ();
 FILLER_ASAP7_75t_R FILLER_141_927 ();
 DECAPx4_ASAP7_75t_R FILLER_141_935 ();
 FILLER_ASAP7_75t_R FILLER_141_945 ();
 FILLER_ASAP7_75t_R FILLER_141_950 ();
 DECAPx4_ASAP7_75t_R FILLER_141_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_968 ();
 DECAPx4_ASAP7_75t_R FILLER_141_975 ();
 FILLER_ASAP7_75t_R FILLER_141_989 ();
 DECAPx10_ASAP7_75t_R FILLER_141_997 ();
 FILLER_ASAP7_75t_R FILLER_141_1019 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1027 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_1037 ();
 FILLER_ASAP7_75t_R FILLER_141_1046 ();
 DECAPx6_ASAP7_75t_R FILLER_141_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1068 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1092 ();
 FILLER_ASAP7_75t_R FILLER_141_1096 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1106 ();
 FILLER_ASAP7_75t_R FILLER_141_1124 ();
 FILLER_ASAP7_75t_R FILLER_141_1132 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1140 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1155 ();
 FILLER_ASAP7_75t_R FILLER_141_1165 ();
 FILLER_ASAP7_75t_R FILLER_141_1193 ();
 FILLER_ASAP7_75t_R FILLER_141_1221 ();
 FILLER_ASAP7_75t_R FILLER_141_1229 ();
 FILLER_ASAP7_75t_R FILLER_141_1257 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_141_1273 ();
 DECAPx4_ASAP7_75t_R FILLER_141_1295 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1305 ();
 DECAPx2_ASAP7_75t_R FILLER_141_1314 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_1320 ();
 DECAPx6_ASAP7_75t_R FILLER_141_1326 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_1340 ();
 FILLER_ASAP7_75t_R FILLER_141_1347 ();
 FILLER_ASAP7_75t_R FILLER_141_1375 ();
 FILLER_ASAP7_75t_R FILLER_142_2 ();
 DECAPx1_ASAP7_75t_R FILLER_142_30 ();
 DECAPx1_ASAP7_75t_R FILLER_142_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_44 ();
 FILLER_ASAP7_75t_R FILLER_142_71 ();
 FILLER_ASAP7_75t_R FILLER_142_81 ();
 DECAPx1_ASAP7_75t_R FILLER_142_89 ();
 DECAPx1_ASAP7_75t_R FILLER_142_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_103 ();
 FILLER_ASAP7_75t_R FILLER_142_130 ();
 FILLER_ASAP7_75t_R FILLER_142_142 ();
 DECAPx6_ASAP7_75t_R FILLER_142_150 ();
 DECAPx2_ASAP7_75t_R FILLER_142_164 ();
 DECAPx1_ASAP7_75t_R FILLER_142_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_180 ();
 DECAPx1_ASAP7_75t_R FILLER_142_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_188 ();
 FILLER_ASAP7_75t_R FILLER_142_195 ();
 DECAPx2_ASAP7_75t_R FILLER_142_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_211 ();
 DECAPx1_ASAP7_75t_R FILLER_142_218 ();
 DECAPx4_ASAP7_75t_R FILLER_142_225 ();
 FILLER_ASAP7_75t_R FILLER_142_241 ();
 DECAPx1_ASAP7_75t_R FILLER_142_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_250 ();
 FILLER_ASAP7_75t_R FILLER_142_277 ();
 DECAPx1_ASAP7_75t_R FILLER_142_286 ();
 DECAPx6_ASAP7_75t_R FILLER_142_316 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_142_330 ();
 DECAPx6_ASAP7_75t_R FILLER_142_339 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_142_353 ();
 DECAPx2_ASAP7_75t_R FILLER_142_362 ();
 DECAPx6_ASAP7_75t_R FILLER_142_371 ();
 FILLER_ASAP7_75t_R FILLER_142_385 ();
 DECAPx1_ASAP7_75t_R FILLER_142_393 ();
 DECAPx6_ASAP7_75t_R FILLER_142_415 ();
 DECAPx1_ASAP7_75t_R FILLER_142_429 ();
 FILLER_ASAP7_75t_R FILLER_142_440 ();
 DECAPx2_ASAP7_75t_R FILLER_142_448 ();
 FILLER_ASAP7_75t_R FILLER_142_460 ();
 FILLER_ASAP7_75t_R FILLER_142_464 ();
 DECAPx2_ASAP7_75t_R FILLER_142_476 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_142_482 ();
 DECAPx1_ASAP7_75t_R FILLER_142_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_499 ();
 DECAPx2_ASAP7_75t_R FILLER_142_506 ();
 DECAPx10_ASAP7_75t_R FILLER_142_515 ();
 DECAPx2_ASAP7_75t_R FILLER_142_537 ();
 DECAPx2_ASAP7_75t_R FILLER_142_550 ();
 DECAPx6_ASAP7_75t_R FILLER_142_559 ();
 DECAPx2_ASAP7_75t_R FILLER_142_573 ();
 DECAPx6_ASAP7_75t_R FILLER_142_585 ();
 FILLER_ASAP7_75t_R FILLER_142_607 ();
 DECAPx10_ASAP7_75t_R FILLER_142_615 ();
 DECAPx10_ASAP7_75t_R FILLER_142_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_659 ();
 FILLER_ASAP7_75t_R FILLER_142_666 ();
 DECAPx4_ASAP7_75t_R FILLER_142_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_684 ();
 DECAPx10_ASAP7_75t_R FILLER_142_693 ();
 DECAPx10_ASAP7_75t_R FILLER_142_715 ();
 DECAPx4_ASAP7_75t_R FILLER_142_737 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_142_747 ();
 DECAPx1_ASAP7_75t_R FILLER_142_756 ();
 DECAPx1_ASAP7_75t_R FILLER_142_767 ();
 DECAPx4_ASAP7_75t_R FILLER_142_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_788 ();
 DECAPx10_ASAP7_75t_R FILLER_142_797 ();
 DECAPx10_ASAP7_75t_R FILLER_142_819 ();
 DECAPx6_ASAP7_75t_R FILLER_142_841 ();
 FILLER_ASAP7_75t_R FILLER_142_855 ();
 FILLER_ASAP7_75t_R FILLER_142_863 ();
 DECAPx10_ASAP7_75t_R FILLER_142_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_897 ();
 FILLER_ASAP7_75t_R FILLER_142_905 ();
 DECAPx4_ASAP7_75t_R FILLER_142_914 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_142_930 ();
 DECAPx2_ASAP7_75t_R FILLER_142_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_949 ();
 FILLER_ASAP7_75t_R FILLER_142_958 ();
 DECAPx4_ASAP7_75t_R FILLER_142_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_973 ();
 DECAPx6_ASAP7_75t_R FILLER_142_980 ();
 DECAPx1_ASAP7_75t_R FILLER_142_994 ();
 DECAPx4_ASAP7_75t_R FILLER_142_1004 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_142_1014 ();
 FILLER_ASAP7_75t_R FILLER_142_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_142_1035 ();
 FILLER_ASAP7_75t_R FILLER_142_1042 ();
 DECAPx6_ASAP7_75t_R FILLER_142_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1068 ();
 FILLER_ASAP7_75t_R FILLER_142_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_142_1139 ();
 DECAPx6_ASAP7_75t_R FILLER_142_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1181 ();
 FILLER_ASAP7_75t_R FILLER_142_1185 ();
 DECAPx1_ASAP7_75t_R FILLER_142_1191 ();
 FILLER_ASAP7_75t_R FILLER_142_1201 ();
 DECAPx1_ASAP7_75t_R FILLER_142_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1210 ();
 DECAPx6_ASAP7_75t_R FILLER_142_1219 ();
 DECAPx6_ASAP7_75t_R FILLER_142_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1255 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_142_1282 ();
 FILLER_ASAP7_75t_R FILLER_142_1293 ();
 DECAPx6_ASAP7_75t_R FILLER_142_1303 ();
 DECAPx4_ASAP7_75t_R FILLER_142_1323 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_142_1333 ();
 DECAPx4_ASAP7_75t_R FILLER_142_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1354 ();
 DECAPx2_ASAP7_75t_R FILLER_142_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_1369 ();
 FILLER_ASAP7_75t_R FILLER_142_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_143_2 ();
 FILLER_ASAP7_75t_R FILLER_143_14 ();
 FILLER_ASAP7_75t_R FILLER_143_21 ();
 FILLER_ASAP7_75t_R FILLER_143_26 ();
 DECAPx1_ASAP7_75t_R FILLER_143_34 ();
 DECAPx2_ASAP7_75t_R FILLER_143_41 ();
 FILLER_ASAP7_75t_R FILLER_143_47 ();
 DECAPx1_ASAP7_75t_R FILLER_143_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_59 ();
 DECAPx2_ASAP7_75t_R FILLER_143_63 ();
 FILLER_ASAP7_75t_R FILLER_143_75 ();
 DECAPx6_ASAP7_75t_R FILLER_143_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_99 ();
 DECAPx2_ASAP7_75t_R FILLER_143_103 ();
 FILLER_ASAP7_75t_R FILLER_143_109 ();
 FILLER_ASAP7_75t_R FILLER_143_117 ();
 DECAPx2_ASAP7_75t_R FILLER_143_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_128 ();
 FILLER_ASAP7_75t_R FILLER_143_135 ();
 DECAPx6_ASAP7_75t_R FILLER_143_163 ();
 DECAPx1_ASAP7_75t_R FILLER_143_177 ();
 DECAPx2_ASAP7_75t_R FILLER_143_191 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_197 ();
 DECAPx6_ASAP7_75t_R FILLER_143_206 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_226 ();
 DECAPx10_ASAP7_75t_R FILLER_143_235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_263 ();
 DECAPx1_ASAP7_75t_R FILLER_143_272 ();
 FILLER_ASAP7_75t_R FILLER_143_283 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_291 ();
 DECAPx1_ASAP7_75t_R FILLER_143_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_304 ();
 DECAPx6_ASAP7_75t_R FILLER_143_308 ();
 DECAPx2_ASAP7_75t_R FILLER_143_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_328 ();
 FILLER_ASAP7_75t_R FILLER_143_337 ();
 DECAPx2_ASAP7_75t_R FILLER_143_347 ();
 DECAPx1_ASAP7_75t_R FILLER_143_379 ();
 DECAPx6_ASAP7_75t_R FILLER_143_389 ();
 DECAPx1_ASAP7_75t_R FILLER_143_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_413 ();
 DECAPx2_ASAP7_75t_R FILLER_143_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_426 ();
 FILLER_ASAP7_75t_R FILLER_143_453 ();
 DECAPx6_ASAP7_75t_R FILLER_143_458 ();
 FILLER_ASAP7_75t_R FILLER_143_472 ();
 FILLER_ASAP7_75t_R FILLER_143_481 ();
 FILLER_ASAP7_75t_R FILLER_143_495 ();
 DECAPx1_ASAP7_75t_R FILLER_143_504 ();
 FILLER_ASAP7_75t_R FILLER_143_516 ();
 FILLER_ASAP7_75t_R FILLER_143_526 ();
 DECAPx1_ASAP7_75t_R FILLER_143_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_540 ();
 DECAPx1_ASAP7_75t_R FILLER_143_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_571 ();
 FILLER_ASAP7_75t_R FILLER_143_578 ();
 DECAPx2_ASAP7_75t_R FILLER_143_587 ();
 FILLER_ASAP7_75t_R FILLER_143_603 ();
 FILLER_ASAP7_75t_R FILLER_143_611 ();
 DECAPx1_ASAP7_75t_R FILLER_143_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_623 ();
 DECAPx1_ASAP7_75t_R FILLER_143_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_636 ();
 FILLER_ASAP7_75t_R FILLER_143_643 ();
 DECAPx6_ASAP7_75t_R FILLER_143_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_666 ();
 DECAPx4_ASAP7_75t_R FILLER_143_673 ();
 FILLER_ASAP7_75t_R FILLER_143_689 ();
 DECAPx2_ASAP7_75t_R FILLER_143_697 ();
 FILLER_ASAP7_75t_R FILLER_143_713 ();
 DECAPx2_ASAP7_75t_R FILLER_143_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_727 ();
 DECAPx4_ASAP7_75t_R FILLER_143_736 ();
 FILLER_ASAP7_75t_R FILLER_143_746 ();
 FILLER_ASAP7_75t_R FILLER_143_756 ();
 FILLER_ASAP7_75t_R FILLER_143_766 ();
 FILLER_ASAP7_75t_R FILLER_143_774 ();
 DECAPx1_ASAP7_75t_R FILLER_143_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_790 ();
 DECAPx6_ASAP7_75t_R FILLER_143_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_815 ();
 DECAPx1_ASAP7_75t_R FILLER_143_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_830 ();
 DECAPx6_ASAP7_75t_R FILLER_143_837 ();
 DECAPx1_ASAP7_75t_R FILLER_143_851 ();
 DECAPx4_ASAP7_75t_R FILLER_143_864 ();
 DECAPx4_ASAP7_75t_R FILLER_143_880 ();
 DECAPx10_ASAP7_75t_R FILLER_143_897 ();
 DECAPx2_ASAP7_75t_R FILLER_143_919 ();
 DECAPx1_ASAP7_75t_R FILLER_143_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_931 ();
 DECAPx2_ASAP7_75t_R FILLER_143_937 ();
 FILLER_ASAP7_75t_R FILLER_143_943 ();
 FILLER_ASAP7_75t_R FILLER_143_954 ();
 DECAPx1_ASAP7_75t_R FILLER_143_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_966 ();
 DECAPx6_ASAP7_75t_R FILLER_143_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_992 ();
 FILLER_ASAP7_75t_R FILLER_143_1002 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1023 ();
 DECAPx6_ASAP7_75t_R FILLER_143_1032 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_1046 ();
 FILLER_ASAP7_75t_R FILLER_143_1058 ();
 DECAPx4_ASAP7_75t_R FILLER_143_1070 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_1080 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_1086 ();
 DECAPx6_ASAP7_75t_R FILLER_143_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1109 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_143_1130 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1152 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_143_1177 ();
 DECAPx4_ASAP7_75t_R FILLER_143_1199 ();
 FILLER_ASAP7_75t_R FILLER_143_1209 ();
 DECAPx6_ASAP7_75t_R FILLER_143_1214 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1234 ();
 FILLER_ASAP7_75t_R FILLER_143_1241 ();
 DECAPx4_ASAP7_75t_R FILLER_143_1249 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_143_1270 ();
 FILLER_ASAP7_75t_R FILLER_143_1280 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1308 ();
 FILLER_ASAP7_75t_R FILLER_143_1314 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1326 ();
 FILLER_ASAP7_75t_R FILLER_143_1336 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1344 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_1350 ();
 DECAPx1_ASAP7_75t_R FILLER_143_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_1365 ();
 DECAPx2_ASAP7_75t_R FILLER_143_1369 ();
 FILLER_ASAP7_75t_R FILLER_143_1375 ();
 FILLER_ASAP7_75t_R FILLER_144_2 ();
 DECAPx2_ASAP7_75t_R FILLER_144_10 ();
 DECAPx6_ASAP7_75t_R FILLER_144_22 ();
 DECAPx1_ASAP7_75t_R FILLER_144_36 ();
 DECAPx10_ASAP7_75t_R FILLER_144_46 ();
 DECAPx6_ASAP7_75t_R FILLER_144_68 ();
 DECAPx2_ASAP7_75t_R FILLER_144_82 ();
 DECAPx6_ASAP7_75t_R FILLER_144_96 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_110 ();
 DECAPx10_ASAP7_75t_R FILLER_144_116 ();
 DECAPx1_ASAP7_75t_R FILLER_144_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_142 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_149 ();
 FILLER_ASAP7_75t_R FILLER_144_155 ();
 DECAPx6_ASAP7_75t_R FILLER_144_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_181 ();
 DECAPx2_ASAP7_75t_R FILLER_144_188 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_194 ();
 DECAPx6_ASAP7_75t_R FILLER_144_203 ();
 DECAPx10_ASAP7_75t_R FILLER_144_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_265 ();
 FILLER_ASAP7_75t_R FILLER_144_272 ();
 FILLER_ASAP7_75t_R FILLER_144_280 ();
 DECAPx6_ASAP7_75t_R FILLER_144_285 ();
 DECAPx1_ASAP7_75t_R FILLER_144_305 ();
 DECAPx2_ASAP7_75t_R FILLER_144_315 ();
 DECAPx2_ASAP7_75t_R FILLER_144_324 ();
 FILLER_ASAP7_75t_R FILLER_144_330 ();
 DECAPx6_ASAP7_75t_R FILLER_144_338 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_352 ();
 DECAPx2_ASAP7_75t_R FILLER_144_361 ();
 FILLER_ASAP7_75t_R FILLER_144_367 ();
 DECAPx2_ASAP7_75t_R FILLER_144_395 ();
 FILLER_ASAP7_75t_R FILLER_144_401 ();
 DECAPx1_ASAP7_75t_R FILLER_144_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_413 ();
 DECAPx6_ASAP7_75t_R FILLER_144_422 ();
 DECAPx2_ASAP7_75t_R FILLER_144_436 ();
 DECAPx2_ASAP7_75t_R FILLER_144_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_451 ();
 FILLER_ASAP7_75t_R FILLER_144_460 ();
 FILLER_ASAP7_75t_R FILLER_144_464 ();
 DECAPx1_ASAP7_75t_R FILLER_144_472 ();
 DECAPx10_ASAP7_75t_R FILLER_144_482 ();
 DECAPx4_ASAP7_75t_R FILLER_144_504 ();
 FILLER_ASAP7_75t_R FILLER_144_522 ();
 FILLER_ASAP7_75t_R FILLER_144_530 ();
 DECAPx6_ASAP7_75t_R FILLER_144_538 ();
 DECAPx2_ASAP7_75t_R FILLER_144_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_558 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_567 ();
 DECAPx10_ASAP7_75t_R FILLER_144_576 ();
 DECAPx2_ASAP7_75t_R FILLER_144_598 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_604 ();
 FILLER_ASAP7_75t_R FILLER_144_615 ();
 FILLER_ASAP7_75t_R FILLER_144_629 ();
 DECAPx2_ASAP7_75t_R FILLER_144_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_645 ();
 FILLER_ASAP7_75t_R FILLER_144_652 ();
 DECAPx1_ASAP7_75t_R FILLER_144_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_666 ();
 DECAPx2_ASAP7_75t_R FILLER_144_674 ();
 FILLER_ASAP7_75t_R FILLER_144_680 ();
 FILLER_ASAP7_75t_R FILLER_144_688 ();
 DECAPx2_ASAP7_75t_R FILLER_144_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_702 ();
 DECAPx2_ASAP7_75t_R FILLER_144_711 ();
 FILLER_ASAP7_75t_R FILLER_144_723 ();
 FILLER_ASAP7_75t_R FILLER_144_733 ();
 FILLER_ASAP7_75t_R FILLER_144_742 ();
 DECAPx10_ASAP7_75t_R FILLER_144_750 ();
 DECAPx10_ASAP7_75t_R FILLER_144_772 ();
 DECAPx2_ASAP7_75t_R FILLER_144_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_800 ();
 FILLER_ASAP7_75t_R FILLER_144_807 ();
 FILLER_ASAP7_75t_R FILLER_144_818 ();
 FILLER_ASAP7_75t_R FILLER_144_823 ();
 DECAPx1_ASAP7_75t_R FILLER_144_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_855 ();
 DECAPx6_ASAP7_75t_R FILLER_144_864 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_878 ();
 DECAPx1_ASAP7_75t_R FILLER_144_889 ();
 DECAPx2_ASAP7_75t_R FILLER_144_899 ();
 DECAPx2_ASAP7_75t_R FILLER_144_919 ();
 FILLER_ASAP7_75t_R FILLER_144_925 ();
 FILLER_ASAP7_75t_R FILLER_144_934 ();
 DECAPx6_ASAP7_75t_R FILLER_144_943 ();
 DECAPx1_ASAP7_75t_R FILLER_144_965 ();
 DECAPx2_ASAP7_75t_R FILLER_144_983 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_989 ();
 DECAPx1_ASAP7_75t_R FILLER_144_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_999 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1013 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1035 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1049 ();
 FILLER_ASAP7_75t_R FILLER_144_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1067 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1084 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1098 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1120 ();
 FILLER_ASAP7_75t_R FILLER_144_1143 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1157 ();
 DECAPx1_ASAP7_75t_R FILLER_144_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1176 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1230 ();
 DECAPx4_ASAP7_75t_R FILLER_144_1252 ();
 FILLER_ASAP7_75t_R FILLER_144_1262 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1270 ();
 FILLER_ASAP7_75t_R FILLER_144_1284 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1289 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_1295 ();
 DECAPx2_ASAP7_75t_R FILLER_144_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_144_1313 ();
 DECAPx6_ASAP7_75t_R FILLER_144_1335 ();
 FILLER_ASAP7_75t_R FILLER_144_1375 ();
 DECAPx1_ASAP7_75t_R FILLER_145_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_6 ();
 DECAPx2_ASAP7_75t_R FILLER_145_33 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_39 ();
 FILLER_ASAP7_75t_R FILLER_145_50 ();
 DECAPx4_ASAP7_75t_R FILLER_145_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_68 ();
 DECAPx6_ASAP7_75t_R FILLER_145_75 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_89 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_102 ();
 DECAPx1_ASAP7_75t_R FILLER_145_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_115 ();
 FILLER_ASAP7_75t_R FILLER_145_124 ();
 DECAPx6_ASAP7_75t_R FILLER_145_132 ();
 DECAPx2_ASAP7_75t_R FILLER_145_146 ();
 DECAPx1_ASAP7_75t_R FILLER_145_155 ();
 DECAPx2_ASAP7_75t_R FILLER_145_165 ();
 DECAPx1_ASAP7_75t_R FILLER_145_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_181 ();
 DECAPx1_ASAP7_75t_R FILLER_145_188 ();
 FILLER_ASAP7_75t_R FILLER_145_195 ();
 DECAPx4_ASAP7_75t_R FILLER_145_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_215 ();
 DECAPx1_ASAP7_75t_R FILLER_145_222 ();
 FILLER_ASAP7_75t_R FILLER_145_232 ();
 DECAPx1_ASAP7_75t_R FILLER_145_237 ();
 DECAPx1_ASAP7_75t_R FILLER_145_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_271 ();
 FILLER_ASAP7_75t_R FILLER_145_278 ();
 DECAPx4_ASAP7_75t_R FILLER_145_283 ();
 DECAPx1_ASAP7_75t_R FILLER_145_319 ();
 FILLER_ASAP7_75t_R FILLER_145_329 ();
 DECAPx6_ASAP7_75t_R FILLER_145_337 ();
 DECAPx6_ASAP7_75t_R FILLER_145_357 ();
 DECAPx1_ASAP7_75t_R FILLER_145_371 ();
 FILLER_ASAP7_75t_R FILLER_145_381 ();
 DECAPx1_ASAP7_75t_R FILLER_145_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_390 ();
 DECAPx6_ASAP7_75t_R FILLER_145_394 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_408 ();
 DECAPx6_ASAP7_75t_R FILLER_145_414 ();
 FILLER_ASAP7_75t_R FILLER_145_434 ();
 DECAPx4_ASAP7_75t_R FILLER_145_439 ();
 FILLER_ASAP7_75t_R FILLER_145_455 ();
 DECAPx1_ASAP7_75t_R FILLER_145_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_467 ();
 FILLER_ASAP7_75t_R FILLER_145_478 ();
 DECAPx4_ASAP7_75t_R FILLER_145_490 ();
 FILLER_ASAP7_75t_R FILLER_145_500 ();
 FILLER_ASAP7_75t_R FILLER_145_505 ();
 FILLER_ASAP7_75t_R FILLER_145_513 ();
 DECAPx10_ASAP7_75t_R FILLER_145_521 ();
 FILLER_ASAP7_75t_R FILLER_145_543 ();
 DECAPx6_ASAP7_75t_R FILLER_145_551 ();
 FILLER_ASAP7_75t_R FILLER_145_565 ();
 DECAPx4_ASAP7_75t_R FILLER_145_573 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_583 ();
 DECAPx4_ASAP7_75t_R FILLER_145_592 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_602 ();
 DECAPx6_ASAP7_75t_R FILLER_145_611 ();
 DECAPx1_ASAP7_75t_R FILLER_145_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_629 ();
 DECAPx1_ASAP7_75t_R FILLER_145_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_641 ();
 DECAPx2_ASAP7_75t_R FILLER_145_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_660 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_667 ();
 DECAPx10_ASAP7_75t_R FILLER_145_677 ();
 DECAPx1_ASAP7_75t_R FILLER_145_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_703 ();
 FILLER_ASAP7_75t_R FILLER_145_712 ();
 DECAPx1_ASAP7_75t_R FILLER_145_720 ();
 DECAPx6_ASAP7_75t_R FILLER_145_730 ();
 DECAPx2_ASAP7_75t_R FILLER_145_744 ();
 DECAPx6_ASAP7_75t_R FILLER_145_758 ();
 DECAPx2_ASAP7_75t_R FILLER_145_772 ();
 FILLER_ASAP7_75t_R FILLER_145_784 ();
 DECAPx2_ASAP7_75t_R FILLER_145_789 ();
 FILLER_ASAP7_75t_R FILLER_145_795 ();
 DECAPx1_ASAP7_75t_R FILLER_145_806 ();
 FILLER_ASAP7_75t_R FILLER_145_818 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_826 ();
 DECAPx1_ASAP7_75t_R FILLER_145_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_839 ();
 DECAPx2_ASAP7_75t_R FILLER_145_843 ();
 FILLER_ASAP7_75t_R FILLER_145_849 ();
 DECAPx4_ASAP7_75t_R FILLER_145_858 ();
 FILLER_ASAP7_75t_R FILLER_145_868 ();
 DECAPx6_ASAP7_75t_R FILLER_145_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_891 ();
 DECAPx2_ASAP7_75t_R FILLER_145_901 ();
 DECAPx2_ASAP7_75t_R FILLER_145_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_924 ();
 DECAPx2_ASAP7_75t_R FILLER_145_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_933 ();
 DECAPx10_ASAP7_75t_R FILLER_145_940 ();
 FILLER_ASAP7_75t_R FILLER_145_962 ();
 DECAPx4_ASAP7_75t_R FILLER_145_971 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_981 ();
 DECAPx6_ASAP7_75t_R FILLER_145_990 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_1004 ();
 FILLER_ASAP7_75t_R FILLER_145_1016 ();
 DECAPx6_ASAP7_75t_R FILLER_145_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1095 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_1101 ();
 FILLER_ASAP7_75t_R FILLER_145_1110 ();
 FILLER_ASAP7_75t_R FILLER_145_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1138 ();
 DECAPx4_ASAP7_75t_R FILLER_145_1165 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_1175 ();
 FILLER_ASAP7_75t_R FILLER_145_1204 ();
 FILLER_ASAP7_75t_R FILLER_145_1212 ();
 FILLER_ASAP7_75t_R FILLER_145_1217 ();
 FILLER_ASAP7_75t_R FILLER_145_1228 ();
 FILLER_ASAP7_75t_R FILLER_145_1256 ();
 FILLER_ASAP7_75t_R FILLER_145_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_145_1272 ();
 FILLER_ASAP7_75t_R FILLER_145_1278 ();
 FILLER_ASAP7_75t_R FILLER_145_1283 ();
 DECAPx1_ASAP7_75t_R FILLER_145_1294 ();
 FILLER_ASAP7_75t_R FILLER_145_1304 ();
 DECAPx4_ASAP7_75t_R FILLER_145_1332 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_1342 ();
 FILLER_ASAP7_75t_R FILLER_145_1346 ();
 FILLER_ASAP7_75t_R FILLER_145_1357 ();
 DECAPx4_ASAP7_75t_R FILLER_145_1367 ();
 DECAPx2_ASAP7_75t_R FILLER_146_2 ();
 FILLER_ASAP7_75t_R FILLER_146_8 ();
 FILLER_ASAP7_75t_R FILLER_146_16 ();
 FILLER_ASAP7_75t_R FILLER_146_24 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_31 ();
 FILLER_ASAP7_75t_R FILLER_146_37 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_42 ();
 DECAPx2_ASAP7_75t_R FILLER_146_53 ();
 FILLER_ASAP7_75t_R FILLER_146_59 ();
 DECAPx2_ASAP7_75t_R FILLER_146_87 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_93 ();
 FILLER_ASAP7_75t_R FILLER_146_102 ();
 DECAPx4_ASAP7_75t_R FILLER_146_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_117 ();
 DECAPx4_ASAP7_75t_R FILLER_146_126 ();
 FILLER_ASAP7_75t_R FILLER_146_136 ();
 DECAPx6_ASAP7_75t_R FILLER_146_148 ();
 DECAPx2_ASAP7_75t_R FILLER_146_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_168 ();
 DECAPx6_ASAP7_75t_R FILLER_146_195 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_209 ();
 FILLER_ASAP7_75t_R FILLER_146_238 ();
 FILLER_ASAP7_75t_R FILLER_146_246 ();
 DECAPx2_ASAP7_75t_R FILLER_146_254 ();
 DECAPx2_ASAP7_75t_R FILLER_146_286 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_292 ();
 DECAPx2_ASAP7_75t_R FILLER_146_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_307 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_311 ();
 FILLER_ASAP7_75t_R FILLER_146_340 ();
 DECAPx2_ASAP7_75t_R FILLER_146_368 ();
 DECAPx6_ASAP7_75t_R FILLER_146_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_394 ();
 FILLER_ASAP7_75t_R FILLER_146_403 ();
 FILLER_ASAP7_75t_R FILLER_146_419 ();
 FILLER_ASAP7_75t_R FILLER_146_427 ();
 FILLER_ASAP7_75t_R FILLER_146_435 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_459 ();
 DECAPx6_ASAP7_75t_R FILLER_146_464 ();
 DECAPx2_ASAP7_75t_R FILLER_146_478 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_494 ();
 FILLER_ASAP7_75t_R FILLER_146_504 ();
 DECAPx6_ASAP7_75t_R FILLER_146_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_523 ();
 DECAPx2_ASAP7_75t_R FILLER_146_530 ();
 FILLER_ASAP7_75t_R FILLER_146_539 ();
 DECAPx2_ASAP7_75t_R FILLER_146_567 ();
 FILLER_ASAP7_75t_R FILLER_146_580 ();
 DECAPx2_ASAP7_75t_R FILLER_146_597 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_603 ();
 FILLER_ASAP7_75t_R FILLER_146_612 ();
 DECAPx4_ASAP7_75t_R FILLER_146_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_630 ();
 DECAPx10_ASAP7_75t_R FILLER_146_637 ();
 DECAPx10_ASAP7_75t_R FILLER_146_659 ();
 DECAPx1_ASAP7_75t_R FILLER_146_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_685 ();
 DECAPx10_ASAP7_75t_R FILLER_146_692 ();
 DECAPx2_ASAP7_75t_R FILLER_146_714 ();
 FILLER_ASAP7_75t_R FILLER_146_720 ();
 DECAPx6_ASAP7_75t_R FILLER_146_728 ();
 DECAPx1_ASAP7_75t_R FILLER_146_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_746 ();
 DECAPx6_ASAP7_75t_R FILLER_146_753 ();
 FILLER_ASAP7_75t_R FILLER_146_773 ();
 FILLER_ASAP7_75t_R FILLER_146_789 ();
 FILLER_ASAP7_75t_R FILLER_146_801 ();
 DECAPx10_ASAP7_75t_R FILLER_146_806 ();
 DECAPx10_ASAP7_75t_R FILLER_146_828 ();
 DECAPx6_ASAP7_75t_R FILLER_146_850 ();
 DECAPx6_ASAP7_75t_R FILLER_146_873 ();
 DECAPx1_ASAP7_75t_R FILLER_146_887 ();
 FILLER_ASAP7_75t_R FILLER_146_898 ();
 FILLER_ASAP7_75t_R FILLER_146_906 ();
 FILLER_ASAP7_75t_R FILLER_146_911 ();
 DECAPx1_ASAP7_75t_R FILLER_146_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_920 ();
 DECAPx2_ASAP7_75t_R FILLER_146_929 ();
 FILLER_ASAP7_75t_R FILLER_146_943 ();
 DECAPx6_ASAP7_75t_R FILLER_146_953 ();
 FILLER_ASAP7_75t_R FILLER_146_967 ();
 DECAPx2_ASAP7_75t_R FILLER_146_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_984 ();
 DECAPx2_ASAP7_75t_R FILLER_146_994 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_1000 ();
 DECAPx4_ASAP7_75t_R FILLER_146_1012 ();
 FILLER_ASAP7_75t_R FILLER_146_1030 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1038 ();
 FILLER_ASAP7_75t_R FILLER_146_1053 ();
 FILLER_ASAP7_75t_R FILLER_146_1059 ();
 DECAPx6_ASAP7_75t_R FILLER_146_1064 ();
 FILLER_ASAP7_75t_R FILLER_146_1078 ();
 FILLER_ASAP7_75t_R FILLER_146_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1091 ();
 FILLER_ASAP7_75t_R FILLER_146_1105 ();
 FILLER_ASAP7_75t_R FILLER_146_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1125 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_1131 ();
 FILLER_ASAP7_75t_R FILLER_146_1137 ();
 FILLER_ASAP7_75t_R FILLER_146_1147 ();
 FILLER_ASAP7_75t_R FILLER_146_1152 ();
 DECAPx6_ASAP7_75t_R FILLER_146_1157 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1171 ();
 FILLER_ASAP7_75t_R FILLER_146_1185 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_1193 ();
 FILLER_ASAP7_75t_R FILLER_146_1206 ();
 FILLER_ASAP7_75t_R FILLER_146_1218 ();
 FILLER_ASAP7_75t_R FILLER_146_1226 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1234 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_1240 ();
 FILLER_ASAP7_75t_R FILLER_146_1249 ();
 FILLER_ASAP7_75t_R FILLER_146_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_146_1262 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1276 ();
 FILLER_ASAP7_75t_R FILLER_146_1286 ();
 FILLER_ASAP7_75t_R FILLER_146_1294 ();
 FILLER_ASAP7_75t_R FILLER_146_1302 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1314 ();
 DECAPx1_ASAP7_75t_R FILLER_146_1323 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1327 ();
 DECAPx4_ASAP7_75t_R FILLER_146_1338 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_1351 ();
 FILLER_ASAP7_75t_R FILLER_146_1360 ();
 DECAPx2_ASAP7_75t_R FILLER_146_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_1376 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_147_2 ();
 DECAPx6_ASAP7_75t_R FILLER_147_31 ();
 DECAPx2_ASAP7_75t_R FILLER_147_45 ();
 DECAPx2_ASAP7_75t_R FILLER_147_57 ();
 FILLER_ASAP7_75t_R FILLER_147_63 ();
 FILLER_ASAP7_75t_R FILLER_147_71 ();
 FILLER_ASAP7_75t_R FILLER_147_79 ();
 DECAPx1_ASAP7_75t_R FILLER_147_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_88 ();
 FILLER_ASAP7_75t_R FILLER_147_95 ();
 FILLER_ASAP7_75t_R FILLER_147_103 ();
 DECAPx4_ASAP7_75t_R FILLER_147_113 ();
 FILLER_ASAP7_75t_R FILLER_147_129 ();
 DECAPx4_ASAP7_75t_R FILLER_147_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_149 ();
 DECAPx6_ASAP7_75t_R FILLER_147_156 ();
 DECAPx2_ASAP7_75t_R FILLER_147_170 ();
 FILLER_ASAP7_75t_R FILLER_147_182 ();
 DECAPx10_ASAP7_75t_R FILLER_147_187 ();
 DECAPx6_ASAP7_75t_R FILLER_147_209 ();
 DECAPx1_ASAP7_75t_R FILLER_147_223 ();
 DECAPx10_ASAP7_75t_R FILLER_147_230 ();
 DECAPx1_ASAP7_75t_R FILLER_147_252 ();
 DECAPx6_ASAP7_75t_R FILLER_147_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_273 ();
 DECAPx1_ASAP7_75t_R FILLER_147_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_281 ();
 DECAPx10_ASAP7_75t_R FILLER_147_308 ();
 DECAPx6_ASAP7_75t_R FILLER_147_333 ();
 DECAPx1_ASAP7_75t_R FILLER_147_353 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_147_360 ();
 DECAPx1_ASAP7_75t_R FILLER_147_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_393 ();
 FILLER_ASAP7_75t_R FILLER_147_402 ();
 DECAPx6_ASAP7_75t_R FILLER_147_410 ();
 DECAPx2_ASAP7_75t_R FILLER_147_424 ();
 FILLER_ASAP7_75t_R FILLER_147_438 ();
 DECAPx10_ASAP7_75t_R FILLER_147_466 ();
 DECAPx2_ASAP7_75t_R FILLER_147_488 ();
 FILLER_ASAP7_75t_R FILLER_147_520 ();
 DECAPx2_ASAP7_75t_R FILLER_147_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_543 ();
 DECAPx2_ASAP7_75t_R FILLER_147_550 ();
 DECAPx6_ASAP7_75t_R FILLER_147_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_573 ();
 DECAPx2_ASAP7_75t_R FILLER_147_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_586 ();
 DECAPx2_ASAP7_75t_R FILLER_147_593 ();
 FILLER_ASAP7_75t_R FILLER_147_599 ();
 FILLER_ASAP7_75t_R FILLER_147_609 ();
 DECAPx2_ASAP7_75t_R FILLER_147_618 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_147_624 ();
 DECAPx6_ASAP7_75t_R FILLER_147_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_649 ();
 DECAPx4_ASAP7_75t_R FILLER_147_656 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_147_666 ();
 DECAPx2_ASAP7_75t_R FILLER_147_675 ();
 FILLER_ASAP7_75t_R FILLER_147_687 ();
 DECAPx6_ASAP7_75t_R FILLER_147_695 ();
 DECAPx2_ASAP7_75t_R FILLER_147_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_715 ();
 DECAPx4_ASAP7_75t_R FILLER_147_722 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_147_738 ();
 FILLER_ASAP7_75t_R FILLER_147_747 ();
 FILLER_ASAP7_75t_R FILLER_147_755 ();
 DECAPx2_ASAP7_75t_R FILLER_147_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_775 ();
 DECAPx4_ASAP7_75t_R FILLER_147_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_793 ();
 DECAPx4_ASAP7_75t_R FILLER_147_800 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_147_810 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_147_821 ();
 DECAPx4_ASAP7_75t_R FILLER_147_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_838 ();
 FILLER_ASAP7_75t_R FILLER_147_845 ();
 DECAPx2_ASAP7_75t_R FILLER_147_855 ();
 DECAPx4_ASAP7_75t_R FILLER_147_869 ();
 DECAPx10_ASAP7_75t_R FILLER_147_887 ();
 DECAPx4_ASAP7_75t_R FILLER_147_909 ();
 FILLER_ASAP7_75t_R FILLER_147_923 ();
 FILLER_ASAP7_75t_R FILLER_147_927 ();
 FILLER_ASAP7_75t_R FILLER_147_938 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_147_954 ();
 FILLER_ASAP7_75t_R FILLER_147_964 ();
 DECAPx6_ASAP7_75t_R FILLER_147_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_987 ();
 DECAPx2_ASAP7_75t_R FILLER_147_994 ();
 DECAPx6_ASAP7_75t_R FILLER_147_1006 ();
 DECAPx1_ASAP7_75t_R FILLER_147_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_147_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1135 ();
 DECAPx6_ASAP7_75t_R FILLER_147_1157 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1171 ();
 DECAPx4_ASAP7_75t_R FILLER_147_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1240 ();
 DECAPx6_ASAP7_75t_R FILLER_147_1262 ();
 FILLER_ASAP7_75t_R FILLER_147_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_147_1284 ();
 DECAPx6_ASAP7_75t_R FILLER_147_1306 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1320 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1326 ();
 FILLER_ASAP7_75t_R FILLER_147_1337 ();
 FILLER_ASAP7_75t_R FILLER_147_1345 ();
 DECAPx1_ASAP7_75t_R FILLER_147_1353 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_1357 ();
 DECAPx2_ASAP7_75t_R FILLER_147_1368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_147_1374 ();
 DECAPx2_ASAP7_75t_R FILLER_148_2 ();
 FILLER_ASAP7_75t_R FILLER_148_8 ();
 FILLER_ASAP7_75t_R FILLER_148_16 ();
 FILLER_ASAP7_75t_R FILLER_148_24 ();
 DECAPx1_ASAP7_75t_R FILLER_148_29 ();
 DECAPx2_ASAP7_75t_R FILLER_148_36 ();
 FILLER_ASAP7_75t_R FILLER_148_42 ();
 DECAPx10_ASAP7_75t_R FILLER_148_52 ();
 DECAPx2_ASAP7_75t_R FILLER_148_74 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_80 ();
 DECAPx4_ASAP7_75t_R FILLER_148_89 ();
 FILLER_ASAP7_75t_R FILLER_148_99 ();
 DECAPx10_ASAP7_75t_R FILLER_148_107 ();
 FILLER_ASAP7_75t_R FILLER_148_129 ();
 DECAPx2_ASAP7_75t_R FILLER_148_140 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_146 ();
 FILLER_ASAP7_75t_R FILLER_148_155 ();
 FILLER_ASAP7_75t_R FILLER_148_165 ();
 DECAPx2_ASAP7_75t_R FILLER_148_173 ();
 FILLER_ASAP7_75t_R FILLER_148_179 ();
 DECAPx1_ASAP7_75t_R FILLER_148_187 ();
 DECAPx6_ASAP7_75t_R FILLER_148_194 ();
 DECAPx1_ASAP7_75t_R FILLER_148_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_212 ();
 DECAPx10_ASAP7_75t_R FILLER_148_219 ();
 DECAPx2_ASAP7_75t_R FILLER_148_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_247 ();
 DECAPx2_ASAP7_75t_R FILLER_148_254 ();
 FILLER_ASAP7_75t_R FILLER_148_260 ();
 FILLER_ASAP7_75t_R FILLER_148_265 ();
 DECAPx6_ASAP7_75t_R FILLER_148_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_287 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_294 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_300 ();
 FILLER_ASAP7_75t_R FILLER_148_306 ();
 FILLER_ASAP7_75t_R FILLER_148_334 ();
 DECAPx10_ASAP7_75t_R FILLER_148_342 ();
 DECAPx1_ASAP7_75t_R FILLER_148_364 ();
 DECAPx1_ASAP7_75t_R FILLER_148_374 ();
 DECAPx4_ASAP7_75t_R FILLER_148_381 ();
 DECAPx1_ASAP7_75t_R FILLER_148_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_401 ();
 FILLER_ASAP7_75t_R FILLER_148_408 ();
 DECAPx6_ASAP7_75t_R FILLER_148_417 ();
 DECAPx1_ASAP7_75t_R FILLER_148_431 ();
 FILLER_ASAP7_75t_R FILLER_148_441 ();
 FILLER_ASAP7_75t_R FILLER_148_449 ();
 DECAPx1_ASAP7_75t_R FILLER_148_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_461 ();
 FILLER_ASAP7_75t_R FILLER_148_464 ();
 FILLER_ASAP7_75t_R FILLER_148_473 ();
 FILLER_ASAP7_75t_R FILLER_148_481 ();
 DECAPx6_ASAP7_75t_R FILLER_148_490 ();
 FILLER_ASAP7_75t_R FILLER_148_512 ();
 DECAPx10_ASAP7_75t_R FILLER_148_517 ();
 DECAPx10_ASAP7_75t_R FILLER_148_539 ();
 DECAPx2_ASAP7_75t_R FILLER_148_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_567 ();
 DECAPx10_ASAP7_75t_R FILLER_148_574 ();
 DECAPx4_ASAP7_75t_R FILLER_148_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_606 ();
 FILLER_ASAP7_75t_R FILLER_148_613 ();
 FILLER_ASAP7_75t_R FILLER_148_621 ();
 FILLER_ASAP7_75t_R FILLER_148_629 ();
 FILLER_ASAP7_75t_R FILLER_148_639 ();
 FILLER_ASAP7_75t_R FILLER_148_649 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_659 ();
 FILLER_ASAP7_75t_R FILLER_148_668 ();
 FILLER_ASAP7_75t_R FILLER_148_677 ();
 DECAPx2_ASAP7_75t_R FILLER_148_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_691 ();
 FILLER_ASAP7_75t_R FILLER_148_699 ();
 DECAPx2_ASAP7_75t_R FILLER_148_709 ();
 DECAPx2_ASAP7_75t_R FILLER_148_721 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_727 ();
 DECAPx1_ASAP7_75t_R FILLER_148_736 ();
 FILLER_ASAP7_75t_R FILLER_148_748 ();
 DECAPx4_ASAP7_75t_R FILLER_148_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_767 ();
 DECAPx4_ASAP7_75t_R FILLER_148_774 ();
 FILLER_ASAP7_75t_R FILLER_148_791 ();
 DECAPx1_ASAP7_75t_R FILLER_148_801 ();
 DECAPx1_ASAP7_75t_R FILLER_148_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_818 ();
 FILLER_ASAP7_75t_R FILLER_148_828 ();
 FILLER_ASAP7_75t_R FILLER_148_836 ();
 FILLER_ASAP7_75t_R FILLER_148_848 ();
 FILLER_ASAP7_75t_R FILLER_148_857 ();
 FILLER_ASAP7_75t_R FILLER_148_865 ();
 DECAPx2_ASAP7_75t_R FILLER_148_873 ();
 FILLER_ASAP7_75t_R FILLER_148_879 ();
 FILLER_ASAP7_75t_R FILLER_148_890 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_901 ();
 DECAPx2_ASAP7_75t_R FILLER_148_912 ();
 FILLER_ASAP7_75t_R FILLER_148_918 ();
 DECAPx6_ASAP7_75t_R FILLER_148_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_940 ();
 FILLER_ASAP7_75t_R FILLER_148_952 ();
 FILLER_ASAP7_75t_R FILLER_148_963 ();
 FILLER_ASAP7_75t_R FILLER_148_973 ();
 FILLER_ASAP7_75t_R FILLER_148_982 ();
 DECAPx6_ASAP7_75t_R FILLER_148_987 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1009 ();
 DECAPx6_ASAP7_75t_R FILLER_148_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1051 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_1057 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1089 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_1095 ();
 FILLER_ASAP7_75t_R FILLER_148_1101 ();
 DECAPx6_ASAP7_75t_R FILLER_148_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1120 ();
 FILLER_ASAP7_75t_R FILLER_148_1124 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1135 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1145 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_1165 ();
 FILLER_ASAP7_75t_R FILLER_148_1171 ();
 FILLER_ASAP7_75t_R FILLER_148_1182 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1208 ();
 FILLER_ASAP7_75t_R FILLER_148_1223 ();
 DECAPx4_ASAP7_75t_R FILLER_148_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1252 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_1258 ();
 FILLER_ASAP7_75t_R FILLER_148_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_148_1276 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1298 ();
 FILLER_ASAP7_75t_R FILLER_148_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_148_1318 ();
 DECAPx2_ASAP7_75t_R FILLER_148_1340 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_1346 ();
 FILLER_ASAP7_75t_R FILLER_148_1375 ();
 DECAPx1_ASAP7_75t_R FILLER_149_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_6 ();
 DECAPx2_ASAP7_75t_R FILLER_149_13 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_149_19 ();
 DECAPx1_ASAP7_75t_R FILLER_149_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_32 ();
 FILLER_ASAP7_75t_R FILLER_149_39 ();
 DECAPx6_ASAP7_75t_R FILLER_149_49 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_149_63 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_149_72 ();
 DECAPx6_ASAP7_75t_R FILLER_149_101 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_149_115 ();
 DECAPx1_ASAP7_75t_R FILLER_149_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_129 ();
 FILLER_ASAP7_75t_R FILLER_149_136 ();
 DECAPx4_ASAP7_75t_R FILLER_149_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_174 ();
 FILLER_ASAP7_75t_R FILLER_149_201 ();
 FILLER_ASAP7_75t_R FILLER_149_229 ();
 FILLER_ASAP7_75t_R FILLER_149_237 ();
 DECAPx2_ASAP7_75t_R FILLER_149_242 ();
 FILLER_ASAP7_75t_R FILLER_149_248 ();
 FILLER_ASAP7_75t_R FILLER_149_256 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_149_264 ();
 FILLER_ASAP7_75t_R FILLER_149_275 ();
 DECAPx2_ASAP7_75t_R FILLER_149_283 ();
 DECAPx6_ASAP7_75t_R FILLER_149_295 ();
 DECAPx1_ASAP7_75t_R FILLER_149_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_313 ();
 DECAPx4_ASAP7_75t_R FILLER_149_320 ();
 FILLER_ASAP7_75t_R FILLER_149_356 ();
 FILLER_ASAP7_75t_R FILLER_149_361 ();
 DECAPx10_ASAP7_75t_R FILLER_149_369 ();
 DECAPx6_ASAP7_75t_R FILLER_149_391 ();
 DECAPx1_ASAP7_75t_R FILLER_149_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_409 ();
 FILLER_ASAP7_75t_R FILLER_149_426 ();
 DECAPx6_ASAP7_75t_R FILLER_149_434 ();
 DECAPx2_ASAP7_75t_R FILLER_149_448 ();
 FILLER_ASAP7_75t_R FILLER_149_480 ();
 DECAPx4_ASAP7_75t_R FILLER_149_508 ();
 DECAPx4_ASAP7_75t_R FILLER_149_526 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_149_536 ();
 DECAPx1_ASAP7_75t_R FILLER_149_545 ();
 DECAPx1_ASAP7_75t_R FILLER_149_552 ();
 DECAPx10_ASAP7_75t_R FILLER_149_582 ();
 DECAPx10_ASAP7_75t_R FILLER_149_604 ();
 DECAPx1_ASAP7_75t_R FILLER_149_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_630 ();
 DECAPx10_ASAP7_75t_R FILLER_149_637 ();
 DECAPx2_ASAP7_75t_R FILLER_149_659 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_149_665 ();
 DECAPx4_ASAP7_75t_R FILLER_149_676 ();
 FILLER_ASAP7_75t_R FILLER_149_692 ();
 DECAPx2_ASAP7_75t_R FILLER_149_700 ();
 FILLER_ASAP7_75t_R FILLER_149_706 ();
 DECAPx2_ASAP7_75t_R FILLER_149_714 ();
 DECAPx4_ASAP7_75t_R FILLER_149_726 ();
 FILLER_ASAP7_75t_R FILLER_149_736 ();
 DECAPx10_ASAP7_75t_R FILLER_149_744 ();
 DECAPx10_ASAP7_75t_R FILLER_149_766 ();
 DECAPx1_ASAP7_75t_R FILLER_149_788 ();
 FILLER_ASAP7_75t_R FILLER_149_804 ();
 FILLER_ASAP7_75t_R FILLER_149_809 ();
 FILLER_ASAP7_75t_R FILLER_149_817 ();
 DECAPx10_ASAP7_75t_R FILLER_149_825 ();
 DECAPx10_ASAP7_75t_R FILLER_149_847 ();
 DECAPx1_ASAP7_75t_R FILLER_149_869 ();
 FILLER_ASAP7_75t_R FILLER_149_879 ();
 DECAPx4_ASAP7_75t_R FILLER_149_891 ();
 DECAPx6_ASAP7_75t_R FILLER_149_909 ();
 FILLER_ASAP7_75t_R FILLER_149_923 ();
 DECAPx10_ASAP7_75t_R FILLER_149_927 ();
 DECAPx4_ASAP7_75t_R FILLER_149_949 ();
 DECAPx10_ASAP7_75t_R FILLER_149_966 ();
 DECAPx10_ASAP7_75t_R FILLER_149_988 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1016 ();
 FILLER_ASAP7_75t_R FILLER_149_1020 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1033 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_149_1056 ();
 FILLER_ASAP7_75t_R FILLER_149_1065 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1070 ();
 DECAPx1_ASAP7_75t_R FILLER_149_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_1114 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1124 ();
 FILLER_ASAP7_75t_R FILLER_149_1136 ();
 FILLER_ASAP7_75t_R FILLER_149_1164 ();
 DECAPx1_ASAP7_75t_R FILLER_149_1176 ();
 FILLER_ASAP7_75t_R FILLER_149_1206 ();
 FILLER_ASAP7_75t_R FILLER_149_1217 ();
 FILLER_ASAP7_75t_R FILLER_149_1222 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1250 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_149_1256 ();
 FILLER_ASAP7_75t_R FILLER_149_1285 ();
 FILLER_ASAP7_75t_R FILLER_149_1295 ();
 DECAPx1_ASAP7_75t_R FILLER_149_1303 ();
 FILLER_ASAP7_75t_R FILLER_149_1310 ();
 DECAPx4_ASAP7_75t_R FILLER_149_1321 ();
 FILLER_ASAP7_75t_R FILLER_149_1331 ();
 DECAPx6_ASAP7_75t_R FILLER_149_1343 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_149_1363 ();
 DECAPx2_ASAP7_75t_R FILLER_149_1369 ();
 FILLER_ASAP7_75t_R FILLER_149_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_150_2 ();
 DECAPx1_ASAP7_75t_R FILLER_150_34 ();
 DECAPx1_ASAP7_75t_R FILLER_150_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_48 ();
 DECAPx1_ASAP7_75t_R FILLER_150_55 ();
 DECAPx6_ASAP7_75t_R FILLER_150_65 ();
 DECAPx1_ASAP7_75t_R FILLER_150_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_89 ();
 DECAPx6_ASAP7_75t_R FILLER_150_93 ();
 FILLER_ASAP7_75t_R FILLER_150_107 ();
 DECAPx1_ASAP7_75t_R FILLER_150_115 ();
 FILLER_ASAP7_75t_R FILLER_150_127 ();
 DECAPx4_ASAP7_75t_R FILLER_150_135 ();
 FILLER_ASAP7_75t_R FILLER_150_151 ();
 DECAPx10_ASAP7_75t_R FILLER_150_156 ();
 DECAPx2_ASAP7_75t_R FILLER_150_184 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_150_190 ();
 DECAPx2_ASAP7_75t_R FILLER_150_199 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_150_205 ();
 DECAPx1_ASAP7_75t_R FILLER_150_214 ();
 FILLER_ASAP7_75t_R FILLER_150_221 ();
 FILLER_ASAP7_75t_R FILLER_150_229 ();
 FILLER_ASAP7_75t_R FILLER_150_240 ();
 FILLER_ASAP7_75t_R FILLER_150_250 ();
 FILLER_ASAP7_75t_R FILLER_150_274 ();
 DECAPx4_ASAP7_75t_R FILLER_150_302 ();
 DECAPx1_ASAP7_75t_R FILLER_150_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_322 ();
 DECAPx4_ASAP7_75t_R FILLER_150_326 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_150_336 ();
 DECAPx2_ASAP7_75t_R FILLER_150_345 ();
 FILLER_ASAP7_75t_R FILLER_150_365 ();
 DECAPx2_ASAP7_75t_R FILLER_150_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_381 ();
 FILLER_ASAP7_75t_R FILLER_150_388 ();
 DECAPx1_ASAP7_75t_R FILLER_150_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_397 ();
 DECAPx4_ASAP7_75t_R FILLER_150_404 ();
 FILLER_ASAP7_75t_R FILLER_150_414 ();
 FILLER_ASAP7_75t_R FILLER_150_422 ();
 DECAPx2_ASAP7_75t_R FILLER_150_432 ();
 DECAPx4_ASAP7_75t_R FILLER_150_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_454 ();
 DECAPx1_ASAP7_75t_R FILLER_150_458 ();
 DECAPx2_ASAP7_75t_R FILLER_150_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_470 ();
 DECAPx4_ASAP7_75t_R FILLER_150_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_484 ();
 DECAPx2_ASAP7_75t_R FILLER_150_491 ();
 DECAPx4_ASAP7_75t_R FILLER_150_500 ();
 FILLER_ASAP7_75t_R FILLER_150_516 ();
 DECAPx2_ASAP7_75t_R FILLER_150_526 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_150_532 ();
 FILLER_ASAP7_75t_R FILLER_150_561 ();
 FILLER_ASAP7_75t_R FILLER_150_569 ();
 FILLER_ASAP7_75t_R FILLER_150_574 ();
 DECAPx2_ASAP7_75t_R FILLER_150_579 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_150_585 ();
 FILLER_ASAP7_75t_R FILLER_150_595 ();
 DECAPx4_ASAP7_75t_R FILLER_150_603 ();
 DECAPx10_ASAP7_75t_R FILLER_150_623 ();
 DECAPx4_ASAP7_75t_R FILLER_150_653 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_150_663 ();
 DECAPx6_ASAP7_75t_R FILLER_150_673 ();
 DECAPx2_ASAP7_75t_R FILLER_150_698 ();
 FILLER_ASAP7_75t_R FILLER_150_704 ();
 DECAPx1_ASAP7_75t_R FILLER_150_713 ();
 DECAPx10_ASAP7_75t_R FILLER_150_723 ();
 DECAPx1_ASAP7_75t_R FILLER_150_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_749 ();
 DECAPx4_ASAP7_75t_R FILLER_150_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_770 ();
 FILLER_ASAP7_75t_R FILLER_150_781 ();
 DECAPx10_ASAP7_75t_R FILLER_150_790 ();
 DECAPx10_ASAP7_75t_R FILLER_150_815 ();
 DECAPx6_ASAP7_75t_R FILLER_150_847 ();
 DECAPx10_ASAP7_75t_R FILLER_150_867 ();
 DECAPx10_ASAP7_75t_R FILLER_150_889 ();
 DECAPx1_ASAP7_75t_R FILLER_150_911 ();
 DECAPx10_ASAP7_75t_R FILLER_150_921 ();
 DECAPx10_ASAP7_75t_R FILLER_150_949 ();
 DECAPx4_ASAP7_75t_R FILLER_150_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_981 ();
 FILLER_ASAP7_75t_R FILLER_150_991 ();
 DECAPx1_ASAP7_75t_R FILLER_150_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1003 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_150_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_150_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1053 ();
 FILLER_ASAP7_75t_R FILLER_150_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_150_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1077 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1092 ();
 FILLER_ASAP7_75t_R FILLER_150_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1107 ();
 FILLER_ASAP7_75t_R FILLER_150_1113 ();
 FILLER_ASAP7_75t_R FILLER_150_1118 ();
 FILLER_ASAP7_75t_R FILLER_150_1129 ();
 FILLER_ASAP7_75t_R FILLER_150_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1147 ();
 DECAPx6_ASAP7_75t_R FILLER_150_1156 ();
 DECAPx1_ASAP7_75t_R FILLER_150_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1174 ();
 DECAPx6_ASAP7_75t_R FILLER_150_1185 ();
 FILLER_ASAP7_75t_R FILLER_150_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1207 ();
 FILLER_ASAP7_75t_R FILLER_150_1213 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1218 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_150_1241 ();
 DECAPx1_ASAP7_75t_R FILLER_150_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1267 ();
 DECAPx6_ASAP7_75t_R FILLER_150_1276 ();
 FILLER_ASAP7_75t_R FILLER_150_1290 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1295 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_150_1301 ();
 FILLER_ASAP7_75t_R FILLER_150_1310 ();
 FILLER_ASAP7_75t_R FILLER_150_1315 ();
 FILLER_ASAP7_75t_R FILLER_150_1343 ();
 DECAPx10_ASAP7_75t_R FILLER_150_1348 ();
 DECAPx2_ASAP7_75t_R FILLER_150_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_1376 ();
 FILLER_ASAP7_75t_R FILLER_151_2 ();
 DECAPx2_ASAP7_75t_R FILLER_151_10 ();
 FILLER_ASAP7_75t_R FILLER_151_22 ();
 FILLER_ASAP7_75t_R FILLER_151_30 ();
 DECAPx10_ASAP7_75t_R FILLER_151_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_57 ();
 FILLER_ASAP7_75t_R FILLER_151_68 ();
 FILLER_ASAP7_75t_R FILLER_151_76 ();
 DECAPx6_ASAP7_75t_R FILLER_151_84 ();
 DECAPx1_ASAP7_75t_R FILLER_151_98 ();
 FILLER_ASAP7_75t_R FILLER_151_110 ();
 FILLER_ASAP7_75t_R FILLER_151_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_143 ();
 DECAPx6_ASAP7_75t_R FILLER_151_172 ();
 DECAPx1_ASAP7_75t_R FILLER_151_186 ();
 DECAPx4_ASAP7_75t_R FILLER_151_216 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_226 ();
 DECAPx6_ASAP7_75t_R FILLER_151_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_249 ();
 DECAPx2_ASAP7_75t_R FILLER_151_276 ();
 FILLER_ASAP7_75t_R FILLER_151_282 ();
 FILLER_ASAP7_75t_R FILLER_151_290 ();
 DECAPx4_ASAP7_75t_R FILLER_151_295 ();
 FILLER_ASAP7_75t_R FILLER_151_313 ();
 DECAPx10_ASAP7_75t_R FILLER_151_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_343 ();
 DECAPx1_ASAP7_75t_R FILLER_151_347 ();
 DECAPx6_ASAP7_75t_R FILLER_151_357 ();
 DECAPx1_ASAP7_75t_R FILLER_151_371 ();
 FILLER_ASAP7_75t_R FILLER_151_401 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_411 ();
 FILLER_ASAP7_75t_R FILLER_151_436 ();
 FILLER_ASAP7_75t_R FILLER_151_446 ();
 DECAPx6_ASAP7_75t_R FILLER_151_454 ();
 DECAPx1_ASAP7_75t_R FILLER_151_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_472 ();
 DECAPx10_ASAP7_75t_R FILLER_151_495 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_517 ();
 DECAPx4_ASAP7_75t_R FILLER_151_526 ();
 FILLER_ASAP7_75t_R FILLER_151_536 ();
 DECAPx6_ASAP7_75t_R FILLER_151_544 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_558 ();
 DECAPx6_ASAP7_75t_R FILLER_151_567 ();
 DECAPx1_ASAP7_75t_R FILLER_151_581 ();
 DECAPx1_ASAP7_75t_R FILLER_151_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_598 ();
 FILLER_ASAP7_75t_R FILLER_151_606 ();
 DECAPx6_ASAP7_75t_R FILLER_151_616 ();
 DECAPx2_ASAP7_75t_R FILLER_151_636 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_642 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_652 ();
 DECAPx2_ASAP7_75t_R FILLER_151_661 ();
 DECAPx6_ASAP7_75t_R FILLER_151_673 ();
 DECAPx10_ASAP7_75t_R FILLER_151_693 ();
 FILLER_ASAP7_75t_R FILLER_151_721 ();
 DECAPx6_ASAP7_75t_R FILLER_151_729 ();
 FILLER_ASAP7_75t_R FILLER_151_749 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_757 ();
 FILLER_ASAP7_75t_R FILLER_151_763 ();
 FILLER_ASAP7_75t_R FILLER_151_774 ();
 DECAPx4_ASAP7_75t_R FILLER_151_782 ();
 FILLER_ASAP7_75t_R FILLER_151_792 ();
 DECAPx6_ASAP7_75t_R FILLER_151_803 ();
 FILLER_ASAP7_75t_R FILLER_151_817 ();
 DECAPx2_ASAP7_75t_R FILLER_151_824 ();
 FILLER_ASAP7_75t_R FILLER_151_830 ();
 DECAPx4_ASAP7_75t_R FILLER_151_846 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_856 ();
 FILLER_ASAP7_75t_R FILLER_151_868 ();
 FILLER_ASAP7_75t_R FILLER_151_878 ();
 DECAPx1_ASAP7_75t_R FILLER_151_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_890 ();
 DECAPx1_ASAP7_75t_R FILLER_151_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_903 ();
 FILLER_ASAP7_75t_R FILLER_151_907 ();
 DECAPx2_ASAP7_75t_R FILLER_151_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_924 ();
 DECAPx6_ASAP7_75t_R FILLER_151_927 ();
 FILLER_ASAP7_75t_R FILLER_151_941 ();
 DECAPx2_ASAP7_75t_R FILLER_151_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_958 ();
 DECAPx4_ASAP7_75t_R FILLER_151_966 ();
 FILLER_ASAP7_75t_R FILLER_151_976 ();
 FILLER_ASAP7_75t_R FILLER_151_981 ();
 FILLER_ASAP7_75t_R FILLER_151_992 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1002 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_1012 ();
 FILLER_ASAP7_75t_R FILLER_151_1022 ();
 FILLER_ASAP7_75t_R FILLER_151_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_151_1038 ();
 FILLER_ASAP7_75t_R FILLER_151_1060 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1068 ();
 FILLER_ASAP7_75t_R FILLER_151_1078 ();
 FILLER_ASAP7_75t_R FILLER_151_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_151_1094 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_151_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_151_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_151_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_151_1179 ();
 DECAPx6_ASAP7_75t_R FILLER_151_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_151_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1221 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1228 ();
 FILLER_ASAP7_75t_R FILLER_151_1238 ();
 FILLER_ASAP7_75t_R FILLER_151_1266 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_1288 ();
 FILLER_ASAP7_75t_R FILLER_151_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_151_1303 ();
 DECAPx1_ASAP7_75t_R FILLER_151_1325 ();
 DECAPx4_ASAP7_75t_R FILLER_151_1339 ();
 FILLER_ASAP7_75t_R FILLER_151_1375 ();
 FILLER_ASAP7_75t_R FILLER_152_2 ();
 FILLER_ASAP7_75t_R FILLER_152_10 ();
 FILLER_ASAP7_75t_R FILLER_152_18 ();
 DECAPx6_ASAP7_75t_R FILLER_152_25 ();
 DECAPx1_ASAP7_75t_R FILLER_152_39 ();
 DECAPx6_ASAP7_75t_R FILLER_152_51 ();
 FILLER_ASAP7_75t_R FILLER_152_91 ();
 DECAPx1_ASAP7_75t_R FILLER_152_96 ();
 FILLER_ASAP7_75t_R FILLER_152_107 ();
 DECAPx2_ASAP7_75t_R FILLER_152_115 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_121 ();
 DECAPx4_ASAP7_75t_R FILLER_152_132 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_142 ();
 FILLER_ASAP7_75t_R FILLER_152_151 ();
 FILLER_ASAP7_75t_R FILLER_152_159 ();
 DECAPx1_ASAP7_75t_R FILLER_152_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_168 ();
 FILLER_ASAP7_75t_R FILLER_152_175 ();
 DECAPx6_ASAP7_75t_R FILLER_152_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_197 ();
 FILLER_ASAP7_75t_R FILLER_152_204 ();
 DECAPx10_ASAP7_75t_R FILLER_152_209 ();
 DECAPx6_ASAP7_75t_R FILLER_152_231 ();
 DECAPx2_ASAP7_75t_R FILLER_152_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_251 ();
 DECAPx2_ASAP7_75t_R FILLER_152_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_264 ();
 DECAPx10_ASAP7_75t_R FILLER_152_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_290 ();
 DECAPx6_ASAP7_75t_R FILLER_152_294 ();
 FILLER_ASAP7_75t_R FILLER_152_316 ();
 DECAPx4_ASAP7_75t_R FILLER_152_324 ();
 DECAPx4_ASAP7_75t_R FILLER_152_340 ();
 DECAPx2_ASAP7_75t_R FILLER_152_356 ();
 DECAPx2_ASAP7_75t_R FILLER_152_370 ();
 FILLER_ASAP7_75t_R FILLER_152_376 ();
 DECAPx4_ASAP7_75t_R FILLER_152_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_394 ();
 FILLER_ASAP7_75t_R FILLER_152_401 ();
 DECAPx1_ASAP7_75t_R FILLER_152_411 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_421 ();
 DECAPx2_ASAP7_75t_R FILLER_152_433 ();
 FILLER_ASAP7_75t_R FILLER_152_439 ();
 DECAPx6_ASAP7_75t_R FILLER_152_444 ();
 DECAPx1_ASAP7_75t_R FILLER_152_458 ();
 FILLER_ASAP7_75t_R FILLER_152_464 ();
 DECAPx1_ASAP7_75t_R FILLER_152_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_476 ();
 DECAPx2_ASAP7_75t_R FILLER_152_503 ();
 FILLER_ASAP7_75t_R FILLER_152_509 ();
 FILLER_ASAP7_75t_R FILLER_152_517 ();
 DECAPx6_ASAP7_75t_R FILLER_152_522 ();
 DECAPx2_ASAP7_75t_R FILLER_152_536 ();
 DECAPx2_ASAP7_75t_R FILLER_152_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_554 ();
 DECAPx2_ASAP7_75t_R FILLER_152_581 ();
 FILLER_ASAP7_75t_R FILLER_152_587 ();
 FILLER_ASAP7_75t_R FILLER_152_595 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_603 ();
 FILLER_ASAP7_75t_R FILLER_152_615 ();
 DECAPx2_ASAP7_75t_R FILLER_152_625 ();
 FILLER_ASAP7_75t_R FILLER_152_637 ();
 DECAPx2_ASAP7_75t_R FILLER_152_645 ();
 FILLER_ASAP7_75t_R FILLER_152_651 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_667 ();
 DECAPx1_ASAP7_75t_R FILLER_152_676 ();
 FILLER_ASAP7_75t_R FILLER_152_686 ();
 FILLER_ASAP7_75t_R FILLER_152_695 ();
 DECAPx10_ASAP7_75t_R FILLER_152_707 ();
 DECAPx1_ASAP7_75t_R FILLER_152_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_742 ();
 DECAPx6_ASAP7_75t_R FILLER_152_749 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_763 ();
 DECAPx2_ASAP7_75t_R FILLER_152_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_780 ();
 FILLER_ASAP7_75t_R FILLER_152_789 ();
 DECAPx4_ASAP7_75t_R FILLER_152_800 ();
 FILLER_ASAP7_75t_R FILLER_152_819 ();
 DECAPx2_ASAP7_75t_R FILLER_152_828 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_834 ();
 FILLER_ASAP7_75t_R FILLER_152_845 ();
 FILLER_ASAP7_75t_R FILLER_152_853 ();
 FILLER_ASAP7_75t_R FILLER_152_858 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_863 ();
 DECAPx1_ASAP7_75t_R FILLER_152_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_879 ();
 DECAPx1_ASAP7_75t_R FILLER_152_887 ();
 FILLER_ASAP7_75t_R FILLER_152_897 ();
 FILLER_ASAP7_75t_R FILLER_152_906 ();
 FILLER_ASAP7_75t_R FILLER_152_916 ();
 FILLER_ASAP7_75t_R FILLER_152_927 ();
 FILLER_ASAP7_75t_R FILLER_152_932 ();
 FILLER_ASAP7_75t_R FILLER_152_942 ();
 DECAPx4_ASAP7_75t_R FILLER_152_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_962 ();
 DECAPx1_ASAP7_75t_R FILLER_152_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_973 ();
 DECAPx1_ASAP7_75t_R FILLER_152_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_985 ();
 FILLER_ASAP7_75t_R FILLER_152_992 ();
 DECAPx6_ASAP7_75t_R FILLER_152_997 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1011 ();
 FILLER_ASAP7_75t_R FILLER_152_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_152_1030 ();
 FILLER_ASAP7_75t_R FILLER_152_1036 ();
 FILLER_ASAP7_75t_R FILLER_152_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1058 ();
 DECAPx4_ASAP7_75t_R FILLER_152_1080 ();
 FILLER_ASAP7_75t_R FILLER_152_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_152_1100 ();
 DECAPx4_ASAP7_75t_R FILLER_152_1109 ();
 FILLER_ASAP7_75t_R FILLER_152_1119 ();
 DECAPx4_ASAP7_75t_R FILLER_152_1127 ();
 FILLER_ASAP7_75t_R FILLER_152_1137 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1145 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1165 ();
 FILLER_ASAP7_75t_R FILLER_152_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1208 ();
 DECAPx4_ASAP7_75t_R FILLER_152_1230 ();
 FILLER_ASAP7_75t_R FILLER_152_1250 ();
 FILLER_ASAP7_75t_R FILLER_152_1260 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1269 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_1276 ();
 DECAPx4_ASAP7_75t_R FILLER_152_1288 ();
 FILLER_ASAP7_75t_R FILLER_152_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_152_1314 ();
 DECAPx6_ASAP7_75t_R FILLER_152_1336 ();
 DECAPx2_ASAP7_75t_R FILLER_152_1353 ();
 FILLER_ASAP7_75t_R FILLER_152_1367 ();
 DECAPx1_ASAP7_75t_R FILLER_152_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_1376 ();
 FILLER_ASAP7_75t_R FILLER_153_2 ();
 DECAPx1_ASAP7_75t_R FILLER_153_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_34 ();
 FILLER_ASAP7_75t_R FILLER_153_38 ();
 FILLER_ASAP7_75t_R FILLER_153_46 ();
 DECAPx10_ASAP7_75t_R FILLER_153_54 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_76 ();
 DECAPx6_ASAP7_75t_R FILLER_153_82 ();
 FILLER_ASAP7_75t_R FILLER_153_96 ();
 DECAPx4_ASAP7_75t_R FILLER_153_104 ();
 FILLER_ASAP7_75t_R FILLER_153_114 ();
 FILLER_ASAP7_75t_R FILLER_153_122 ();
 DECAPx1_ASAP7_75t_R FILLER_153_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_134 ();
 FILLER_ASAP7_75t_R FILLER_153_138 ();
 DECAPx10_ASAP7_75t_R FILLER_153_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_168 ();
 FILLER_ASAP7_75t_R FILLER_153_195 ();
 FILLER_ASAP7_75t_R FILLER_153_200 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_208 ();
 FILLER_ASAP7_75t_R FILLER_153_218 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_226 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_239 ();
 FILLER_ASAP7_75t_R FILLER_153_248 ();
 DECAPx10_ASAP7_75t_R FILLER_153_253 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_275 ();
 DECAPx1_ASAP7_75t_R FILLER_153_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_288 ();
 FILLER_ASAP7_75t_R FILLER_153_295 ();
 DECAPx10_ASAP7_75t_R FILLER_153_303 ();
 DECAPx2_ASAP7_75t_R FILLER_153_325 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_331 ();
 FILLER_ASAP7_75t_R FILLER_153_340 ();
 DECAPx1_ASAP7_75t_R FILLER_153_348 ();
 FILLER_ASAP7_75t_R FILLER_153_374 ();
 DECAPx1_ASAP7_75t_R FILLER_153_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_386 ();
 DECAPx1_ASAP7_75t_R FILLER_153_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_397 ();
 DECAPx1_ASAP7_75t_R FILLER_153_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_405 ();
 DECAPx4_ASAP7_75t_R FILLER_153_428 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_438 ();
 DECAPx2_ASAP7_75t_R FILLER_153_447 ();
 FILLER_ASAP7_75t_R FILLER_153_479 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_484 ();
 FILLER_ASAP7_75t_R FILLER_153_493 ();
 DECAPx1_ASAP7_75t_R FILLER_153_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_502 ();
 FILLER_ASAP7_75t_R FILLER_153_529 ();
 DECAPx2_ASAP7_75t_R FILLER_153_557 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_563 ();
 FILLER_ASAP7_75t_R FILLER_153_572 ();
 DECAPx4_ASAP7_75t_R FILLER_153_577 ();
 FILLER_ASAP7_75t_R FILLER_153_587 ();
 DECAPx4_ASAP7_75t_R FILLER_153_595 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_605 ();
 FILLER_ASAP7_75t_R FILLER_153_614 ();
 DECAPx4_ASAP7_75t_R FILLER_153_622 ();
 DECAPx2_ASAP7_75t_R FILLER_153_639 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_645 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_656 ();
 DECAPx6_ASAP7_75t_R FILLER_153_667 ();
 DECAPx2_ASAP7_75t_R FILLER_153_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_687 ();
 DECAPx10_ASAP7_75t_R FILLER_153_700 ();
 DECAPx2_ASAP7_75t_R FILLER_153_722 ();
 DECAPx4_ASAP7_75t_R FILLER_153_737 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_747 ();
 DECAPx1_ASAP7_75t_R FILLER_153_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_760 ();
 FILLER_ASAP7_75t_R FILLER_153_764 ();
 DECAPx2_ASAP7_75t_R FILLER_153_772 ();
 DECAPx6_ASAP7_75t_R FILLER_153_782 ();
 FILLER_ASAP7_75t_R FILLER_153_796 ();
 FILLER_ASAP7_75t_R FILLER_153_804 ();
 DECAPx2_ASAP7_75t_R FILLER_153_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_818 ();
 FILLER_ASAP7_75t_R FILLER_153_829 ();
 DECAPx10_ASAP7_75t_R FILLER_153_837 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_859 ();
 DECAPx10_ASAP7_75t_R FILLER_153_865 ();
 DECAPx6_ASAP7_75t_R FILLER_153_887 ();
 DECAPx2_ASAP7_75t_R FILLER_153_908 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_914 ();
 FILLER_ASAP7_75t_R FILLER_153_923 ();
 FILLER_ASAP7_75t_R FILLER_153_927 ();
 FILLER_ASAP7_75t_R FILLER_153_939 ();
 DECAPx1_ASAP7_75t_R FILLER_153_948 ();
 FILLER_ASAP7_75t_R FILLER_153_959 ();
 FILLER_ASAP7_75t_R FILLER_153_970 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_978 ();
 DECAPx4_ASAP7_75t_R FILLER_153_990 ();
 DECAPx6_ASAP7_75t_R FILLER_153_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1022 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_1030 ();
 FILLER_ASAP7_75t_R FILLER_153_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1071 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_1081 ();
 FILLER_ASAP7_75t_R FILLER_153_1090 ();
 FILLER_ASAP7_75t_R FILLER_153_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1133 ();
 FILLER_ASAP7_75t_R FILLER_153_1144 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1172 ();
 FILLER_ASAP7_75t_R FILLER_153_1178 ();
 FILLER_ASAP7_75t_R FILLER_153_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1221 ();
 FILLER_ASAP7_75t_R FILLER_153_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1238 ();
 FILLER_ASAP7_75t_R FILLER_153_1245 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_1253 ();
 FILLER_ASAP7_75t_R FILLER_153_1266 ();
 DECAPx2_ASAP7_75t_R FILLER_153_1274 ();
 FILLER_ASAP7_75t_R FILLER_153_1280 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1296 ();
 FILLER_ASAP7_75t_R FILLER_153_1305 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1333 ();
 FILLER_ASAP7_75t_R FILLER_153_1346 ();
 DECAPx1_ASAP7_75t_R FILLER_153_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_1358 ();
 FILLER_ASAP7_75t_R FILLER_153_1367 ();
 FILLER_ASAP7_75t_R FILLER_153_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_154_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_8 ();
 FILLER_ASAP7_75t_R FILLER_154_15 ();
 DECAPx4_ASAP7_75t_R FILLER_154_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_30 ();
 FILLER_ASAP7_75t_R FILLER_154_37 ();
 DECAPx6_ASAP7_75t_R FILLER_154_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_59 ();
 DECAPx10_ASAP7_75t_R FILLER_154_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_88 ();
 DECAPx4_ASAP7_75t_R FILLER_154_95 ();
 FILLER_ASAP7_75t_R FILLER_154_131 ();
 DECAPx4_ASAP7_75t_R FILLER_154_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_169 ();
 DECAPx2_ASAP7_75t_R FILLER_154_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_182 ();
 DECAPx6_ASAP7_75t_R FILLER_154_186 ();
 DECAPx1_ASAP7_75t_R FILLER_154_200 ();
 DECAPx2_ASAP7_75t_R FILLER_154_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_218 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_154_231 ();
 DECAPx2_ASAP7_75t_R FILLER_154_260 ();
 FILLER_ASAP7_75t_R FILLER_154_266 ();
 FILLER_ASAP7_75t_R FILLER_154_294 ();
 DECAPx2_ASAP7_75t_R FILLER_154_302 ();
 DECAPx1_ASAP7_75t_R FILLER_154_316 ();
 FILLER_ASAP7_75t_R FILLER_154_328 ();
 FILLER_ASAP7_75t_R FILLER_154_337 ();
 DECAPx2_ASAP7_75t_R FILLER_154_345 ();
 DECAPx1_ASAP7_75t_R FILLER_154_354 ();
 FILLER_ASAP7_75t_R FILLER_154_364 ();
 DECAPx2_ASAP7_75t_R FILLER_154_369 ();
 DECAPx1_ASAP7_75t_R FILLER_154_401 ();
 FILLER_ASAP7_75t_R FILLER_154_413 ();
 DECAPx2_ASAP7_75t_R FILLER_154_421 ();
 DECAPx2_ASAP7_75t_R FILLER_154_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_154_459 ();
 FILLER_ASAP7_75t_R FILLER_154_464 ();
 DECAPx1_ASAP7_75t_R FILLER_154_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_476 ();
 FILLER_ASAP7_75t_R FILLER_154_480 ();
 DECAPx6_ASAP7_75t_R FILLER_154_488 ();
 DECAPx1_ASAP7_75t_R FILLER_154_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_506 ();
 DECAPx1_ASAP7_75t_R FILLER_154_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_517 ();
 DECAPx6_ASAP7_75t_R FILLER_154_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_535 ();
 DECAPx1_ASAP7_75t_R FILLER_154_542 ();
 DECAPx6_ASAP7_75t_R FILLER_154_549 ();
 DECAPx2_ASAP7_75t_R FILLER_154_563 ();
 DECAPx6_ASAP7_75t_R FILLER_154_575 ();
 FILLER_ASAP7_75t_R FILLER_154_589 ();
 DECAPx10_ASAP7_75t_R FILLER_154_598 ();
 DECAPx4_ASAP7_75t_R FILLER_154_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_630 ();
 FILLER_ASAP7_75t_R FILLER_154_637 ();
 FILLER_ASAP7_75t_R FILLER_154_651 ();
 DECAPx6_ASAP7_75t_R FILLER_154_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_673 ();
 FILLER_ASAP7_75t_R FILLER_154_684 ();
 DECAPx4_ASAP7_75t_R FILLER_154_698 ();
 DECAPx1_ASAP7_75t_R FILLER_154_714 ();
 DECAPx2_ASAP7_75t_R FILLER_154_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_730 ();
 DECAPx4_ASAP7_75t_R FILLER_154_737 ();
 FILLER_ASAP7_75t_R FILLER_154_747 ();
 DECAPx2_ASAP7_75t_R FILLER_154_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_762 ();
 DECAPx10_ASAP7_75t_R FILLER_154_772 ();
 DECAPx10_ASAP7_75t_R FILLER_154_794 ();
 DECAPx10_ASAP7_75t_R FILLER_154_816 ();
 FILLER_ASAP7_75t_R FILLER_154_838 ();
 FILLER_ASAP7_75t_R FILLER_154_849 ();
 DECAPx6_ASAP7_75t_R FILLER_154_858 ();
 FILLER_ASAP7_75t_R FILLER_154_872 ();
 FILLER_ASAP7_75t_R FILLER_154_880 ();
 DECAPx10_ASAP7_75t_R FILLER_154_888 ();
 DECAPx1_ASAP7_75t_R FILLER_154_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_914 ();
 DECAPx10_ASAP7_75t_R FILLER_154_921 ();
 DECAPx10_ASAP7_75t_R FILLER_154_943 ();
 FILLER_ASAP7_75t_R FILLER_154_965 ();
 DECAPx4_ASAP7_75t_R FILLER_154_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_983 ();
 DECAPx2_ASAP7_75t_R FILLER_154_990 ();
 DECAPx4_ASAP7_75t_R FILLER_154_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1016 ();
 DECAPx6_ASAP7_75t_R FILLER_154_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1038 ();
 DECAPx4_ASAP7_75t_R FILLER_154_1048 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_154_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1067 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1089 ();
 DECAPx6_ASAP7_75t_R FILLER_154_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1150 ();
 FILLER_ASAP7_75t_R FILLER_154_1159 ();
 DECAPx1_ASAP7_75t_R FILLER_154_1164 ();
 FILLER_ASAP7_75t_R FILLER_154_1174 ();
 FILLER_ASAP7_75t_R FILLER_154_1182 ();
 DECAPx6_ASAP7_75t_R FILLER_154_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1206 ();
 FILLER_ASAP7_75t_R FILLER_154_1213 ();
 DECAPx6_ASAP7_75t_R FILLER_154_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1242 ();
 DECAPx1_ASAP7_75t_R FILLER_154_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_1268 ();
 DECAPx6_ASAP7_75t_R FILLER_154_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_154_1289 ();
 DECAPx4_ASAP7_75t_R FILLER_154_1311 ();
 DECAPx1_ASAP7_75t_R FILLER_154_1324 ();
 FILLER_ASAP7_75t_R FILLER_154_1338 ();
 FILLER_ASAP7_75t_R FILLER_154_1346 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_154_1354 ();
 FILLER_ASAP7_75t_R FILLER_154_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_154_1371 ();
 DECAPx1_ASAP7_75t_R FILLER_155_2 ();
 DECAPx2_ASAP7_75t_R FILLER_155_12 ();
 DECAPx2_ASAP7_75t_R FILLER_155_44 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_50 ();
 FILLER_ASAP7_75t_R FILLER_155_56 ();
 FILLER_ASAP7_75t_R FILLER_155_66 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_74 ();
 DECAPx2_ASAP7_75t_R FILLER_155_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_109 ();
 DECAPx1_ASAP7_75t_R FILLER_155_116 ();
 DECAPx6_ASAP7_75t_R FILLER_155_123 ();
 DECAPx1_ASAP7_75t_R FILLER_155_143 ();
 DECAPx2_ASAP7_75t_R FILLER_155_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_183 ();
 DECAPx10_ASAP7_75t_R FILLER_155_192 ();
 DECAPx10_ASAP7_75t_R FILLER_155_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_236 ();
 DECAPx2_ASAP7_75t_R FILLER_155_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_249 ();
 FILLER_ASAP7_75t_R FILLER_155_256 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_265 ();
 FILLER_ASAP7_75t_R FILLER_155_278 ();
 FILLER_ASAP7_75t_R FILLER_155_286 ();
 FILLER_ASAP7_75t_R FILLER_155_294 ();
 DECAPx2_ASAP7_75t_R FILLER_155_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_308 ();
 FILLER_ASAP7_75t_R FILLER_155_315 ();
 DECAPx2_ASAP7_75t_R FILLER_155_328 ();
 FILLER_ASAP7_75t_R FILLER_155_334 ();
 DECAPx2_ASAP7_75t_R FILLER_155_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_368 ();
 DECAPx1_ASAP7_75t_R FILLER_155_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_379 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_386 ();
 DECAPx6_ASAP7_75t_R FILLER_155_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_406 ();
 DECAPx6_ASAP7_75t_R FILLER_155_415 ();
 DECAPx1_ASAP7_75t_R FILLER_155_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_433 ();
 FILLER_ASAP7_75t_R FILLER_155_440 ();
 DECAPx1_ASAP7_75t_R FILLER_155_445 ();
 FILLER_ASAP7_75t_R FILLER_155_475 ();
 FILLER_ASAP7_75t_R FILLER_155_483 ();
 FILLER_ASAP7_75t_R FILLER_155_493 ();
 FILLER_ASAP7_75t_R FILLER_155_501 ();
 DECAPx6_ASAP7_75t_R FILLER_155_513 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_527 ();
 DECAPx2_ASAP7_75t_R FILLER_155_536 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_542 ();
 FILLER_ASAP7_75t_R FILLER_155_548 ();
 DECAPx4_ASAP7_75t_R FILLER_155_558 ();
 FILLER_ASAP7_75t_R FILLER_155_568 ();
 FILLER_ASAP7_75t_R FILLER_155_578 ();
 DECAPx1_ASAP7_75t_R FILLER_155_586 ();
 DECAPx6_ASAP7_75t_R FILLER_155_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_611 ();
 DECAPx2_ASAP7_75t_R FILLER_155_619 ();
 DECAPx4_ASAP7_75t_R FILLER_155_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_644 ();
 DECAPx4_ASAP7_75t_R FILLER_155_657 ();
 DECAPx1_ASAP7_75t_R FILLER_155_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_679 ();
 FILLER_ASAP7_75t_R FILLER_155_686 ();
 DECAPx2_ASAP7_75t_R FILLER_155_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_704 ();
 FILLER_ASAP7_75t_R FILLER_155_708 ();
 FILLER_ASAP7_75t_R FILLER_155_719 ();
 DECAPx1_ASAP7_75t_R FILLER_155_729 ();
 DECAPx6_ASAP7_75t_R FILLER_155_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_750 ();
 DECAPx4_ASAP7_75t_R FILLER_155_759 ();
 FILLER_ASAP7_75t_R FILLER_155_769 ();
 DECAPx2_ASAP7_75t_R FILLER_155_779 ();
 FILLER_ASAP7_75t_R FILLER_155_794 ();
 FILLER_ASAP7_75t_R FILLER_155_810 ();
 DECAPx6_ASAP7_75t_R FILLER_155_818 ();
 DECAPx1_ASAP7_75t_R FILLER_155_832 ();
 DECAPx6_ASAP7_75t_R FILLER_155_843 ();
 DECAPx2_ASAP7_75t_R FILLER_155_863 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_869 ();
 FILLER_ASAP7_75t_R FILLER_155_878 ();
 FILLER_ASAP7_75t_R FILLER_155_894 ();
 FILLER_ASAP7_75t_R FILLER_155_903 ();
 FILLER_ASAP7_75t_R FILLER_155_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_922 ();
 DECAPx4_ASAP7_75t_R FILLER_155_927 ();
 FILLER_ASAP7_75t_R FILLER_155_937 ();
 DECAPx4_ASAP7_75t_R FILLER_155_945 ();
 FILLER_ASAP7_75t_R FILLER_155_955 ();
 DECAPx6_ASAP7_75t_R FILLER_155_963 ();
 DECAPx2_ASAP7_75t_R FILLER_155_977 ();
 DECAPx2_ASAP7_75t_R FILLER_155_992 ();
 FILLER_ASAP7_75t_R FILLER_155_998 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1038 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1060 ();
 FILLER_ASAP7_75t_R FILLER_155_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1078 ();
 FILLER_ASAP7_75t_R FILLER_155_1087 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1110 ();
 FILLER_ASAP7_75t_R FILLER_155_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1127 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1136 ();
 FILLER_ASAP7_75t_R FILLER_155_1150 ();
 FILLER_ASAP7_75t_R FILLER_155_1160 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1179 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1189 ();
 FILLER_ASAP7_75t_R FILLER_155_1203 ();
 FILLER_ASAP7_75t_R FILLER_155_1211 ();
 DECAPx4_ASAP7_75t_R FILLER_155_1219 ();
 FILLER_ASAP7_75t_R FILLER_155_1229 ();
 FILLER_ASAP7_75t_R FILLER_155_1234 ();
 DECAPx4_ASAP7_75t_R FILLER_155_1243 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_1253 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1263 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_155_1321 ();
 DECAPx6_ASAP7_75t_R FILLER_155_1343 ();
 DECAPx1_ASAP7_75t_R FILLER_155_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_1361 ();
 DECAPx2_ASAP7_75t_R FILLER_155_1368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_1374 ();
 FILLER_ASAP7_75t_R FILLER_156_2 ();
 DECAPx6_ASAP7_75t_R FILLER_156_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_23 ();
 FILLER_ASAP7_75t_R FILLER_156_30 ();
 DECAPx10_ASAP7_75t_R FILLER_156_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_57 ();
 DECAPx6_ASAP7_75t_R FILLER_156_64 ();
 DECAPx1_ASAP7_75t_R FILLER_156_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_82 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_89 ();
 DECAPx10_ASAP7_75t_R FILLER_156_95 ();
 DECAPx10_ASAP7_75t_R FILLER_156_117 ();
 DECAPx10_ASAP7_75t_R FILLER_156_139 ();
 FILLER_ASAP7_75t_R FILLER_156_161 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_169 ();
 DECAPx4_ASAP7_75t_R FILLER_156_175 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_185 ();
 DECAPx4_ASAP7_75t_R FILLER_156_197 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_207 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_216 ();
 DECAPx10_ASAP7_75t_R FILLER_156_227 ();
 DECAPx2_ASAP7_75t_R FILLER_156_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_255 ();
 DECAPx6_ASAP7_75t_R FILLER_156_262 ();
 DECAPx2_ASAP7_75t_R FILLER_156_276 ();
 DECAPx10_ASAP7_75t_R FILLER_156_285 ();
 DECAPx10_ASAP7_75t_R FILLER_156_307 ();
 DECAPx6_ASAP7_75t_R FILLER_156_329 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_343 ();
 DECAPx6_ASAP7_75t_R FILLER_156_352 ();
 FILLER_ASAP7_75t_R FILLER_156_392 ();
 DECAPx4_ASAP7_75t_R FILLER_156_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_407 ();
 DECAPx6_ASAP7_75t_R FILLER_156_414 ();
 DECAPx6_ASAP7_75t_R FILLER_156_434 ();
 DECAPx2_ASAP7_75t_R FILLER_156_448 ();
 FILLER_ASAP7_75t_R FILLER_156_460 ();
 FILLER_ASAP7_75t_R FILLER_156_464 ();
 DECAPx6_ASAP7_75t_R FILLER_156_472 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_486 ();
 DECAPx10_ASAP7_75t_R FILLER_156_497 ();
 FILLER_ASAP7_75t_R FILLER_156_545 ();
 FILLER_ASAP7_75t_R FILLER_156_553 ();
 DECAPx6_ASAP7_75t_R FILLER_156_563 ();
 DECAPx2_ASAP7_75t_R FILLER_156_585 ();
 FILLER_ASAP7_75t_R FILLER_156_591 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_601 ();
 FILLER_ASAP7_75t_R FILLER_156_613 ();
 DECAPx1_ASAP7_75t_R FILLER_156_623 ();
 FILLER_ASAP7_75t_R FILLER_156_655 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_663 ();
 FILLER_ASAP7_75t_R FILLER_156_674 ();
 DECAPx2_ASAP7_75t_R FILLER_156_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_688 ();
 DECAPx2_ASAP7_75t_R FILLER_156_692 ();
 FILLER_ASAP7_75t_R FILLER_156_698 ();
 DECAPx2_ASAP7_75t_R FILLER_156_709 ();
 DECAPx2_ASAP7_75t_R FILLER_156_718 ();
 FILLER_ASAP7_75t_R FILLER_156_727 ();
 FILLER_ASAP7_75t_R FILLER_156_738 ();
 DECAPx4_ASAP7_75t_R FILLER_156_748 ();
 FILLER_ASAP7_75t_R FILLER_156_758 ();
 DECAPx1_ASAP7_75t_R FILLER_156_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_772 ();
 DECAPx2_ASAP7_75t_R FILLER_156_782 ();
 DECAPx1_ASAP7_75t_R FILLER_156_799 ();
 FILLER_ASAP7_75t_R FILLER_156_812 ();
 DECAPx1_ASAP7_75t_R FILLER_156_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_824 ();
 FILLER_ASAP7_75t_R FILLER_156_832 ();
 FILLER_ASAP7_75t_R FILLER_156_841 ();
 FILLER_ASAP7_75t_R FILLER_156_850 ();
 DECAPx2_ASAP7_75t_R FILLER_156_860 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_866 ();
 FILLER_ASAP7_75t_R FILLER_156_878 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_891 ();
 DECAPx4_ASAP7_75t_R FILLER_156_902 ();
 FILLER_ASAP7_75t_R FILLER_156_912 ();
 DECAPx4_ASAP7_75t_R FILLER_156_923 ();
 FILLER_ASAP7_75t_R FILLER_156_940 ();
 DECAPx2_ASAP7_75t_R FILLER_156_949 ();
 DECAPx4_ASAP7_75t_R FILLER_156_964 ();
 FILLER_ASAP7_75t_R FILLER_156_974 ();
 DECAPx10_ASAP7_75t_R FILLER_156_984 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_156_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_156_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1035 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1045 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_1051 ();
 DECAPx4_ASAP7_75t_R FILLER_156_1063 ();
 FILLER_ASAP7_75t_R FILLER_156_1099 ();
 FILLER_ASAP7_75t_R FILLER_156_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_156_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1149 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_1156 ();
 DECAPx6_ASAP7_75t_R FILLER_156_1168 ();
 DECAPx4_ASAP7_75t_R FILLER_156_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_156_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1208 ();
 DECAPx4_ASAP7_75t_R FILLER_156_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1222 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1229 ();
 FILLER_ASAP7_75t_R FILLER_156_1244 ();
 DECAPx1_ASAP7_75t_R FILLER_156_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_1253 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_1280 ();
 FILLER_ASAP7_75t_R FILLER_156_1289 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_1294 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_1303 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1332 ();
 FILLER_ASAP7_75t_R FILLER_156_1338 ();
 DECAPx2_ASAP7_75t_R FILLER_156_1343 ();
 FILLER_ASAP7_75t_R FILLER_156_1375 ();
 FILLER_ASAP7_75t_R FILLER_157_2 ();
 DECAPx6_ASAP7_75t_R FILLER_157_9 ();
 DECAPx2_ASAP7_75t_R FILLER_157_49 ();
 DECAPx6_ASAP7_75t_R FILLER_157_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_75 ();
 DECAPx10_ASAP7_75t_R FILLER_157_82 ();
 DECAPx1_ASAP7_75t_R FILLER_157_104 ();
 FILLER_ASAP7_75t_R FILLER_157_114 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_126 ();
 FILLER_ASAP7_75t_R FILLER_157_135 ();
 FILLER_ASAP7_75t_R FILLER_157_163 ();
 DECAPx4_ASAP7_75t_R FILLER_157_171 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_181 ();
 FILLER_ASAP7_75t_R FILLER_157_190 ();
 DECAPx6_ASAP7_75t_R FILLER_157_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_209 ();
 FILLER_ASAP7_75t_R FILLER_157_218 ();
 DECAPx6_ASAP7_75t_R FILLER_157_226 ();
 DECAPx2_ASAP7_75t_R FILLER_157_246 ();
 FILLER_ASAP7_75t_R FILLER_157_252 ();
 FILLER_ASAP7_75t_R FILLER_157_257 ();
 DECAPx6_ASAP7_75t_R FILLER_157_267 ();
 FILLER_ASAP7_75t_R FILLER_157_281 ();
 DECAPx10_ASAP7_75t_R FILLER_157_289 ();
 DECAPx2_ASAP7_75t_R FILLER_157_311 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_317 ();
 DECAPx4_ASAP7_75t_R FILLER_157_326 ();
 DECAPx4_ASAP7_75t_R FILLER_157_362 ();
 FILLER_ASAP7_75t_R FILLER_157_372 ();
 FILLER_ASAP7_75t_R FILLER_157_380 ();
 DECAPx6_ASAP7_75t_R FILLER_157_385 ();
 DECAPx2_ASAP7_75t_R FILLER_157_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_405 ();
 DECAPx2_ASAP7_75t_R FILLER_157_412 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_418 ();
 DECAPx6_ASAP7_75t_R FILLER_157_447 ();
 FILLER_ASAP7_75t_R FILLER_157_461 ();
 DECAPx2_ASAP7_75t_R FILLER_157_466 ();
 DECAPx10_ASAP7_75t_R FILLER_157_475 ();
 DECAPx6_ASAP7_75t_R FILLER_157_497 ();
 DECAPx2_ASAP7_75t_R FILLER_157_517 ();
 DECAPx1_ASAP7_75t_R FILLER_157_529 ();
 FILLER_ASAP7_75t_R FILLER_157_536 ();
 DECAPx4_ASAP7_75t_R FILLER_157_541 ();
 FILLER_ASAP7_75t_R FILLER_157_551 ();
 DECAPx4_ASAP7_75t_R FILLER_157_559 ();
 DECAPx10_ASAP7_75t_R FILLER_157_575 ();
 DECAPx2_ASAP7_75t_R FILLER_157_603 ();
 FILLER_ASAP7_75t_R FILLER_157_609 ();
 DECAPx2_ASAP7_75t_R FILLER_157_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_620 ();
 DECAPx2_ASAP7_75t_R FILLER_157_627 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_633 ();
 DECAPx6_ASAP7_75t_R FILLER_157_646 ();
 DECAPx2_ASAP7_75t_R FILLER_157_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_666 ();
 DECAPx6_ASAP7_75t_R FILLER_157_673 ();
 DECAPx10_ASAP7_75t_R FILLER_157_693 ();
 DECAPx10_ASAP7_75t_R FILLER_157_715 ();
 DECAPx6_ASAP7_75t_R FILLER_157_743 ();
 DECAPx6_ASAP7_75t_R FILLER_157_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_778 ();
 DECAPx6_ASAP7_75t_R FILLER_157_785 ();
 DECAPx1_ASAP7_75t_R FILLER_157_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_803 ();
 FILLER_ASAP7_75t_R FILLER_157_812 ();
 DECAPx2_ASAP7_75t_R FILLER_157_821 ();
 DECAPx1_ASAP7_75t_R FILLER_157_834 ();
 DECAPx10_ASAP7_75t_R FILLER_157_848 ();
 DECAPx1_ASAP7_75t_R FILLER_157_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_874 ();
 DECAPx2_ASAP7_75t_R FILLER_157_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_884 ();
 DECAPx2_ASAP7_75t_R FILLER_157_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_894 ();
 DECAPx1_ASAP7_75t_R FILLER_157_902 ();
 DECAPx4_ASAP7_75t_R FILLER_157_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_924 ();
 FILLER_ASAP7_75t_R FILLER_157_927 ();
 FILLER_ASAP7_75t_R FILLER_157_939 ();
 FILLER_ASAP7_75t_R FILLER_157_947 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_952 ();
 DECAPx2_ASAP7_75t_R FILLER_157_961 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_967 ();
 DECAPx6_ASAP7_75t_R FILLER_157_980 ();
 DECAPx1_ASAP7_75t_R FILLER_157_994 ();
 FILLER_ASAP7_75t_R FILLER_157_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1013 ();
 FILLER_ASAP7_75t_R FILLER_157_1019 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1027 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1042 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_1051 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_1057 ();
 DECAPx4_ASAP7_75t_R FILLER_157_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1076 ();
 FILLER_ASAP7_75t_R FILLER_157_1087 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1092 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_1098 ();
 DECAPx1_ASAP7_75t_R FILLER_157_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1126 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_1132 ();
 FILLER_ASAP7_75t_R FILLER_157_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1154 ();
 FILLER_ASAP7_75t_R FILLER_157_1179 ();
 FILLER_ASAP7_75t_R FILLER_157_1189 ();
 DECAPx6_ASAP7_75t_R FILLER_157_1197 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_1211 ();
 DECAPx6_ASAP7_75t_R FILLER_157_1215 ();
 FILLER_ASAP7_75t_R FILLER_157_1229 ();
 FILLER_ASAP7_75t_R FILLER_157_1237 ();
 DECAPx4_ASAP7_75t_R FILLER_157_1247 ();
 FILLER_ASAP7_75t_R FILLER_157_1265 ();
 FILLER_ASAP7_75t_R FILLER_157_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_157_1278 ();
 FILLER_ASAP7_75t_R FILLER_157_1293 ();
 FILLER_ASAP7_75t_R FILLER_157_1298 ();
 FILLER_ASAP7_75t_R FILLER_157_1309 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_157_1323 ();
 DECAPx4_ASAP7_75t_R FILLER_157_1345 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_1355 ();
 FILLER_ASAP7_75t_R FILLER_157_1368 ();
 FILLER_ASAP7_75t_R FILLER_157_1375 ();
 FILLER_ASAP7_75t_R FILLER_158_2 ();
 DECAPx6_ASAP7_75t_R FILLER_158_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_23 ();
 FILLER_ASAP7_75t_R FILLER_158_30 ();
 DECAPx1_ASAP7_75t_R FILLER_158_38 ();
 FILLER_ASAP7_75t_R FILLER_158_68 ();
 FILLER_ASAP7_75t_R FILLER_158_96 ();
 DECAPx2_ASAP7_75t_R FILLER_158_104 ();
 DECAPx6_ASAP7_75t_R FILLER_158_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_130 ();
 DECAPx2_ASAP7_75t_R FILLER_158_137 ();
 DECAPx1_ASAP7_75t_R FILLER_158_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_153 ();
 DECAPx1_ASAP7_75t_R FILLER_158_180 ();
 DECAPx6_ASAP7_75t_R FILLER_158_192 ();
 FILLER_ASAP7_75t_R FILLER_158_206 ();
 DECAPx6_ASAP7_75t_R FILLER_158_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_228 ();
 DECAPx6_ASAP7_75t_R FILLER_158_255 ();
 FILLER_ASAP7_75t_R FILLER_158_275 ();
 DECAPx1_ASAP7_75t_R FILLER_158_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_284 ();
 DECAPx2_ASAP7_75t_R FILLER_158_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_302 ();
 DECAPx1_ASAP7_75t_R FILLER_158_309 ();
 FILLER_ASAP7_75t_R FILLER_158_316 ();
 DECAPx6_ASAP7_75t_R FILLER_158_326 ();
 DECAPx1_ASAP7_75t_R FILLER_158_346 ();
 DECAPx2_ASAP7_75t_R FILLER_158_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_359 ();
 DECAPx4_ASAP7_75t_R FILLER_158_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_376 ();
 DECAPx4_ASAP7_75t_R FILLER_158_385 ();
 FILLER_ASAP7_75t_R FILLER_158_395 ();
 FILLER_ASAP7_75t_R FILLER_158_403 ();
 DECAPx6_ASAP7_75t_R FILLER_158_411 ();
 DECAPx1_ASAP7_75t_R FILLER_158_431 ();
 DECAPx4_ASAP7_75t_R FILLER_158_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_448 ();
 DECAPx2_ASAP7_75t_R FILLER_158_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_461 ();
 DECAPx1_ASAP7_75t_R FILLER_158_464 ();
 FILLER_ASAP7_75t_R FILLER_158_474 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_158_484 ();
 DECAPx1_ASAP7_75t_R FILLER_158_493 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_158_503 ();
 DECAPx2_ASAP7_75t_R FILLER_158_532 ();
 DECAPx10_ASAP7_75t_R FILLER_158_541 ();
 DECAPx4_ASAP7_75t_R FILLER_158_563 ();
 DECAPx4_ASAP7_75t_R FILLER_158_579 ();
 FILLER_ASAP7_75t_R FILLER_158_589 ();
 DECAPx10_ASAP7_75t_R FILLER_158_597 ();
 DECAPx10_ASAP7_75t_R FILLER_158_619 ();
 DECAPx1_ASAP7_75t_R FILLER_158_641 ();
 DECAPx10_ASAP7_75t_R FILLER_158_653 ();
 DECAPx10_ASAP7_75t_R FILLER_158_675 ();
 DECAPx1_ASAP7_75t_R FILLER_158_697 ();
 DECAPx10_ASAP7_75t_R FILLER_158_708 ();
 FILLER_ASAP7_75t_R FILLER_158_736 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_158_746 ();
 DECAPx2_ASAP7_75t_R FILLER_158_759 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_158_765 ();
 DECAPx10_ASAP7_75t_R FILLER_158_775 ();
 DECAPx4_ASAP7_75t_R FILLER_158_797 ();
 FILLER_ASAP7_75t_R FILLER_158_807 ();
 FILLER_ASAP7_75t_R FILLER_158_816 ();
 DECAPx4_ASAP7_75t_R FILLER_158_825 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_158_835 ();
 DECAPx10_ASAP7_75t_R FILLER_158_844 ();
 DECAPx10_ASAP7_75t_R FILLER_158_866 ();
 FILLER_ASAP7_75t_R FILLER_158_888 ();
 DECAPx10_ASAP7_75t_R FILLER_158_896 ();
 DECAPx10_ASAP7_75t_R FILLER_158_918 ();
 DECAPx4_ASAP7_75t_R FILLER_158_940 ();
 DECAPx4_ASAP7_75t_R FILLER_158_960 ();
 FILLER_ASAP7_75t_R FILLER_158_976 ();
 FILLER_ASAP7_75t_R FILLER_158_988 ();
 DECAPx4_ASAP7_75t_R FILLER_158_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1010 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1023 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1035 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1049 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1062 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_158_1076 ();
 FILLER_ASAP7_75t_R FILLER_158_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_158_1090 ();
 FILLER_ASAP7_75t_R FILLER_158_1096 ();
 FILLER_ASAP7_75t_R FILLER_158_1124 ();
 FILLER_ASAP7_75t_R FILLER_158_1152 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_158_1157 ();
 FILLER_ASAP7_75t_R FILLER_158_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_158_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1180 ();
 FILLER_ASAP7_75t_R FILLER_158_1189 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1208 ();
 FILLER_ASAP7_75t_R FILLER_158_1221 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1240 ();
 DECAPx2_ASAP7_75t_R FILLER_158_1249 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1265 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1279 ();
 DECAPx4_ASAP7_75t_R FILLER_158_1286 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_158_1296 ();
 DECAPx4_ASAP7_75t_R FILLER_158_1305 ();
 FILLER_ASAP7_75t_R FILLER_158_1315 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1329 ();
 FILLER_ASAP7_75t_R FILLER_158_1333 ();
 DECAPx6_ASAP7_75t_R FILLER_158_1344 ();
 FILLER_ASAP7_75t_R FILLER_158_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_158_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_1376 ();
 FILLER_ASAP7_75t_R FILLER_159_2 ();
 FILLER_ASAP7_75t_R FILLER_159_9 ();
 DECAPx10_ASAP7_75t_R FILLER_159_16 ();
 DECAPx2_ASAP7_75t_R FILLER_159_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_47 ();
 FILLER_ASAP7_75t_R FILLER_159_54 ();
 DECAPx6_ASAP7_75t_R FILLER_159_59 ();
 FILLER_ASAP7_75t_R FILLER_159_79 ();
 FILLER_ASAP7_75t_R FILLER_159_84 ();
 FILLER_ASAP7_75t_R FILLER_159_112 ();
 DECAPx2_ASAP7_75t_R FILLER_159_122 ();
 DECAPx2_ASAP7_75t_R FILLER_159_136 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_148 ();
 DECAPx2_ASAP7_75t_R FILLER_159_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_160 ();
 FILLER_ASAP7_75t_R FILLER_159_167 ();
 DECAPx2_ASAP7_75t_R FILLER_159_172 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_178 ();
 DECAPx1_ASAP7_75t_R FILLER_159_187 ();
 FILLER_ASAP7_75t_R FILLER_159_197 ();
 DECAPx2_ASAP7_75t_R FILLER_159_225 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_231 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_240 ();
 DECAPx4_ASAP7_75t_R FILLER_159_246 ();
 FILLER_ASAP7_75t_R FILLER_159_256 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_264 ();
 DECAPx2_ASAP7_75t_R FILLER_159_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_288 ();
 DECAPx1_ASAP7_75t_R FILLER_159_315 ();
 FILLER_ASAP7_75t_R FILLER_159_327 ();
 DECAPx10_ASAP7_75t_R FILLER_159_335 ();
 DECAPx2_ASAP7_75t_R FILLER_159_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_370 ();
 FILLER_ASAP7_75t_R FILLER_159_381 ();
 FILLER_ASAP7_75t_R FILLER_159_391 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_419 ();
 DECAPx2_ASAP7_75t_R FILLER_159_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_432 ();
 FILLER_ASAP7_75t_R FILLER_159_439 ();
 DECAPx2_ASAP7_75t_R FILLER_159_467 ();
 FILLER_ASAP7_75t_R FILLER_159_495 ();
 FILLER_ASAP7_75t_R FILLER_159_507 ();
 DECAPx2_ASAP7_75t_R FILLER_159_515 ();
 DECAPx1_ASAP7_75t_R FILLER_159_543 ();
 FILLER_ASAP7_75t_R FILLER_159_553 ();
 DECAPx2_ASAP7_75t_R FILLER_159_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_569 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_576 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_585 ();
 DECAPx2_ASAP7_75t_R FILLER_159_596 ();
 FILLER_ASAP7_75t_R FILLER_159_602 ();
 FILLER_ASAP7_75t_R FILLER_159_610 ();
 DECAPx1_ASAP7_75t_R FILLER_159_618 ();
 DECAPx4_ASAP7_75t_R FILLER_159_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_641 ();
 DECAPx2_ASAP7_75t_R FILLER_159_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_655 ();
 DECAPx2_ASAP7_75t_R FILLER_159_682 ();
 DECAPx4_ASAP7_75t_R FILLER_159_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_701 ();
 FILLER_ASAP7_75t_R FILLER_159_709 ();
 DECAPx4_ASAP7_75t_R FILLER_159_723 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_733 ();
 DECAPx6_ASAP7_75t_R FILLER_159_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_760 ();
 DECAPx4_ASAP7_75t_R FILLER_159_770 ();
 DECAPx2_ASAP7_75t_R FILLER_159_789 ();
 FILLER_ASAP7_75t_R FILLER_159_795 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_806 ();
 FILLER_ASAP7_75t_R FILLER_159_815 ();
 DECAPx6_ASAP7_75t_R FILLER_159_823 ();
 DECAPx1_ASAP7_75t_R FILLER_159_837 ();
 FILLER_ASAP7_75t_R FILLER_159_847 ();
 FILLER_ASAP7_75t_R FILLER_159_859 ();
 FILLER_ASAP7_75t_R FILLER_159_873 ();
 FILLER_ASAP7_75t_R FILLER_159_883 ();
 DECAPx2_ASAP7_75t_R FILLER_159_891 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_897 ();
 DECAPx2_ASAP7_75t_R FILLER_159_908 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_922 ();
 FILLER_ASAP7_75t_R FILLER_159_927 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_939 ();
 DECAPx2_ASAP7_75t_R FILLER_159_949 ();
 FILLER_ASAP7_75t_R FILLER_159_955 ();
 FILLER_ASAP7_75t_R FILLER_159_960 ();
 DECAPx1_ASAP7_75t_R FILLER_159_988 ();
 DECAPx4_ASAP7_75t_R FILLER_159_998 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1041 ();
 DECAPx6_ASAP7_75t_R FILLER_159_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1069 ();
 DECAPx4_ASAP7_75t_R FILLER_159_1091 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_1101 ();
 FILLER_ASAP7_75t_R FILLER_159_1110 ();
 DECAPx6_ASAP7_75t_R FILLER_159_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1129 ();
 FILLER_ASAP7_75t_R FILLER_159_1143 ();
 DECAPx4_ASAP7_75t_R FILLER_159_1148 ();
 DECAPx4_ASAP7_75t_R FILLER_159_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1176 ();
 FILLER_ASAP7_75t_R FILLER_159_1203 ();
 DECAPx4_ASAP7_75t_R FILLER_159_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1221 ();
 DECAPx4_ASAP7_75t_R FILLER_159_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_159_1266 ();
 DECAPx4_ASAP7_75t_R FILLER_159_1288 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_1298 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1307 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_1313 ();
 DECAPx1_ASAP7_75t_R FILLER_159_1340 ();
 DECAPx4_ASAP7_75t_R FILLER_159_1354 ();
 FILLER_ASAP7_75t_R FILLER_159_1364 ();
 DECAPx2_ASAP7_75t_R FILLER_159_1369 ();
 FILLER_ASAP7_75t_R FILLER_159_1375 ();
 FILLER_ASAP7_75t_R FILLER_160_2 ();
 FILLER_ASAP7_75t_R FILLER_160_9 ();
 DECAPx2_ASAP7_75t_R FILLER_160_16 ();
 FILLER_ASAP7_75t_R FILLER_160_48 ();
 FILLER_ASAP7_75t_R FILLER_160_56 ();
 DECAPx10_ASAP7_75t_R FILLER_160_64 ();
 DECAPx4_ASAP7_75t_R FILLER_160_86 ();
 FILLER_ASAP7_75t_R FILLER_160_102 ();
 FILLER_ASAP7_75t_R FILLER_160_107 ();
 FILLER_ASAP7_75t_R FILLER_160_115 ();
 DECAPx2_ASAP7_75t_R FILLER_160_120 ();
 FILLER_ASAP7_75t_R FILLER_160_126 ();
 DECAPx10_ASAP7_75t_R FILLER_160_134 ();
 DECAPx10_ASAP7_75t_R FILLER_160_156 ();
 DECAPx4_ASAP7_75t_R FILLER_160_178 ();
 FILLER_ASAP7_75t_R FILLER_160_188 ();
 DECAPx2_ASAP7_75t_R FILLER_160_196 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_160_202 ();
 FILLER_ASAP7_75t_R FILLER_160_211 ();
 FILLER_ASAP7_75t_R FILLER_160_219 ();
 DECAPx2_ASAP7_75t_R FILLER_160_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_230 ();
 DECAPx2_ASAP7_75t_R FILLER_160_237 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_160_243 ();
 DECAPx1_ASAP7_75t_R FILLER_160_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_276 ();
 DECAPx1_ASAP7_75t_R FILLER_160_285 ();
 FILLER_ASAP7_75t_R FILLER_160_295 ();
 FILLER_ASAP7_75t_R FILLER_160_303 ();
 DECAPx2_ASAP7_75t_R FILLER_160_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_314 ();
 FILLER_ASAP7_75t_R FILLER_160_321 ();
 DECAPx2_ASAP7_75t_R FILLER_160_329 ();
 FILLER_ASAP7_75t_R FILLER_160_335 ();
 DECAPx4_ASAP7_75t_R FILLER_160_343 ();
 FILLER_ASAP7_75t_R FILLER_160_360 ();
 DECAPx10_ASAP7_75t_R FILLER_160_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_406 ();
 DECAPx2_ASAP7_75t_R FILLER_160_410 ();
 FILLER_ASAP7_75t_R FILLER_160_438 ();
 FILLER_ASAP7_75t_R FILLER_160_447 ();
 FILLER_ASAP7_75t_R FILLER_160_455 ();
 FILLER_ASAP7_75t_R FILLER_160_460 ();
 DECAPx1_ASAP7_75t_R FILLER_160_464 ();
 FILLER_ASAP7_75t_R FILLER_160_474 ();
 DECAPx6_ASAP7_75t_R FILLER_160_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_498 ();
 DECAPx6_ASAP7_75t_R FILLER_160_505 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_160_545 ();
 FILLER_ASAP7_75t_R FILLER_160_556 ();
 DECAPx10_ASAP7_75t_R FILLER_160_564 ();
 DECAPx2_ASAP7_75t_R FILLER_160_586 ();
 DECAPx1_ASAP7_75t_R FILLER_160_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_602 ();
 DECAPx1_ASAP7_75t_R FILLER_160_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_633 ();
 DECAPx4_ASAP7_75t_R FILLER_160_640 ();
 FILLER_ASAP7_75t_R FILLER_160_650 ();
 FILLER_ASAP7_75t_R FILLER_160_658 ();
 FILLER_ASAP7_75t_R FILLER_160_666 ();
 FILLER_ASAP7_75t_R FILLER_160_671 ();
 DECAPx2_ASAP7_75t_R FILLER_160_699 ();
 FILLER_ASAP7_75t_R FILLER_160_708 ();
 DECAPx1_ASAP7_75t_R FILLER_160_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_722 ();
 DECAPx4_ASAP7_75t_R FILLER_160_732 ();
 FILLER_ASAP7_75t_R FILLER_160_742 ();
 DECAPx1_ASAP7_75t_R FILLER_160_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_757 ();
 DECAPx6_ASAP7_75t_R FILLER_160_764 ();
 FILLER_ASAP7_75t_R FILLER_160_786 ();
 FILLER_ASAP7_75t_R FILLER_160_796 ();
 FILLER_ASAP7_75t_R FILLER_160_801 ();
 DECAPx6_ASAP7_75t_R FILLER_160_817 ();
 FILLER_ASAP7_75t_R FILLER_160_831 ();
 DECAPx1_ASAP7_75t_R FILLER_160_859 ();
 DECAPx1_ASAP7_75t_R FILLER_160_871 ();
 FILLER_ASAP7_75t_R FILLER_160_881 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_160_891 ();
 FILLER_ASAP7_75t_R FILLER_160_904 ();
 FILLER_ASAP7_75t_R FILLER_160_932 ();
 DECAPx2_ASAP7_75t_R FILLER_160_941 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_160_947 ();
 FILLER_ASAP7_75t_R FILLER_160_960 ();
 DECAPx2_ASAP7_75t_R FILLER_160_969 ();
 FILLER_ASAP7_75t_R FILLER_160_975 ();
 DECAPx4_ASAP7_75t_R FILLER_160_980 ();
 FILLER_ASAP7_75t_R FILLER_160_990 ();
 FILLER_ASAP7_75t_R FILLER_160_998 ();
 FILLER_ASAP7_75t_R FILLER_160_1010 ();
 DECAPx4_ASAP7_75t_R FILLER_160_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1041 ();
 DECAPx4_ASAP7_75t_R FILLER_160_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1093 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_160_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_160_1130 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_160_1176 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1198 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1204 ();
 FILLER_ASAP7_75t_R FILLER_160_1215 ();
 FILLER_ASAP7_75t_R FILLER_160_1223 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_160_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_160_1257 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1271 ();
 FILLER_ASAP7_75t_R FILLER_160_1283 ();
 FILLER_ASAP7_75t_R FILLER_160_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1299 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1303 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1312 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1328 ();
 DECAPx2_ASAP7_75t_R FILLER_160_1332 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_1338 ();
 DECAPx1_ASAP7_75t_R FILLER_160_1345 ();
 FILLER_ASAP7_75t_R FILLER_160_1375 ();
 FILLER_ASAP7_75t_R FILLER_161_2 ();
 DECAPx6_ASAP7_75t_R FILLER_161_9 ();
 FILLER_ASAP7_75t_R FILLER_161_29 ();
 DECAPx2_ASAP7_75t_R FILLER_161_37 ();
 DECAPx2_ASAP7_75t_R FILLER_161_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_75 ();
 DECAPx1_ASAP7_75t_R FILLER_161_82 ();
 DECAPx10_ASAP7_75t_R FILLER_161_89 ();
 DECAPx2_ASAP7_75t_R FILLER_161_111 ();
 FILLER_ASAP7_75t_R FILLER_161_123 ();
 DECAPx10_ASAP7_75t_R FILLER_161_128 ();
 DECAPx6_ASAP7_75t_R FILLER_161_150 ();
 FILLER_ASAP7_75t_R FILLER_161_164 ();
 FILLER_ASAP7_75t_R FILLER_161_172 ();
 DECAPx1_ASAP7_75t_R FILLER_161_177 ();
 FILLER_ASAP7_75t_R FILLER_161_187 ();
 DECAPx10_ASAP7_75t_R FILLER_161_192 ();
 DECAPx2_ASAP7_75t_R FILLER_161_214 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_220 ();
 FILLER_ASAP7_75t_R FILLER_161_249 ();
 DECAPx1_ASAP7_75t_R FILLER_161_257 ();
 DECAPx10_ASAP7_75t_R FILLER_161_264 ();
 DECAPx10_ASAP7_75t_R FILLER_161_286 ();
 DECAPx6_ASAP7_75t_R FILLER_161_308 ();
 DECAPx1_ASAP7_75t_R FILLER_161_322 ();
 DECAPx1_ASAP7_75t_R FILLER_161_352 ();
 DECAPx2_ASAP7_75t_R FILLER_161_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_372 ();
 FILLER_ASAP7_75t_R FILLER_161_380 ();
 DECAPx4_ASAP7_75t_R FILLER_161_388 ();
 DECAPx2_ASAP7_75t_R FILLER_161_405 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_411 ();
 FILLER_ASAP7_75t_R FILLER_161_424 ();
 DECAPx6_ASAP7_75t_R FILLER_161_438 ();
 FILLER_ASAP7_75t_R FILLER_161_452 ();
 DECAPx1_ASAP7_75t_R FILLER_161_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_484 ();
 DECAPx4_ASAP7_75t_R FILLER_161_493 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_509 ();
 DECAPx2_ASAP7_75t_R FILLER_161_515 ();
 FILLER_ASAP7_75t_R FILLER_161_521 ();
 FILLER_ASAP7_75t_R FILLER_161_529 ();
 FILLER_ASAP7_75t_R FILLER_161_537 ();
 DECAPx2_ASAP7_75t_R FILLER_161_542 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_548 ();
 DECAPx6_ASAP7_75t_R FILLER_161_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_571 ();
 DECAPx1_ASAP7_75t_R FILLER_161_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_582 ();
 FILLER_ASAP7_75t_R FILLER_161_586 ();
 DECAPx10_ASAP7_75t_R FILLER_161_596 ();
 DECAPx4_ASAP7_75t_R FILLER_161_621 ();
 FILLER_ASAP7_75t_R FILLER_161_631 ();
 FILLER_ASAP7_75t_R FILLER_161_640 ();
 FILLER_ASAP7_75t_R FILLER_161_646 ();
 FILLER_ASAP7_75t_R FILLER_161_654 ();
 FILLER_ASAP7_75t_R FILLER_161_664 ();
 DECAPx2_ASAP7_75t_R FILLER_161_669 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_675 ();
 DECAPx4_ASAP7_75t_R FILLER_161_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_696 ();
 FILLER_ASAP7_75t_R FILLER_161_706 ();
 FILLER_ASAP7_75t_R FILLER_161_714 ();
 FILLER_ASAP7_75t_R FILLER_161_722 ();
 FILLER_ASAP7_75t_R FILLER_161_732 ();
 DECAPx6_ASAP7_75t_R FILLER_161_740 ();
 DECAPx1_ASAP7_75t_R FILLER_161_754 ();
 DECAPx2_ASAP7_75t_R FILLER_161_767 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_773 ();
 DECAPx6_ASAP7_75t_R FILLER_161_782 ();
 DECAPx1_ASAP7_75t_R FILLER_161_796 ();
 DECAPx6_ASAP7_75t_R FILLER_161_803 ();
 DECAPx1_ASAP7_75t_R FILLER_161_817 ();
 FILLER_ASAP7_75t_R FILLER_161_827 ();
 DECAPx2_ASAP7_75t_R FILLER_161_837 ();
 FILLER_ASAP7_75t_R FILLER_161_843 ();
 FILLER_ASAP7_75t_R FILLER_161_853 ();
 DECAPx1_ASAP7_75t_R FILLER_161_858 ();
 DECAPx10_ASAP7_75t_R FILLER_161_888 ();
 FILLER_ASAP7_75t_R FILLER_161_918 ();
 FILLER_ASAP7_75t_R FILLER_161_923 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_927 ();
 DECAPx1_ASAP7_75t_R FILLER_161_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_941 ();
 DECAPx10_ASAP7_75t_R FILLER_161_949 ();
 DECAPx2_ASAP7_75t_R FILLER_161_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_977 ();
 DECAPx10_ASAP7_75t_R FILLER_161_986 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1022 ();
 FILLER_ASAP7_75t_R FILLER_161_1037 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1046 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_1052 ();
 FILLER_ASAP7_75t_R FILLER_161_1064 ();
 DECAPx4_ASAP7_75t_R FILLER_161_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1084 ();
 FILLER_ASAP7_75t_R FILLER_161_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1104 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_1118 ();
 FILLER_ASAP7_75t_R FILLER_161_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_161_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1158 ();
 FILLER_ASAP7_75t_R FILLER_161_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_161_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1194 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_1200 ();
 FILLER_ASAP7_75t_R FILLER_161_1229 ();
 FILLER_ASAP7_75t_R FILLER_161_1239 ();
 DECAPx6_ASAP7_75t_R FILLER_161_1244 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1258 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1288 ();
 FILLER_ASAP7_75t_R FILLER_161_1294 ();
 FILLER_ASAP7_75t_R FILLER_161_1304 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1332 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_1338 ();
 FILLER_ASAP7_75t_R FILLER_161_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_161_1355 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_1361 ();
 FILLER_ASAP7_75t_R FILLER_161_1368 ();
 DECAPx1_ASAP7_75t_R FILLER_161_1373 ();
 FILLER_ASAP7_75t_R FILLER_162_2 ();
 DECAPx10_ASAP7_75t_R FILLER_162_9 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_162_31 ();
 FILLER_ASAP7_75t_R FILLER_162_37 ();
 FILLER_ASAP7_75t_R FILLER_162_46 ();
 FILLER_ASAP7_75t_R FILLER_162_55 ();
 FILLER_ASAP7_75t_R FILLER_162_64 ();
 FILLER_ASAP7_75t_R FILLER_162_69 ();
 DECAPx2_ASAP7_75t_R FILLER_162_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_103 ();
 DECAPx1_ASAP7_75t_R FILLER_162_110 ();
 DECAPx6_ASAP7_75t_R FILLER_162_120 ();
 FILLER_ASAP7_75t_R FILLER_162_134 ();
 FILLER_ASAP7_75t_R FILLER_162_142 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_162_150 ();
 DECAPx2_ASAP7_75t_R FILLER_162_179 ();
 DECAPx4_ASAP7_75t_R FILLER_162_193 ();
 FILLER_ASAP7_75t_R FILLER_162_203 ();
 FILLER_ASAP7_75t_R FILLER_162_211 ();
 DECAPx4_ASAP7_75t_R FILLER_162_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_226 ();
 DECAPx1_ASAP7_75t_R FILLER_162_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_237 ();
 DECAPx10_ASAP7_75t_R FILLER_162_241 ();
 DECAPx10_ASAP7_75t_R FILLER_162_263 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_162_285 ();
 FILLER_ASAP7_75t_R FILLER_162_294 ();
 DECAPx4_ASAP7_75t_R FILLER_162_302 ();
 DECAPx6_ASAP7_75t_R FILLER_162_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_334 ();
 FILLER_ASAP7_75t_R FILLER_162_341 ();
 DECAPx4_ASAP7_75t_R FILLER_162_346 ();
 DECAPx1_ASAP7_75t_R FILLER_162_366 ();
 DECAPx1_ASAP7_75t_R FILLER_162_392 ();
 FILLER_ASAP7_75t_R FILLER_162_404 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_162_413 ();
 DECAPx6_ASAP7_75t_R FILLER_162_422 ();
 DECAPx2_ASAP7_75t_R FILLER_162_436 ();
 DECAPx2_ASAP7_75t_R FILLER_162_448 ();
 FILLER_ASAP7_75t_R FILLER_162_460 ();
 FILLER_ASAP7_75t_R FILLER_162_464 ();
 FILLER_ASAP7_75t_R FILLER_162_472 ();
 DECAPx1_ASAP7_75t_R FILLER_162_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_481 ();
 FILLER_ASAP7_75t_R FILLER_162_488 ();
 DECAPx1_ASAP7_75t_R FILLER_162_493 ();
 FILLER_ASAP7_75t_R FILLER_162_523 ();
 DECAPx10_ASAP7_75t_R FILLER_162_531 ();
 DECAPx2_ASAP7_75t_R FILLER_162_553 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_162_559 ();
 FILLER_ASAP7_75t_R FILLER_162_588 ();
 DECAPx6_ASAP7_75t_R FILLER_162_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_610 ();
 DECAPx6_ASAP7_75t_R FILLER_162_617 ();
 DECAPx1_ASAP7_75t_R FILLER_162_631 ();
 DECAPx10_ASAP7_75t_R FILLER_162_642 ();
 DECAPx4_ASAP7_75t_R FILLER_162_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_674 ();
 DECAPx6_ASAP7_75t_R FILLER_162_683 ();
 FILLER_ASAP7_75t_R FILLER_162_697 ();
 FILLER_ASAP7_75t_R FILLER_162_702 ();
 DECAPx1_ASAP7_75t_R FILLER_162_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_711 ();
 DECAPx4_ASAP7_75t_R FILLER_162_721 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_162_731 ();
 DECAPx4_ASAP7_75t_R FILLER_162_744 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_162_754 ();
 DECAPx10_ASAP7_75t_R FILLER_162_763 ();
 DECAPx10_ASAP7_75t_R FILLER_162_785 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_162_807 ();
 DECAPx2_ASAP7_75t_R FILLER_162_821 ();
 DECAPx2_ASAP7_75t_R FILLER_162_834 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_162_840 ();
 DECAPx10_ASAP7_75t_R FILLER_162_851 ();
 DECAPx1_ASAP7_75t_R FILLER_162_873 ();
 DECAPx10_ASAP7_75t_R FILLER_162_880 ();
 DECAPx2_ASAP7_75t_R FILLER_162_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_908 ();
 DECAPx10_ASAP7_75t_R FILLER_162_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_937 ();
 DECAPx6_ASAP7_75t_R FILLER_162_945 ();
 FILLER_ASAP7_75t_R FILLER_162_959 ();
 DECAPx6_ASAP7_75t_R FILLER_162_987 ();
 FILLER_ASAP7_75t_R FILLER_162_1001 ();
 DECAPx4_ASAP7_75t_R FILLER_162_1010 ();
 FILLER_ASAP7_75t_R FILLER_162_1020 ();
 FILLER_ASAP7_75t_R FILLER_162_1030 ();
 FILLER_ASAP7_75t_R FILLER_162_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1049 ();
 FILLER_ASAP7_75t_R FILLER_162_1058 ();
 FILLER_ASAP7_75t_R FILLER_162_1063 ();
 FILLER_ASAP7_75t_R FILLER_162_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1076 ();
 FILLER_ASAP7_75t_R FILLER_162_1085 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1148 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_162_1154 ();
 DECAPx6_ASAP7_75t_R FILLER_162_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1177 ();
 DECAPx6_ASAP7_75t_R FILLER_162_1189 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1207 ();
 FILLER_ASAP7_75t_R FILLER_162_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1221 ();
 FILLER_ASAP7_75t_R FILLER_162_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_162_1253 ();
 FILLER_ASAP7_75t_R FILLER_162_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1280 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1290 ();
 DECAPx6_ASAP7_75t_R FILLER_162_1299 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1313 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_1319 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1323 ();
 DECAPx6_ASAP7_75t_R FILLER_162_1337 ();
 DECAPx1_ASAP7_75t_R FILLER_162_1351 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_162_1363 ();
 DECAPx2_ASAP7_75t_R FILLER_162_1369 ();
 FILLER_ASAP7_75t_R FILLER_162_1375 ();
 FILLER_ASAP7_75t_R FILLER_163_2 ();
 DECAPx6_ASAP7_75t_R FILLER_163_9 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_163_23 ();
 DECAPx2_ASAP7_75t_R FILLER_163_32 ();
 FILLER_ASAP7_75t_R FILLER_163_38 ();
 FILLER_ASAP7_75t_R FILLER_163_46 ();
 FILLER_ASAP7_75t_R FILLER_163_55 ();
 FILLER_ASAP7_75t_R FILLER_163_64 ();
 DECAPx1_ASAP7_75t_R FILLER_163_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_73 ();
 DECAPx6_ASAP7_75t_R FILLER_163_80 ();
 DECAPx1_ASAP7_75t_R FILLER_163_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_98 ();
 DECAPx1_ASAP7_75t_R FILLER_163_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_129 ();
 DECAPx1_ASAP7_75t_R FILLER_163_156 ();
 FILLER_ASAP7_75t_R FILLER_163_166 ();
 FILLER_ASAP7_75t_R FILLER_163_190 ();
 FILLER_ASAP7_75t_R FILLER_163_218 ();
 DECAPx4_ASAP7_75t_R FILLER_163_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_233 ();
 DECAPx1_ASAP7_75t_R FILLER_163_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_244 ();
 DECAPx1_ASAP7_75t_R FILLER_163_251 ();
 DECAPx4_ASAP7_75t_R FILLER_163_261 ();
 DECAPx1_ASAP7_75t_R FILLER_163_277 ();
 FILLER_ASAP7_75t_R FILLER_163_307 ();
 DECAPx1_ASAP7_75t_R FILLER_163_312 ();
 DECAPx10_ASAP7_75t_R FILLER_163_324 ();
 DECAPx2_ASAP7_75t_R FILLER_163_346 ();
 FILLER_ASAP7_75t_R FILLER_163_352 ();
 FILLER_ASAP7_75t_R FILLER_163_364 ();
 DECAPx2_ASAP7_75t_R FILLER_163_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_378 ();
 FILLER_ASAP7_75t_R FILLER_163_391 ();
 DECAPx2_ASAP7_75t_R FILLER_163_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_406 ();
 FILLER_ASAP7_75t_R FILLER_163_413 ();
 DECAPx4_ASAP7_75t_R FILLER_163_423 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_163_433 ();
 FILLER_ASAP7_75t_R FILLER_163_448 ();
 DECAPx10_ASAP7_75t_R FILLER_163_457 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_163_479 ();
 DECAPx4_ASAP7_75t_R FILLER_163_488 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_163_498 ();
 DECAPx2_ASAP7_75t_R FILLER_163_507 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_163_513 ();
 FILLER_ASAP7_75t_R FILLER_163_542 ();
 DECAPx6_ASAP7_75t_R FILLER_163_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_566 ();
 DECAPx1_ASAP7_75t_R FILLER_163_573 ();
 DECAPx6_ASAP7_75t_R FILLER_163_580 ();
 FILLER_ASAP7_75t_R FILLER_163_594 ();
 FILLER_ASAP7_75t_R FILLER_163_602 ();
 FILLER_ASAP7_75t_R FILLER_163_630 ();
 DECAPx6_ASAP7_75t_R FILLER_163_639 ();
 DECAPx1_ASAP7_75t_R FILLER_163_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_657 ();
 DECAPx2_ASAP7_75t_R FILLER_163_666 ();
 DECAPx10_ASAP7_75t_R FILLER_163_682 ();
 DECAPx10_ASAP7_75t_R FILLER_163_704 ();
 DECAPx6_ASAP7_75t_R FILLER_163_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_740 ();
 DECAPx6_ASAP7_75t_R FILLER_163_747 ();
 DECAPx2_ASAP7_75t_R FILLER_163_761 ();
 FILLER_ASAP7_75t_R FILLER_163_775 ();
 FILLER_ASAP7_75t_R FILLER_163_784 ();
 DECAPx1_ASAP7_75t_R FILLER_163_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_797 ();
 DECAPx6_ASAP7_75t_R FILLER_163_805 ();
 DECAPx10_ASAP7_75t_R FILLER_163_828 ();
 DECAPx4_ASAP7_75t_R FILLER_163_850 ();
 FILLER_ASAP7_75t_R FILLER_163_860 ();
 DECAPx6_ASAP7_75t_R FILLER_163_868 ();
 DECAPx2_ASAP7_75t_R FILLER_163_882 ();
 FILLER_ASAP7_75t_R FILLER_163_898 ();
 DECAPx6_ASAP7_75t_R FILLER_163_908 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_163_922 ();
 DECAPx6_ASAP7_75t_R FILLER_163_927 ();
 DECAPx1_ASAP7_75t_R FILLER_163_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_945 ();
 DECAPx4_ASAP7_75t_R FILLER_163_958 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_163_968 ();
 FILLER_ASAP7_75t_R FILLER_163_977 ();
 DECAPx4_ASAP7_75t_R FILLER_163_987 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1009 ();
 FILLER_ASAP7_75t_R FILLER_163_1022 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1035 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1045 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1055 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1070 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1088 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_163_1105 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1123 ();
 FILLER_ASAP7_75t_R FILLER_163_1153 ();
 DECAPx4_ASAP7_75t_R FILLER_163_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1206 ();
 FILLER_ASAP7_75t_R FILLER_163_1229 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_1243 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1270 ();
 DECAPx2_ASAP7_75t_R FILLER_163_1284 ();
 FILLER_ASAP7_75t_R FILLER_163_1293 ();
 FILLER_ASAP7_75t_R FILLER_163_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_163_1309 ();
 DECAPx6_ASAP7_75t_R FILLER_163_1331 ();
 DECAPx1_ASAP7_75t_R FILLER_163_1345 ();
 FILLER_ASAP7_75t_R FILLER_163_1375 ();
 FILLER_ASAP7_75t_R FILLER_164_2 ();
 DECAPx2_ASAP7_75t_R FILLER_164_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_15 ();
 DECAPx2_ASAP7_75t_R FILLER_164_42 ();
 FILLER_ASAP7_75t_R FILLER_164_48 ();
 FILLER_ASAP7_75t_R FILLER_164_58 ();
 DECAPx1_ASAP7_75t_R FILLER_164_66 ();
 DECAPx1_ASAP7_75t_R FILLER_164_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_80 ();
 FILLER_ASAP7_75t_R FILLER_164_89 ();
 DECAPx6_ASAP7_75t_R FILLER_164_97 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_111 ();
 DECAPx10_ASAP7_75t_R FILLER_164_117 ();
 DECAPx2_ASAP7_75t_R FILLER_164_139 ();
 DECAPx1_ASAP7_75t_R FILLER_164_148 ();
 DECAPx10_ASAP7_75t_R FILLER_164_155 ();
 FILLER_ASAP7_75t_R FILLER_164_183 ();
 DECAPx2_ASAP7_75t_R FILLER_164_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_197 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_204 ();
 FILLER_ASAP7_75t_R FILLER_164_213 ();
 DECAPx2_ASAP7_75t_R FILLER_164_221 ();
 FILLER_ASAP7_75t_R FILLER_164_227 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_232 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_243 ();
 DECAPx2_ASAP7_75t_R FILLER_164_254 ();
 DECAPx2_ASAP7_75t_R FILLER_164_286 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_292 ();
 DECAPx4_ASAP7_75t_R FILLER_164_298 ();
 FILLER_ASAP7_75t_R FILLER_164_308 ();
 FILLER_ASAP7_75t_R FILLER_164_316 ();
 DECAPx4_ASAP7_75t_R FILLER_164_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_334 ();
 DECAPx6_ASAP7_75t_R FILLER_164_341 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_355 ();
 DECAPx10_ASAP7_75t_R FILLER_164_368 ();
 DECAPx4_ASAP7_75t_R FILLER_164_390 ();
 DECAPx2_ASAP7_75t_R FILLER_164_408 ();
 FILLER_ASAP7_75t_R FILLER_164_426 ();
 DECAPx4_ASAP7_75t_R FILLER_164_436 ();
 DECAPx4_ASAP7_75t_R FILLER_164_450 ();
 FILLER_ASAP7_75t_R FILLER_164_460 ();
 DECAPx2_ASAP7_75t_R FILLER_164_464 ();
 FILLER_ASAP7_75t_R FILLER_164_470 ();
 DECAPx2_ASAP7_75t_R FILLER_164_478 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_490 ();
 DECAPx6_ASAP7_75t_R FILLER_164_503 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_517 ();
 DECAPx1_ASAP7_75t_R FILLER_164_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_530 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_534 ();
 FILLER_ASAP7_75t_R FILLER_164_543 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_553 ();
 DECAPx4_ASAP7_75t_R FILLER_164_562 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_572 ();
 DECAPx4_ASAP7_75t_R FILLER_164_581 ();
 DECAPx4_ASAP7_75t_R FILLER_164_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_607 ();
 FILLER_ASAP7_75t_R FILLER_164_616 ();
 DECAPx6_ASAP7_75t_R FILLER_164_621 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_635 ();
 DECAPx4_ASAP7_75t_R FILLER_164_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_674 ();
 FILLER_ASAP7_75t_R FILLER_164_701 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_710 ();
 DECAPx1_ASAP7_75t_R FILLER_164_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_724 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_733 ();
 DECAPx2_ASAP7_75t_R FILLER_164_746 ();
 DECAPx1_ASAP7_75t_R FILLER_164_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_763 ();
 DECAPx1_ASAP7_75t_R FILLER_164_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_775 ();
 DECAPx2_ASAP7_75t_R FILLER_164_788 ();
 FILLER_ASAP7_75t_R FILLER_164_794 ();
 DECAPx4_ASAP7_75t_R FILLER_164_806 ();
 FILLER_ASAP7_75t_R FILLER_164_816 ();
 DECAPx6_ASAP7_75t_R FILLER_164_826 ();
 DECAPx1_ASAP7_75t_R FILLER_164_840 ();
 FILLER_ASAP7_75t_R FILLER_164_854 ();
 DECAPx1_ASAP7_75t_R FILLER_164_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_867 ();
 DECAPx4_ASAP7_75t_R FILLER_164_875 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_888 ();
 DECAPx4_ASAP7_75t_R FILLER_164_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_927 ();
 DECAPx4_ASAP7_75t_R FILLER_164_931 ();
 FILLER_ASAP7_75t_R FILLER_164_941 ();
 FILLER_ASAP7_75t_R FILLER_164_953 ();
 DECAPx4_ASAP7_75t_R FILLER_164_965 ();
 DECAPx6_ASAP7_75t_R FILLER_164_978 ();
 FILLER_ASAP7_75t_R FILLER_164_992 ();
 DECAPx6_ASAP7_75t_R FILLER_164_1000 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_1014 ();
 FILLER_ASAP7_75t_R FILLER_164_1026 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_164_1070 ();
 DECAPx6_ASAP7_75t_R FILLER_164_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1106 ();
 FILLER_ASAP7_75t_R FILLER_164_1118 ();
 FILLER_ASAP7_75t_R FILLER_164_1129 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1145 ();
 FILLER_ASAP7_75t_R FILLER_164_1157 ();
 DECAPx2_ASAP7_75t_R FILLER_164_1165 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_1171 ();
 FILLER_ASAP7_75t_R FILLER_164_1184 ();
 FILLER_ASAP7_75t_R FILLER_164_1194 ();
 DECAPx6_ASAP7_75t_R FILLER_164_1202 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1216 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_1246 ();
 FILLER_ASAP7_75t_R FILLER_164_1257 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1262 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_1272 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1281 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_164_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1304 ();
 DECAPx6_ASAP7_75t_R FILLER_164_1314 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1328 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_1339 ();
 FILLER_ASAP7_75t_R FILLER_164_1345 ();
 FILLER_ASAP7_75t_R FILLER_164_1356 ();
 DECAPx4_ASAP7_75t_R FILLER_164_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_1376 ();
 FILLER_ASAP7_75t_R FILLER_165_2 ();
 DECAPx4_ASAP7_75t_R FILLER_165_9 ();
 FILLER_ASAP7_75t_R FILLER_165_19 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_27 ();
 DECAPx4_ASAP7_75t_R FILLER_165_33 ();
 DECAPx1_ASAP7_75t_R FILLER_165_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_50 ();
 DECAPx2_ASAP7_75t_R FILLER_165_59 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_65 ();
 DECAPx10_ASAP7_75t_R FILLER_165_76 ();
 DECAPx4_ASAP7_75t_R FILLER_165_98 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_134 ();
 FILLER_ASAP7_75t_R FILLER_165_143 ();
 DECAPx1_ASAP7_75t_R FILLER_165_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_152 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_159 ();
 FILLER_ASAP7_75t_R FILLER_165_168 ();
 DECAPx2_ASAP7_75t_R FILLER_165_196 ();
 DECAPx2_ASAP7_75t_R FILLER_165_228 ();
 DECAPx6_ASAP7_75t_R FILLER_165_246 ();
 DECAPx1_ASAP7_75t_R FILLER_165_260 ();
 DECAPx1_ASAP7_75t_R FILLER_165_270 ();
 DECAPx1_ASAP7_75t_R FILLER_165_277 ();
 DECAPx10_ASAP7_75t_R FILLER_165_284 ();
 FILLER_ASAP7_75t_R FILLER_165_312 ();
 DECAPx4_ASAP7_75t_R FILLER_165_320 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_330 ();
 FILLER_ASAP7_75t_R FILLER_165_339 ();
 FILLER_ASAP7_75t_R FILLER_165_347 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_353 ();
 DECAPx6_ASAP7_75t_R FILLER_165_362 ();
 DECAPx1_ASAP7_75t_R FILLER_165_376 ();
 FILLER_ASAP7_75t_R FILLER_165_388 ();
 DECAPx1_ASAP7_75t_R FILLER_165_396 ();
 DECAPx2_ASAP7_75t_R FILLER_165_410 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_416 ();
 FILLER_ASAP7_75t_R FILLER_165_431 ();
 DECAPx10_ASAP7_75t_R FILLER_165_439 ();
 DECAPx4_ASAP7_75t_R FILLER_165_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_497 ();
 DECAPx6_ASAP7_75t_R FILLER_165_504 ();
 DECAPx1_ASAP7_75t_R FILLER_165_518 ();
 DECAPx2_ASAP7_75t_R FILLER_165_528 ();
 FILLER_ASAP7_75t_R FILLER_165_534 ();
 FILLER_ASAP7_75t_R FILLER_165_539 ();
 FILLER_ASAP7_75t_R FILLER_165_547 ();
 FILLER_ASAP7_75t_R FILLER_165_555 ();
 FILLER_ASAP7_75t_R FILLER_165_563 ();
 FILLER_ASAP7_75t_R FILLER_165_571 ();
 DECAPx6_ASAP7_75t_R FILLER_165_579 ();
 DECAPx4_ASAP7_75t_R FILLER_165_599 ();
 FILLER_ASAP7_75t_R FILLER_165_617 ();
 FILLER_ASAP7_75t_R FILLER_165_625 ();
 DECAPx1_ASAP7_75t_R FILLER_165_645 ();
 FILLER_ASAP7_75t_R FILLER_165_655 ();
 DECAPx4_ASAP7_75t_R FILLER_165_665 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_675 ();
 DECAPx1_ASAP7_75t_R FILLER_165_685 ();
 DECAPx2_ASAP7_75t_R FILLER_165_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_698 ();
 FILLER_ASAP7_75t_R FILLER_165_706 ();
 DECAPx2_ASAP7_75t_R FILLER_165_720 ();
 FILLER_ASAP7_75t_R FILLER_165_726 ();
 FILLER_ASAP7_75t_R FILLER_165_740 ();
 DECAPx2_ASAP7_75t_R FILLER_165_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_754 ();
 FILLER_ASAP7_75t_R FILLER_165_765 ();
 DECAPx2_ASAP7_75t_R FILLER_165_777 ();
 DECAPx1_ASAP7_75t_R FILLER_165_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_793 ();
 DECAPx4_ASAP7_75t_R FILLER_165_806 ();
 FILLER_ASAP7_75t_R FILLER_165_822 ();
 DECAPx2_ASAP7_75t_R FILLER_165_832 ();
 FILLER_ASAP7_75t_R FILLER_165_838 ();
 FILLER_ASAP7_75t_R FILLER_165_843 ();
 DECAPx6_ASAP7_75t_R FILLER_165_855 ();
 DECAPx1_ASAP7_75t_R FILLER_165_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_873 ();
 DECAPx1_ASAP7_75t_R FILLER_165_884 ();
 DECAPx2_ASAP7_75t_R FILLER_165_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_904 ();
 DECAPx2_ASAP7_75t_R FILLER_165_908 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_922 ();
 FILLER_ASAP7_75t_R FILLER_165_927 ();
 DECAPx10_ASAP7_75t_R FILLER_165_939 ();
 DECAPx1_ASAP7_75t_R FILLER_165_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_965 ();
 FILLER_ASAP7_75t_R FILLER_165_972 ();
 FILLER_ASAP7_75t_R FILLER_165_980 ();
 DECAPx1_ASAP7_75t_R FILLER_165_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_992 ();
 FILLER_ASAP7_75t_R FILLER_165_1001 ();
 DECAPx4_ASAP7_75t_R FILLER_165_1006 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_1019 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1032 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_1046 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1069 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1101 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_1107 ();
 FILLER_ASAP7_75t_R FILLER_165_1113 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1118 ();
 FILLER_ASAP7_75t_R FILLER_165_1132 ();
 FILLER_ASAP7_75t_R FILLER_165_1160 ();
 FILLER_ASAP7_75t_R FILLER_165_1169 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1174 ();
 FILLER_ASAP7_75t_R FILLER_165_1188 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1193 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1202 ();
 DECAPx1_ASAP7_75t_R FILLER_165_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1220 ();
 DECAPx1_ASAP7_75t_R FILLER_165_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1233 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1237 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_1251 ();
 FILLER_ASAP7_75t_R FILLER_165_1257 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1268 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_1274 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1299 ();
 FILLER_ASAP7_75t_R FILLER_165_1306 ();
 FILLER_ASAP7_75t_R FILLER_165_1334 ();
 FILLER_ASAP7_75t_R FILLER_165_1342 ();
 DECAPx6_ASAP7_75t_R FILLER_165_1350 ();
 DECAPx2_ASAP7_75t_R FILLER_165_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_1376 ();
 FILLER_ASAP7_75t_R FILLER_166_2 ();
 FILLER_ASAP7_75t_R FILLER_166_9 ();
 DECAPx1_ASAP7_75t_R FILLER_166_16 ();
 FILLER_ASAP7_75t_R FILLER_166_26 ();
 DECAPx10_ASAP7_75t_R FILLER_166_34 ();
 DECAPx6_ASAP7_75t_R FILLER_166_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_70 ();
 DECAPx2_ASAP7_75t_R FILLER_166_77 ();
 FILLER_ASAP7_75t_R FILLER_166_83 ();
 FILLER_ASAP7_75t_R FILLER_166_91 ();
 FILLER_ASAP7_75t_R FILLER_166_101 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_111 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_120 ();
 DECAPx1_ASAP7_75t_R FILLER_166_126 ();
 FILLER_ASAP7_75t_R FILLER_166_156 ();
 DECAPx4_ASAP7_75t_R FILLER_166_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_174 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_181 ();
 DECAPx6_ASAP7_75t_R FILLER_166_187 ();
 DECAPx2_ASAP7_75t_R FILLER_166_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_207 ();
 FILLER_ASAP7_75t_R FILLER_166_211 ();
 DECAPx1_ASAP7_75t_R FILLER_166_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_223 ();
 FILLER_ASAP7_75t_R FILLER_166_231 ();
 FILLER_ASAP7_75t_R FILLER_166_240 ();
 DECAPx10_ASAP7_75t_R FILLER_166_248 ();
 DECAPx6_ASAP7_75t_R FILLER_166_270 ();
 DECAPx1_ASAP7_75t_R FILLER_166_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_296 ();
 FILLER_ASAP7_75t_R FILLER_166_323 ();
 DECAPx2_ASAP7_75t_R FILLER_166_351 ();
 FILLER_ASAP7_75t_R FILLER_166_357 ();
 DECAPx2_ASAP7_75t_R FILLER_166_369 ();
 FILLER_ASAP7_75t_R FILLER_166_375 ();
 DECAPx2_ASAP7_75t_R FILLER_166_389 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_395 ();
 DECAPx10_ASAP7_75t_R FILLER_166_406 ();
 DECAPx4_ASAP7_75t_R FILLER_166_428 ();
 FILLER_ASAP7_75t_R FILLER_166_443 ();
 DECAPx1_ASAP7_75t_R FILLER_166_451 ();
 DECAPx1_ASAP7_75t_R FILLER_166_458 ();
 FILLER_ASAP7_75t_R FILLER_166_464 ();
 DECAPx1_ASAP7_75t_R FILLER_166_472 ();
 DECAPx6_ASAP7_75t_R FILLER_166_479 ();
 FILLER_ASAP7_75t_R FILLER_166_500 ();
 FILLER_ASAP7_75t_R FILLER_166_509 ();
 DECAPx10_ASAP7_75t_R FILLER_166_537 ();
 DECAPx6_ASAP7_75t_R FILLER_166_559 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_573 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_584 ();
 DECAPx6_ASAP7_75t_R FILLER_166_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_609 ();
 DECAPx4_ASAP7_75t_R FILLER_166_616 ();
 FILLER_ASAP7_75t_R FILLER_166_626 ();
 FILLER_ASAP7_75t_R FILLER_166_637 ();
 DECAPx2_ASAP7_75t_R FILLER_166_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_652 ();
 FILLER_ASAP7_75t_R FILLER_166_659 ();
 DECAPx2_ASAP7_75t_R FILLER_166_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_670 ();
 FILLER_ASAP7_75t_R FILLER_166_681 ();
 DECAPx1_ASAP7_75t_R FILLER_166_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_690 ();
 FILLER_ASAP7_75t_R FILLER_166_701 ();
 DECAPx2_ASAP7_75t_R FILLER_166_710 ();
 FILLER_ASAP7_75t_R FILLER_166_724 ();
 DECAPx6_ASAP7_75t_R FILLER_166_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_747 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_756 ();
 DECAPx2_ASAP7_75t_R FILLER_166_781 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_787 ();
 FILLER_ASAP7_75t_R FILLER_166_796 ();
 FILLER_ASAP7_75t_R FILLER_166_804 ();
 DECAPx2_ASAP7_75t_R FILLER_166_809 ();
 FILLER_ASAP7_75t_R FILLER_166_815 ();
 FILLER_ASAP7_75t_R FILLER_166_823 ();
 DECAPx6_ASAP7_75t_R FILLER_166_851 ();
 DECAPx1_ASAP7_75t_R FILLER_166_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_869 ();
 DECAPx10_ASAP7_75t_R FILLER_166_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_902 ();
 FILLER_ASAP7_75t_R FILLER_166_911 ();
 DECAPx1_ASAP7_75t_R FILLER_166_939 ();
 DECAPx4_ASAP7_75t_R FILLER_166_952 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_962 ();
 DECAPx2_ASAP7_75t_R FILLER_166_973 ();
 DECAPx2_ASAP7_75t_R FILLER_166_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_993 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1008 ();
 FILLER_ASAP7_75t_R FILLER_166_1012 ();
 FILLER_ASAP7_75t_R FILLER_166_1028 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1041 ();
 FILLER_ASAP7_75t_R FILLER_166_1047 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1055 ();
 FILLER_ASAP7_75t_R FILLER_166_1068 ();
 FILLER_ASAP7_75t_R FILLER_166_1073 ();
 FILLER_ASAP7_75t_R FILLER_166_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1124 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1152 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1166 ();
 FILLER_ASAP7_75t_R FILLER_166_1176 ();
 DECAPx4_ASAP7_75t_R FILLER_166_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1194 ();
 FILLER_ASAP7_75t_R FILLER_166_1204 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1212 ();
 FILLER_ASAP7_75t_R FILLER_166_1225 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1230 ();
 FILLER_ASAP7_75t_R FILLER_166_1236 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1248 ();
 FILLER_ASAP7_75t_R FILLER_166_1257 ();
 FILLER_ASAP7_75t_R FILLER_166_1279 ();
 FILLER_ASAP7_75t_R FILLER_166_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_166_1299 ();
 FILLER_ASAP7_75t_R FILLER_166_1306 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1316 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_166_1326 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1348 ();
 FILLER_ASAP7_75t_R FILLER_166_1360 ();
 DECAPx2_ASAP7_75t_R FILLER_166_1368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_1374 ();
 FILLER_ASAP7_75t_R FILLER_167_2 ();
 DECAPx1_ASAP7_75t_R FILLER_167_9 ();
 FILLER_ASAP7_75t_R FILLER_167_39 ();
 DECAPx1_ASAP7_75t_R FILLER_167_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_48 ();
 FILLER_ASAP7_75t_R FILLER_167_57 ();
 FILLER_ASAP7_75t_R FILLER_167_65 ();
 FILLER_ASAP7_75t_R FILLER_167_73 ();
 DECAPx2_ASAP7_75t_R FILLER_167_81 ();
 FILLER_ASAP7_75t_R FILLER_167_93 ();
 FILLER_ASAP7_75t_R FILLER_167_101 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_167_109 ();
 FILLER_ASAP7_75t_R FILLER_167_118 ();
 DECAPx4_ASAP7_75t_R FILLER_167_123 ();
 DECAPx6_ASAP7_75t_R FILLER_167_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_153 ();
 FILLER_ASAP7_75t_R FILLER_167_162 ();
 DECAPx2_ASAP7_75t_R FILLER_167_172 ();
 DECAPx1_ASAP7_75t_R FILLER_167_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_188 ();
 DECAPx6_ASAP7_75t_R FILLER_167_195 ();
 DECAPx2_ASAP7_75t_R FILLER_167_209 ();
 FILLER_ASAP7_75t_R FILLER_167_222 ();
 FILLER_ASAP7_75t_R FILLER_167_231 ();
 FILLER_ASAP7_75t_R FILLER_167_240 ();
 DECAPx1_ASAP7_75t_R FILLER_167_245 ();
 FILLER_ASAP7_75t_R FILLER_167_257 ();
 FILLER_ASAP7_75t_R FILLER_167_265 ();
 FILLER_ASAP7_75t_R FILLER_167_273 ();
 FILLER_ASAP7_75t_R FILLER_167_281 ();
 FILLER_ASAP7_75t_R FILLER_167_291 ();
 FILLER_ASAP7_75t_R FILLER_167_299 ();
 FILLER_ASAP7_75t_R FILLER_167_309 ();
 FILLER_ASAP7_75t_R FILLER_167_318 ();
 DECAPx6_ASAP7_75t_R FILLER_167_323 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_167_337 ();
 DECAPx2_ASAP7_75t_R FILLER_167_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_349 ();
 DECAPx1_ASAP7_75t_R FILLER_167_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_357 ();
 FILLER_ASAP7_75t_R FILLER_167_364 ();
 DECAPx2_ASAP7_75t_R FILLER_167_373 ();
 DECAPx6_ASAP7_75t_R FILLER_167_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_405 ();
 DECAPx10_ASAP7_75t_R FILLER_167_412 ();
 DECAPx2_ASAP7_75t_R FILLER_167_434 ();
 FILLER_ASAP7_75t_R FILLER_167_466 ();
 FILLER_ASAP7_75t_R FILLER_167_474 ();
 DECAPx2_ASAP7_75t_R FILLER_167_484 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_167_496 ();
 FILLER_ASAP7_75t_R FILLER_167_521 ();
 FILLER_ASAP7_75t_R FILLER_167_529 ();
 DECAPx4_ASAP7_75t_R FILLER_167_534 ();
 FILLER_ASAP7_75t_R FILLER_167_544 ();
 DECAPx6_ASAP7_75t_R FILLER_167_554 ();
 DECAPx2_ASAP7_75t_R FILLER_167_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_574 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_167_581 ();
 FILLER_ASAP7_75t_R FILLER_167_590 ();
 FILLER_ASAP7_75t_R FILLER_167_614 ();
 DECAPx6_ASAP7_75t_R FILLER_167_619 ();
 DECAPx1_ASAP7_75t_R FILLER_167_633 ();
 DECAPx10_ASAP7_75t_R FILLER_167_645 ();
 DECAPx2_ASAP7_75t_R FILLER_167_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_673 ();
 DECAPx2_ASAP7_75t_R FILLER_167_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_686 ();
 FILLER_ASAP7_75t_R FILLER_167_694 ();
 DECAPx10_ASAP7_75t_R FILLER_167_718 ();
 DECAPx6_ASAP7_75t_R FILLER_167_750 ();
 DECAPx1_ASAP7_75t_R FILLER_167_764 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_167_774 ();
 DECAPx6_ASAP7_75t_R FILLER_167_783 ();
 FILLER_ASAP7_75t_R FILLER_167_797 ();
 DECAPx6_ASAP7_75t_R FILLER_167_811 ();
 DECAPx1_ASAP7_75t_R FILLER_167_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_829 ();
 FILLER_ASAP7_75t_R FILLER_167_838 ();
 DECAPx6_ASAP7_75t_R FILLER_167_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_857 ();
 DECAPx10_ASAP7_75t_R FILLER_167_884 ();
 DECAPx6_ASAP7_75t_R FILLER_167_906 ();
 DECAPx1_ASAP7_75t_R FILLER_167_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_924 ();
 FILLER_ASAP7_75t_R FILLER_167_927 ();
 DECAPx4_ASAP7_75t_R FILLER_167_939 ();
 DECAPx2_ASAP7_75t_R FILLER_167_956 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_167_962 ();
 DECAPx2_ASAP7_75t_R FILLER_167_975 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_167_981 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1023 ();
 FILLER_ASAP7_75t_R FILLER_167_1043 ();
 FILLER_ASAP7_75t_R FILLER_167_1048 ();
 FILLER_ASAP7_75t_R FILLER_167_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1088 ();
 FILLER_ASAP7_75t_R FILLER_167_1092 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1111 ();
 FILLER_ASAP7_75t_R FILLER_167_1138 ();
 FILLER_ASAP7_75t_R FILLER_167_1150 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1158 ();
 DECAPx1_ASAP7_75t_R FILLER_167_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1176 ();
 FILLER_ASAP7_75t_R FILLER_167_1187 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1195 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1204 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_167_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_167_1219 ();
 DECAPx4_ASAP7_75t_R FILLER_167_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1251 ();
 DECAPx4_ASAP7_75t_R FILLER_167_1262 ();
 FILLER_ASAP7_75t_R FILLER_167_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_167_1300 ();
 DECAPx6_ASAP7_75t_R FILLER_167_1322 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_1342 ();
 DECAPx4_ASAP7_75t_R FILLER_167_1349 ();
 DECAPx2_ASAP7_75t_R FILLER_167_1369 ();
 FILLER_ASAP7_75t_R FILLER_167_1375 ();
 FILLER_ASAP7_75t_R FILLER_168_2 ();
 DECAPx6_ASAP7_75t_R FILLER_168_9 ();
 DECAPx1_ASAP7_75t_R FILLER_168_23 ();
 DECAPx6_ASAP7_75t_R FILLER_168_30 ();
 DECAPx2_ASAP7_75t_R FILLER_168_44 ();
 DECAPx10_ASAP7_75t_R FILLER_168_58 ();
 DECAPx10_ASAP7_75t_R FILLER_168_80 ();
 DECAPx6_ASAP7_75t_R FILLER_168_102 ();
 DECAPx1_ASAP7_75t_R FILLER_168_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_120 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_127 ();
 DECAPx2_ASAP7_75t_R FILLER_168_136 ();
 FILLER_ASAP7_75t_R FILLER_168_149 ();
 FILLER_ASAP7_75t_R FILLER_168_158 ();
 DECAPx2_ASAP7_75t_R FILLER_168_167 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_199 ();
 FILLER_ASAP7_75t_R FILLER_168_228 ();
 DECAPx1_ASAP7_75t_R FILLER_168_237 ();
 DECAPx1_ASAP7_75t_R FILLER_168_247 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_254 ();
 DECAPx2_ASAP7_75t_R FILLER_168_283 ();
 DECAPx6_ASAP7_75t_R FILLER_168_311 ();
 DECAPx1_ASAP7_75t_R FILLER_168_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_329 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_336 ();
 DECAPx1_ASAP7_75t_R FILLER_168_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_349 ();
 FILLER_ASAP7_75t_R FILLER_168_356 ();
 FILLER_ASAP7_75t_R FILLER_168_364 ();
 FILLER_ASAP7_75t_R FILLER_168_373 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_378 ();
 DECAPx6_ASAP7_75t_R FILLER_168_388 ();
 DECAPx1_ASAP7_75t_R FILLER_168_402 ();
 DECAPx4_ASAP7_75t_R FILLER_168_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_424 ();
 DECAPx4_ASAP7_75t_R FILLER_168_431 ();
 FILLER_ASAP7_75t_R FILLER_168_441 ();
 DECAPx4_ASAP7_75t_R FILLER_168_449 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_459 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_464 ();
 DECAPx2_ASAP7_75t_R FILLER_168_470 ();
 FILLER_ASAP7_75t_R FILLER_168_476 ();
 DECAPx10_ASAP7_75t_R FILLER_168_500 ();
 DECAPx6_ASAP7_75t_R FILLER_168_522 ();
 DECAPx1_ASAP7_75t_R FILLER_168_536 ();
 FILLER_ASAP7_75t_R FILLER_168_546 ();
 DECAPx1_ASAP7_75t_R FILLER_168_556 ();
 FILLER_ASAP7_75t_R FILLER_168_566 ();
 DECAPx1_ASAP7_75t_R FILLER_168_574 ();
 DECAPx4_ASAP7_75t_R FILLER_168_581 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_591 ();
 DECAPx2_ASAP7_75t_R FILLER_168_600 ();
 DECAPx1_ASAP7_75t_R FILLER_168_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_613 ();
 FILLER_ASAP7_75t_R FILLER_168_621 ();
 DECAPx2_ASAP7_75t_R FILLER_168_629 ();
 FILLER_ASAP7_75t_R FILLER_168_638 ();
 DECAPx6_ASAP7_75t_R FILLER_168_647 ();
 DECAPx2_ASAP7_75t_R FILLER_168_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_693 ();
 DECAPx10_ASAP7_75t_R FILLER_168_700 ();
 DECAPx6_ASAP7_75t_R FILLER_168_722 ();
 DECAPx1_ASAP7_75t_R FILLER_168_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_740 ();
 DECAPx4_ASAP7_75t_R FILLER_168_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_759 ();
 DECAPx2_ASAP7_75t_R FILLER_168_772 ();
 FILLER_ASAP7_75t_R FILLER_168_778 ();
 DECAPx2_ASAP7_75t_R FILLER_168_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_794 ();
 DECAPx10_ASAP7_75t_R FILLER_168_801 ();
 DECAPx10_ASAP7_75t_R FILLER_168_823 ();
 DECAPx2_ASAP7_75t_R FILLER_168_845 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_851 ();
 FILLER_ASAP7_75t_R FILLER_168_860 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_870 ();
 FILLER_ASAP7_75t_R FILLER_168_876 ();
 DECAPx2_ASAP7_75t_R FILLER_168_888 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_894 ();
 FILLER_ASAP7_75t_R FILLER_168_907 ();
 DECAPx1_ASAP7_75t_R FILLER_168_915 ();
 FILLER_ASAP7_75t_R FILLER_168_945 ();
 DECAPx2_ASAP7_75t_R FILLER_168_955 ();
 FILLER_ASAP7_75t_R FILLER_168_961 ();
 DECAPx6_ASAP7_75t_R FILLER_168_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_985 ();
 DECAPx1_ASAP7_75t_R FILLER_168_994 ();
 DECAPx10_ASAP7_75t_R FILLER_168_1001 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1023 ();
 FILLER_ASAP7_75t_R FILLER_168_1033 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_168_1057 ();
 DECAPx6_ASAP7_75t_R FILLER_168_1079 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1099 ();
 DECAPx6_ASAP7_75t_R FILLER_168_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1120 ();
 DECAPx6_ASAP7_75t_R FILLER_168_1129 ();
 DECAPx1_ASAP7_75t_R FILLER_168_1143 ();
 FILLER_ASAP7_75t_R FILLER_168_1150 ();
 DECAPx6_ASAP7_75t_R FILLER_168_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_1175 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1202 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_1212 ();
 DECAPx2_ASAP7_75t_R FILLER_168_1218 ();
 FILLER_ASAP7_75t_R FILLER_168_1224 ();
 FILLER_ASAP7_75t_R FILLER_168_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_168_1240 ();
 DECAPx1_ASAP7_75t_R FILLER_168_1262 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1276 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_1286 ();
 DECAPx6_ASAP7_75t_R FILLER_168_1292 ();
 DECAPx4_ASAP7_75t_R FILLER_168_1314 ();
 FILLER_ASAP7_75t_R FILLER_168_1333 ();
 FILLER_ASAP7_75t_R FILLER_168_1338 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_1346 ();
 FILLER_ASAP7_75t_R FILLER_168_1375 ();
 FILLER_ASAP7_75t_R FILLER_169_2 ();
 FILLER_ASAP7_75t_R FILLER_169_9 ();
 DECAPx4_ASAP7_75t_R FILLER_169_16 ();
 DECAPx6_ASAP7_75t_R FILLER_169_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_46 ();
 FILLER_ASAP7_75t_R FILLER_169_53 ();
 DECAPx4_ASAP7_75t_R FILLER_169_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_71 ();
 DECAPx6_ASAP7_75t_R FILLER_169_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_92 ();
 FILLER_ASAP7_75t_R FILLER_169_99 ();
 DECAPx2_ASAP7_75t_R FILLER_169_107 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_113 ();
 DECAPx2_ASAP7_75t_R FILLER_169_142 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_148 ();
 FILLER_ASAP7_75t_R FILLER_169_158 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_167 ();
 DECAPx4_ASAP7_75t_R FILLER_169_176 ();
 FILLER_ASAP7_75t_R FILLER_169_186 ();
 DECAPx6_ASAP7_75t_R FILLER_169_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_205 ();
 DECAPx1_ASAP7_75t_R FILLER_169_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_216 ();
 DECAPx6_ASAP7_75t_R FILLER_169_220 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_234 ();
 FILLER_ASAP7_75t_R FILLER_169_263 ();
 FILLER_ASAP7_75t_R FILLER_169_271 ();
 DECAPx6_ASAP7_75t_R FILLER_169_276 ();
 DECAPx2_ASAP7_75t_R FILLER_169_290 ();
 DECAPx6_ASAP7_75t_R FILLER_169_302 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_322 ();
 DECAPx2_ASAP7_75t_R FILLER_169_351 ();
 FILLER_ASAP7_75t_R FILLER_169_357 ();
 FILLER_ASAP7_75t_R FILLER_169_367 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_376 ();
 DECAPx2_ASAP7_75t_R FILLER_169_387 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_393 ();
 FILLER_ASAP7_75t_R FILLER_169_403 ();
 DECAPx2_ASAP7_75t_R FILLER_169_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_419 ();
 DECAPx2_ASAP7_75t_R FILLER_169_430 ();
 FILLER_ASAP7_75t_R FILLER_169_436 ();
 DECAPx1_ASAP7_75t_R FILLER_169_464 ();
 FILLER_ASAP7_75t_R FILLER_169_474 ();
 FILLER_ASAP7_75t_R FILLER_169_484 ();
 DECAPx1_ASAP7_75t_R FILLER_169_492 ();
 DECAPx1_ASAP7_75t_R FILLER_169_522 ();
 FILLER_ASAP7_75t_R FILLER_169_532 ();
 FILLER_ASAP7_75t_R FILLER_169_537 ();
 FILLER_ASAP7_75t_R FILLER_169_542 ();
 DECAPx2_ASAP7_75t_R FILLER_169_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_556 ();
 FILLER_ASAP7_75t_R FILLER_169_583 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_588 ();
 DECAPx2_ASAP7_75t_R FILLER_169_617 ();
 FILLER_ASAP7_75t_R FILLER_169_635 ();
 DECAPx1_ASAP7_75t_R FILLER_169_643 ();
 FILLER_ASAP7_75t_R FILLER_169_659 ();
 FILLER_ASAP7_75t_R FILLER_169_665 ();
 FILLER_ASAP7_75t_R FILLER_169_677 ();
 DECAPx4_ASAP7_75t_R FILLER_169_682 ();
 FILLER_ASAP7_75t_R FILLER_169_700 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_710 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_716 ();
 DECAPx4_ASAP7_75t_R FILLER_169_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_735 ();
 DECAPx6_ASAP7_75t_R FILLER_169_762 ();
 DECAPx2_ASAP7_75t_R FILLER_169_786 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_792 ();
 DECAPx1_ASAP7_75t_R FILLER_169_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_808 ();
 DECAPx2_ASAP7_75t_R FILLER_169_812 ();
 FILLER_ASAP7_75t_R FILLER_169_818 ();
 FILLER_ASAP7_75t_R FILLER_169_846 ();
 DECAPx2_ASAP7_75t_R FILLER_169_854 ();
 DECAPx4_ASAP7_75t_R FILLER_169_868 ();
 FILLER_ASAP7_75t_R FILLER_169_904 ();
 DECAPx2_ASAP7_75t_R FILLER_169_916 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_922 ();
 FILLER_ASAP7_75t_R FILLER_169_927 ();
 FILLER_ASAP7_75t_R FILLER_169_937 ();
 DECAPx2_ASAP7_75t_R FILLER_169_942 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_948 ();
 DECAPx10_ASAP7_75t_R FILLER_169_977 ();
 DECAPx10_ASAP7_75t_R FILLER_169_999 ();
 DECAPx6_ASAP7_75t_R FILLER_169_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_169_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1059 ();
 DECAPx4_ASAP7_75t_R FILLER_169_1063 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_1073 ();
 FILLER_ASAP7_75t_R FILLER_169_1083 ();
 DECAPx1_ASAP7_75t_R FILLER_169_1088 ();
 DECAPx1_ASAP7_75t_R FILLER_169_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1142 ();
 FILLER_ASAP7_75t_R FILLER_169_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1158 ();
 FILLER_ASAP7_75t_R FILLER_169_1188 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_1193 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_1206 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1219 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_1225 ();
 FILLER_ASAP7_75t_R FILLER_169_1238 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_169_1262 ();
 DECAPx1_ASAP7_75t_R FILLER_169_1284 ();
 DECAPx4_ASAP7_75t_R FILLER_169_1298 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_1316 ();
 FILLER_ASAP7_75t_R FILLER_169_1322 ();
 FILLER_ASAP7_75t_R FILLER_169_1333 ();
 FILLER_ASAP7_75t_R FILLER_169_1341 ();
 FILLER_ASAP7_75t_R FILLER_169_1353 ();
 DECAPx1_ASAP7_75t_R FILLER_169_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_1365 ();
 DECAPx2_ASAP7_75t_R FILLER_169_1369 ();
 FILLER_ASAP7_75t_R FILLER_169_1375 ();
 FILLER_ASAP7_75t_R FILLER_170_2 ();
 DECAPx2_ASAP7_75t_R FILLER_170_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_15 ();
 DECAPx10_ASAP7_75t_R FILLER_170_42 ();
 DECAPx1_ASAP7_75t_R FILLER_170_90 ();
 DECAPx4_ASAP7_75t_R FILLER_170_120 ();
 DECAPx2_ASAP7_75t_R FILLER_170_133 ();
 FILLER_ASAP7_75t_R FILLER_170_139 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_144 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_155 ();
 DECAPx2_ASAP7_75t_R FILLER_170_164 ();
 FILLER_ASAP7_75t_R FILLER_170_170 ();
 DECAPx4_ASAP7_75t_R FILLER_170_179 ();
 FILLER_ASAP7_75t_R FILLER_170_189 ();
 DECAPx10_ASAP7_75t_R FILLER_170_197 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_225 ();
 DECAPx2_ASAP7_75t_R FILLER_170_231 ();
 FILLER_ASAP7_75t_R FILLER_170_237 ();
 DECAPx10_ASAP7_75t_R FILLER_170_245 ();
 DECAPx6_ASAP7_75t_R FILLER_170_267 ();
 DECAPx2_ASAP7_75t_R FILLER_170_281 ();
 FILLER_ASAP7_75t_R FILLER_170_295 ();
 DECAPx1_ASAP7_75t_R FILLER_170_305 ();
 DECAPx1_ASAP7_75t_R FILLER_170_335 ();
 DECAPx1_ASAP7_75t_R FILLER_170_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_346 ();
 FILLER_ASAP7_75t_R FILLER_170_355 ();
 FILLER_ASAP7_75t_R FILLER_170_379 ();
 DECAPx2_ASAP7_75t_R FILLER_170_395 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_401 ();
 DECAPx1_ASAP7_75t_R FILLER_170_412 ();
 FILLER_ASAP7_75t_R FILLER_170_423 ();
 FILLER_ASAP7_75t_R FILLER_170_447 ();
 FILLER_ASAP7_75t_R FILLER_170_455 ();
 FILLER_ASAP7_75t_R FILLER_170_460 ();
 DECAPx2_ASAP7_75t_R FILLER_170_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_470 ();
 FILLER_ASAP7_75t_R FILLER_170_479 ();
 DECAPx2_ASAP7_75t_R FILLER_170_487 ();
 FILLER_ASAP7_75t_R FILLER_170_499 ();
 FILLER_ASAP7_75t_R FILLER_170_507 ();
 FILLER_ASAP7_75t_R FILLER_170_512 ();
 DECAPx6_ASAP7_75t_R FILLER_170_540 ();
 DECAPx6_ASAP7_75t_R FILLER_170_560 ();
 DECAPx4_ASAP7_75t_R FILLER_170_580 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_590 ();
 DECAPx10_ASAP7_75t_R FILLER_170_599 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_621 ();
 FILLER_ASAP7_75t_R FILLER_170_631 ();
 FILLER_ASAP7_75t_R FILLER_170_657 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_665 ();
 DECAPx10_ASAP7_75t_R FILLER_170_674 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_696 ();
 FILLER_ASAP7_75t_R FILLER_170_725 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_735 ();
 DECAPx1_ASAP7_75t_R FILLER_170_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_750 ();
 DECAPx4_ASAP7_75t_R FILLER_170_754 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_764 ();
 DECAPx4_ASAP7_75t_R FILLER_170_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_789 ();
 DECAPx2_ASAP7_75t_R FILLER_170_796 ();
 FILLER_ASAP7_75t_R FILLER_170_828 ();
 FILLER_ASAP7_75t_R FILLER_170_840 ();
 DECAPx10_ASAP7_75t_R FILLER_170_852 ();
 DECAPx4_ASAP7_75t_R FILLER_170_874 ();
 FILLER_ASAP7_75t_R FILLER_170_892 ();
 DECAPx6_ASAP7_75t_R FILLER_170_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_911 ();
 FILLER_ASAP7_75t_R FILLER_170_918 ();
 DECAPx10_ASAP7_75t_R FILLER_170_928 ();
 DECAPx6_ASAP7_75t_R FILLER_170_950 ();
 FILLER_ASAP7_75t_R FILLER_170_964 ();
 DECAPx4_ASAP7_75t_R FILLER_170_969 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_979 ();
 DECAPx2_ASAP7_75t_R FILLER_170_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_996 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1013 ();
 FILLER_ASAP7_75t_R FILLER_170_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1029 ();
 FILLER_ASAP7_75t_R FILLER_170_1035 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_1043 ();
 FILLER_ASAP7_75t_R FILLER_170_1072 ();
 DECAPx4_ASAP7_75t_R FILLER_170_1100 ();
 FILLER_ASAP7_75t_R FILLER_170_1110 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1125 ();
 DECAPx4_ASAP7_75t_R FILLER_170_1152 ();
 FILLER_ASAP7_75t_R FILLER_170_1162 ();
 FILLER_ASAP7_75t_R FILLER_170_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_170_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1198 ();
 DECAPx6_ASAP7_75t_R FILLER_170_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_1222 ();
 FILLER_ASAP7_75t_R FILLER_170_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_170_1277 ();
 FILLER_ASAP7_75t_R FILLER_170_1299 ();
 FILLER_ASAP7_75t_R FILLER_170_1327 ();
 DECAPx1_ASAP7_75t_R FILLER_170_1339 ();
 DECAPx2_ASAP7_75t_R FILLER_170_1369 ();
 FILLER_ASAP7_75t_R FILLER_170_1375 ();
 FILLER_ASAP7_75t_R FILLER_171_2 ();
 FILLER_ASAP7_75t_R FILLER_171_9 ();
 DECAPx1_ASAP7_75t_R FILLER_171_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_20 ();
 DECAPx1_ASAP7_75t_R FILLER_171_27 ();
 DECAPx6_ASAP7_75t_R FILLER_171_34 ();
 DECAPx6_ASAP7_75t_R FILLER_171_54 ();
 DECAPx1_ASAP7_75t_R FILLER_171_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_78 ();
 DECAPx6_ASAP7_75t_R FILLER_171_82 ();
 FILLER_ASAP7_75t_R FILLER_171_96 ();
 DECAPx1_ASAP7_75t_R FILLER_171_104 ();
 DECAPx4_ASAP7_75t_R FILLER_171_111 ();
 FILLER_ASAP7_75t_R FILLER_171_121 ();
 DECAPx4_ASAP7_75t_R FILLER_171_129 ();
 FILLER_ASAP7_75t_R FILLER_171_145 ();
 DECAPx2_ASAP7_75t_R FILLER_171_155 ();
 FILLER_ASAP7_75t_R FILLER_171_161 ();
 DECAPx6_ASAP7_75t_R FILLER_171_169 ();
 FILLER_ASAP7_75t_R FILLER_171_183 ();
 FILLER_ASAP7_75t_R FILLER_171_191 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_201 ();
 FILLER_ASAP7_75t_R FILLER_171_211 ();
 DECAPx6_ASAP7_75t_R FILLER_171_239 ();
 DECAPx1_ASAP7_75t_R FILLER_171_253 ();
 DECAPx4_ASAP7_75t_R FILLER_171_263 ();
 FILLER_ASAP7_75t_R FILLER_171_276 ();
 DECAPx1_ASAP7_75t_R FILLER_171_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_288 ();
 DECAPx6_ASAP7_75t_R FILLER_171_295 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_309 ();
 DECAPx2_ASAP7_75t_R FILLER_171_318 ();
 DECAPx4_ASAP7_75t_R FILLER_171_327 ();
 FILLER_ASAP7_75t_R FILLER_171_337 ();
 FILLER_ASAP7_75t_R FILLER_171_342 ();
 FILLER_ASAP7_75t_R FILLER_171_350 ();
 FILLER_ASAP7_75t_R FILLER_171_358 ();
 FILLER_ASAP7_75t_R FILLER_171_367 ();
 DECAPx2_ASAP7_75t_R FILLER_171_391 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_397 ();
 FILLER_ASAP7_75t_R FILLER_171_410 ();
 FILLER_ASAP7_75t_R FILLER_171_434 ();
 FILLER_ASAP7_75t_R FILLER_171_442 ();
 DECAPx6_ASAP7_75t_R FILLER_171_450 ();
 DECAPx2_ASAP7_75t_R FILLER_171_464 ();
 DECAPx6_ASAP7_75t_R FILLER_171_478 ();
 DECAPx2_ASAP7_75t_R FILLER_171_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_498 ();
 DECAPx6_ASAP7_75t_R FILLER_171_505 ();
 DECAPx2_ASAP7_75t_R FILLER_171_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_531 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_538 ();
 DECAPx1_ASAP7_75t_R FILLER_171_547 ();
 DECAPx2_ASAP7_75t_R FILLER_171_558 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_564 ();
 DECAPx2_ASAP7_75t_R FILLER_171_593 ();
 FILLER_ASAP7_75t_R FILLER_171_599 ();
 DECAPx2_ASAP7_75t_R FILLER_171_607 ();
 FILLER_ASAP7_75t_R FILLER_171_613 ();
 FILLER_ASAP7_75t_R FILLER_171_637 ();
 FILLER_ASAP7_75t_R FILLER_171_651 ();
 DECAPx6_ASAP7_75t_R FILLER_171_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_674 ();
 DECAPx4_ASAP7_75t_R FILLER_171_678 ();
 DECAPx6_ASAP7_75t_R FILLER_171_694 ();
 DECAPx2_ASAP7_75t_R FILLER_171_708 ();
 DECAPx2_ASAP7_75t_R FILLER_171_717 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_723 ();
 DECAPx2_ASAP7_75t_R FILLER_171_729 ();
 DECAPx6_ASAP7_75t_R FILLER_171_741 ();
 DECAPx1_ASAP7_75t_R FILLER_171_755 ();
 DECAPx2_ASAP7_75t_R FILLER_171_768 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_774 ();
 DECAPx6_ASAP7_75t_R FILLER_171_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_803 ();
 DECAPx2_ASAP7_75t_R FILLER_171_810 ();
 FILLER_ASAP7_75t_R FILLER_171_819 ();
 DECAPx1_ASAP7_75t_R FILLER_171_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_833 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_837 ();
 DECAPx2_ASAP7_75t_R FILLER_171_849 ();
 DECAPx2_ASAP7_75t_R FILLER_171_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_871 ();
 DECAPx6_ASAP7_75t_R FILLER_171_882 ();
 DECAPx2_ASAP7_75t_R FILLER_171_896 ();
 DECAPx4_ASAP7_75t_R FILLER_171_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_922 ();
 DECAPx2_ASAP7_75t_R FILLER_171_927 ();
 DECAPx1_ASAP7_75t_R FILLER_171_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_943 ();
 DECAPx2_ASAP7_75t_R FILLER_171_954 ();
 FILLER_ASAP7_75t_R FILLER_171_960 ();
 FILLER_ASAP7_75t_R FILLER_171_970 ();
 DECAPx2_ASAP7_75t_R FILLER_171_978 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1023 ();
 FILLER_ASAP7_75t_R FILLER_171_1032 ();
 FILLER_ASAP7_75t_R FILLER_171_1040 ();
 DECAPx1_ASAP7_75t_R FILLER_171_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1049 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_1060 ();
 FILLER_ASAP7_75t_R FILLER_171_1070 ();
 FILLER_ASAP7_75t_R FILLER_171_1078 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1105 ();
 FILLER_ASAP7_75t_R FILLER_171_1111 ();
 DECAPx6_ASAP7_75t_R FILLER_171_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1140 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_1154 ();
 FILLER_ASAP7_75t_R FILLER_171_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_171_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1205 ();
 DECAPx4_ASAP7_75t_R FILLER_171_1227 ();
 FILLER_ASAP7_75t_R FILLER_171_1240 ();
 FILLER_ASAP7_75t_R FILLER_171_1248 ();
 FILLER_ASAP7_75t_R FILLER_171_1260 ();
 FILLER_ASAP7_75t_R FILLER_171_1265 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_1270 ();
 DECAPx1_ASAP7_75t_R FILLER_171_1282 ();
 FILLER_ASAP7_75t_R FILLER_171_1292 ();
 FILLER_ASAP7_75t_R FILLER_171_1297 ();
 DECAPx6_ASAP7_75t_R FILLER_171_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_171_1319 ();
 DECAPx6_ASAP7_75t_R FILLER_171_1341 ();
 FILLER_ASAP7_75t_R FILLER_171_1355 ();
 DECAPx6_ASAP7_75t_R FILLER_171_1360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_1374 ();
 FILLER_ASAP7_75t_R FILLER_172_2 ();
 DECAPx6_ASAP7_75t_R FILLER_172_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_23 ();
 DECAPx4_ASAP7_75t_R FILLER_172_30 ();
 DECAPx6_ASAP7_75t_R FILLER_172_66 ();
 DECAPx1_ASAP7_75t_R FILLER_172_80 ();
 DECAPx10_ASAP7_75t_R FILLER_172_90 ();
 FILLER_ASAP7_75t_R FILLER_172_112 ();
 DECAPx1_ASAP7_75t_R FILLER_172_140 ();
 DECAPx2_ASAP7_75t_R FILLER_172_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_156 ();
 DECAPx6_ASAP7_75t_R FILLER_172_163 ();
 DECAPx1_ASAP7_75t_R FILLER_172_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_187 ();
 FILLER_ASAP7_75t_R FILLER_172_191 ();
 FILLER_ASAP7_75t_R FILLER_172_201 ();
 DECAPx2_ASAP7_75t_R FILLER_172_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_215 ();
 DECAPx2_ASAP7_75t_R FILLER_172_222 ();
 FILLER_ASAP7_75t_R FILLER_172_228 ();
 DECAPx1_ASAP7_75t_R FILLER_172_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_244 ();
 FILLER_ASAP7_75t_R FILLER_172_271 ();
 DECAPx10_ASAP7_75t_R FILLER_172_299 ();
 FILLER_ASAP7_75t_R FILLER_172_321 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_329 ();
 DECAPx6_ASAP7_75t_R FILLER_172_338 ();
 DECAPx2_ASAP7_75t_R FILLER_172_360 ();
 FILLER_ASAP7_75t_R FILLER_172_374 ();
 DECAPx1_ASAP7_75t_R FILLER_172_382 ();
 FILLER_ASAP7_75t_R FILLER_172_408 ();
 DECAPx1_ASAP7_75t_R FILLER_172_418 ();
 FILLER_ASAP7_75t_R FILLER_172_432 ();
 FILLER_ASAP7_75t_R FILLER_172_460 ();
 DECAPx2_ASAP7_75t_R FILLER_172_464 ();
 FILLER_ASAP7_75t_R FILLER_172_478 ();
 FILLER_ASAP7_75t_R FILLER_172_502 ();
 DECAPx6_ASAP7_75t_R FILLER_172_510 ();
 FILLER_ASAP7_75t_R FILLER_172_524 ();
 FILLER_ASAP7_75t_R FILLER_172_552 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_561 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_567 ();
 DECAPx1_ASAP7_75t_R FILLER_172_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_580 ();
 DECAPx2_ASAP7_75t_R FILLER_172_584 ();
 FILLER_ASAP7_75t_R FILLER_172_590 ();
 FILLER_ASAP7_75t_R FILLER_172_598 ();
 DECAPx10_ASAP7_75t_R FILLER_172_626 ();
 DECAPx1_ASAP7_75t_R FILLER_172_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_652 ();
 DECAPx4_ASAP7_75t_R FILLER_172_663 ();
 DECAPx2_ASAP7_75t_R FILLER_172_683 ();
 FILLER_ASAP7_75t_R FILLER_172_689 ();
 DECAPx10_ASAP7_75t_R FILLER_172_705 ();
 DECAPx10_ASAP7_75t_R FILLER_172_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_749 ();
 FILLER_ASAP7_75t_R FILLER_172_762 ();
 DECAPx2_ASAP7_75t_R FILLER_172_772 ();
 FILLER_ASAP7_75t_R FILLER_172_792 ();
 DECAPx10_ASAP7_75t_R FILLER_172_800 ();
 DECAPx10_ASAP7_75t_R FILLER_172_822 ();
 DECAPx2_ASAP7_75t_R FILLER_172_851 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_857 ();
 DECAPx4_ASAP7_75t_R FILLER_172_886 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_896 ();
 DECAPx2_ASAP7_75t_R FILLER_172_909 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_915 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_924 ();
 FILLER_ASAP7_75t_R FILLER_172_935 ();
 DECAPx6_ASAP7_75t_R FILLER_172_963 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_983 ();
 DECAPx1_ASAP7_75t_R FILLER_172_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_998 ();
 DECAPx6_ASAP7_75t_R FILLER_172_1002 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1027 ();
 FILLER_ASAP7_75t_R FILLER_172_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1107 ();
 FILLER_ASAP7_75t_R FILLER_172_1114 ();
 DECAPx1_ASAP7_75t_R FILLER_172_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_1128 ();
 FILLER_ASAP7_75t_R FILLER_172_1155 ();
 FILLER_ASAP7_75t_R FILLER_172_1160 ();
 FILLER_ASAP7_75t_R FILLER_172_1171 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1185 ();
 FILLER_ASAP7_75t_R FILLER_172_1210 ();
 FILLER_ASAP7_75t_R FILLER_172_1215 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1220 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_1226 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_172_1257 ();
 DECAPx1_ASAP7_75t_R FILLER_172_1271 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1281 ();
 FILLER_ASAP7_75t_R FILLER_172_1287 ();
 FILLER_ASAP7_75t_R FILLER_172_1298 ();
 FILLER_ASAP7_75t_R FILLER_172_1303 ();
 FILLER_ASAP7_75t_R FILLER_172_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_172_1346 ();
 DECAPx2_ASAP7_75t_R FILLER_172_1368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_1374 ();
 FILLER_ASAP7_75t_R FILLER_173_2 ();
 DECAPx2_ASAP7_75t_R FILLER_173_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_15 ();
 FILLER_ASAP7_75t_R FILLER_173_42 ();
 DECAPx1_ASAP7_75t_R FILLER_173_50 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_57 ();
 DECAPx1_ASAP7_75t_R FILLER_173_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_70 ();
 FILLER_ASAP7_75t_R FILLER_173_77 ();
 FILLER_ASAP7_75t_R FILLER_173_82 ();
 DECAPx10_ASAP7_75t_R FILLER_173_92 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_114 ();
 DECAPx1_ASAP7_75t_R FILLER_173_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_127 ();
 DECAPx10_ASAP7_75t_R FILLER_173_131 ();
 DECAPx4_ASAP7_75t_R FILLER_173_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_163 ();
 DECAPx10_ASAP7_75t_R FILLER_173_190 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_212 ();
 DECAPx2_ASAP7_75t_R FILLER_173_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_228 ();
 DECAPx6_ASAP7_75t_R FILLER_173_235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_249 ();
 DECAPx1_ASAP7_75t_R FILLER_173_258 ();
 DECAPx4_ASAP7_75t_R FILLER_173_265 ();
 DECAPx2_ASAP7_75t_R FILLER_173_281 ();
 DECAPx4_ASAP7_75t_R FILLER_173_290 ();
 DECAPx1_ASAP7_75t_R FILLER_173_306 ();
 DECAPx2_ASAP7_75t_R FILLER_173_313 ();
 DECAPx1_ASAP7_75t_R FILLER_173_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_349 ();
 FILLER_ASAP7_75t_R FILLER_173_356 ();
 FILLER_ASAP7_75t_R FILLER_173_364 ();
 DECAPx2_ASAP7_75t_R FILLER_173_373 ();
 FILLER_ASAP7_75t_R FILLER_173_379 ();
 FILLER_ASAP7_75t_R FILLER_173_407 ();
 DECAPx1_ASAP7_75t_R FILLER_173_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_419 ();
 FILLER_ASAP7_75t_R FILLER_173_427 ();
 DECAPx2_ASAP7_75t_R FILLER_173_435 ();
 DECAPx2_ASAP7_75t_R FILLER_173_447 ();
 DECAPx4_ASAP7_75t_R FILLER_173_456 ();
 FILLER_ASAP7_75t_R FILLER_173_472 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_480 ();
 FILLER_ASAP7_75t_R FILLER_173_489 ();
 FILLER_ASAP7_75t_R FILLER_173_499 ();
 DECAPx4_ASAP7_75t_R FILLER_173_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_517 ();
 DECAPx6_ASAP7_75t_R FILLER_173_524 ();
 FILLER_ASAP7_75t_R FILLER_173_538 ();
 DECAPx2_ASAP7_75t_R FILLER_173_543 ();
 DECAPx1_ASAP7_75t_R FILLER_173_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_579 ();
 DECAPx2_ASAP7_75t_R FILLER_173_583 ();
 FILLER_ASAP7_75t_R FILLER_173_589 ();
 FILLER_ASAP7_75t_R FILLER_173_599 ();
 FILLER_ASAP7_75t_R FILLER_173_615 ();
 DECAPx4_ASAP7_75t_R FILLER_173_620 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_630 ();
 DECAPx2_ASAP7_75t_R FILLER_173_639 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_645 ();
 FILLER_ASAP7_75t_R FILLER_173_674 ();
 DECAPx2_ASAP7_75t_R FILLER_173_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_689 ();
 DECAPx2_ASAP7_75t_R FILLER_173_698 ();
 FILLER_ASAP7_75t_R FILLER_173_712 ();
 DECAPx1_ASAP7_75t_R FILLER_173_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_725 ();
 DECAPx1_ASAP7_75t_R FILLER_173_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_738 ();
 DECAPx2_ASAP7_75t_R FILLER_173_747 ();
 FILLER_ASAP7_75t_R FILLER_173_753 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_761 ();
 DECAPx6_ASAP7_75t_R FILLER_173_776 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_790 ();
 FILLER_ASAP7_75t_R FILLER_173_801 ();
 DECAPx4_ASAP7_75t_R FILLER_173_813 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_823 ();
 DECAPx2_ASAP7_75t_R FILLER_173_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_842 ();
 DECAPx2_ASAP7_75t_R FILLER_173_850 ();
 FILLER_ASAP7_75t_R FILLER_173_866 ();
 FILLER_ASAP7_75t_R FILLER_173_876 ();
 DECAPx4_ASAP7_75t_R FILLER_173_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_891 ();
 DECAPx2_ASAP7_75t_R FILLER_173_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_924 ();
 FILLER_ASAP7_75t_R FILLER_173_927 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_937 ();
 DECAPx1_ASAP7_75t_R FILLER_173_948 ();
 DECAPx2_ASAP7_75t_R FILLER_173_955 ();
 DECAPx2_ASAP7_75t_R FILLER_173_968 ();
 FILLER_ASAP7_75t_R FILLER_173_974 ();
 FILLER_ASAP7_75t_R FILLER_173_983 ();
 FILLER_ASAP7_75t_R FILLER_173_991 ();
 DECAPx4_ASAP7_75t_R FILLER_173_996 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1043 ();
 FILLER_ASAP7_75t_R FILLER_173_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_173_1080 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_1086 ();
 FILLER_ASAP7_75t_R FILLER_173_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_173_1103 ();
 FILLER_ASAP7_75t_R FILLER_173_1109 ();
 DECAPx4_ASAP7_75t_R FILLER_173_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1127 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1154 ();
 FILLER_ASAP7_75t_R FILLER_173_1176 ();
 FILLER_ASAP7_75t_R FILLER_173_1181 ();
 DECAPx4_ASAP7_75t_R FILLER_173_1191 ();
 FILLER_ASAP7_75t_R FILLER_173_1209 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1229 ();
 FILLER_ASAP7_75t_R FILLER_173_1251 ();
 DECAPx4_ASAP7_75t_R FILLER_173_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_173_1276 ();
 DECAPx4_ASAP7_75t_R FILLER_173_1288 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_1298 ();
 FILLER_ASAP7_75t_R FILLER_173_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_173_1335 ();
 DECAPx6_ASAP7_75t_R FILLER_173_1357 ();
 DECAPx2_ASAP7_75t_R FILLER_173_1371 ();
 DECAPx6_ASAP7_75t_R FILLER_174_2 ();
 DECAPx1_ASAP7_75t_R FILLER_174_16 ();
 DECAPx1_ASAP7_75t_R FILLER_174_26 ();
 DECAPx4_ASAP7_75t_R FILLER_174_33 ();
 FILLER_ASAP7_75t_R FILLER_174_43 ();
 DECAPx4_ASAP7_75t_R FILLER_174_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_58 ();
 FILLER_ASAP7_75t_R FILLER_174_67 ();
 DECAPx1_ASAP7_75t_R FILLER_174_77 ();
 FILLER_ASAP7_75t_R FILLER_174_87 ();
 FILLER_ASAP7_75t_R FILLER_174_95 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_174_106 ();
 DECAPx1_ASAP7_75t_R FILLER_174_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_119 ();
 FILLER_ASAP7_75t_R FILLER_174_123 ();
 DECAPx6_ASAP7_75t_R FILLER_174_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_145 ();
 DECAPx2_ASAP7_75t_R FILLER_174_154 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_174_160 ();
 FILLER_ASAP7_75t_R FILLER_174_169 ();
 FILLER_ASAP7_75t_R FILLER_174_177 ();
 DECAPx6_ASAP7_75t_R FILLER_174_182 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_174_196 ();
 FILLER_ASAP7_75t_R FILLER_174_205 ();
 FILLER_ASAP7_75t_R FILLER_174_214 ();
 DECAPx1_ASAP7_75t_R FILLER_174_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_230 ();
 DECAPx2_ASAP7_75t_R FILLER_174_237 ();
 FILLER_ASAP7_75t_R FILLER_174_243 ();
 DECAPx6_ASAP7_75t_R FILLER_174_251 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_174_265 ();
 DECAPx1_ASAP7_75t_R FILLER_174_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_278 ();
 DECAPx4_ASAP7_75t_R FILLER_174_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_295 ();
 DECAPx4_ASAP7_75t_R FILLER_174_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_332 ();
 DECAPx10_ASAP7_75t_R FILLER_174_336 ();
 DECAPx4_ASAP7_75t_R FILLER_174_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_374 ();
 DECAPx1_ASAP7_75t_R FILLER_174_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_385 ();
 FILLER_ASAP7_75t_R FILLER_174_408 ();
 DECAPx4_ASAP7_75t_R FILLER_174_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_446 ();
 DECAPx2_ASAP7_75t_R FILLER_174_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_174_459 ();
 FILLER_ASAP7_75t_R FILLER_174_464 ();
 DECAPx1_ASAP7_75t_R FILLER_174_469 ();
 DECAPx2_ASAP7_75t_R FILLER_174_479 ();
 DECAPx1_ASAP7_75t_R FILLER_174_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_492 ();
 DECAPx2_ASAP7_75t_R FILLER_174_501 ();
 FILLER_ASAP7_75t_R FILLER_174_507 ();
 DECAPx2_ASAP7_75t_R FILLER_174_535 ();
 FILLER_ASAP7_75t_R FILLER_174_541 ();
 FILLER_ASAP7_75t_R FILLER_174_549 ();
 FILLER_ASAP7_75t_R FILLER_174_558 ();
 DECAPx10_ASAP7_75t_R FILLER_174_567 ();
 FILLER_ASAP7_75t_R FILLER_174_589 ();
 FILLER_ASAP7_75t_R FILLER_174_599 ();
 DECAPx2_ASAP7_75t_R FILLER_174_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_613 ();
 FILLER_ASAP7_75t_R FILLER_174_624 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_174_632 ();
 DECAPx2_ASAP7_75t_R FILLER_174_645 ();
 DECAPx1_ASAP7_75t_R FILLER_174_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_661 ();
 DECAPx2_ASAP7_75t_R FILLER_174_665 ();
 FILLER_ASAP7_75t_R FILLER_174_671 ();
 DECAPx6_ASAP7_75t_R FILLER_174_676 ();
 DECAPx1_ASAP7_75t_R FILLER_174_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_694 ();
 FILLER_ASAP7_75t_R FILLER_174_702 ();
 DECAPx1_ASAP7_75t_R FILLER_174_710 ();
 FILLER_ASAP7_75t_R FILLER_174_740 ();
 DECAPx4_ASAP7_75t_R FILLER_174_751 ();
 DECAPx2_ASAP7_75t_R FILLER_174_773 ();
 DECAPx6_ASAP7_75t_R FILLER_174_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_801 ();
 FILLER_ASAP7_75t_R FILLER_174_828 ();
 FILLER_ASAP7_75t_R FILLER_174_838 ();
 DECAPx10_ASAP7_75t_R FILLER_174_848 ();
 DECAPx2_ASAP7_75t_R FILLER_174_870 ();
 FILLER_ASAP7_75t_R FILLER_174_876 ();
 DECAPx4_ASAP7_75t_R FILLER_174_886 ();
 FILLER_ASAP7_75t_R FILLER_174_904 ();
 DECAPx10_ASAP7_75t_R FILLER_174_909 ();
 DECAPx4_ASAP7_75t_R FILLER_174_931 ();
 DECAPx2_ASAP7_75t_R FILLER_174_944 ();
 DECAPx6_ASAP7_75t_R FILLER_174_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_970 ();
 FILLER_ASAP7_75t_R FILLER_174_983 ();
 FILLER_ASAP7_75t_R FILLER_174_991 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1019 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_174_1025 ();
 FILLER_ASAP7_75t_R FILLER_174_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1065 ();
 FILLER_ASAP7_75t_R FILLER_174_1071 ();
 FILLER_ASAP7_75t_R FILLER_174_1081 ();
 DECAPx4_ASAP7_75t_R FILLER_174_1091 ();
 FILLER_ASAP7_75t_R FILLER_174_1107 ();
 DECAPx6_ASAP7_75t_R FILLER_174_1115 ();
 DECAPx1_ASAP7_75t_R FILLER_174_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1141 ();
 FILLER_ASAP7_75t_R FILLER_174_1145 ();
 DECAPx6_ASAP7_75t_R FILLER_174_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1170 ();
 FILLER_ASAP7_75t_R FILLER_174_1177 ();
 FILLER_ASAP7_75t_R FILLER_174_1188 ();
 DECAPx4_ASAP7_75t_R FILLER_174_1193 ();
 FILLER_ASAP7_75t_R FILLER_174_1209 ();
 DECAPx4_ASAP7_75t_R FILLER_174_1217 ();
 FILLER_ASAP7_75t_R FILLER_174_1235 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_1249 ();
 FILLER_ASAP7_75t_R FILLER_174_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_174_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1277 ();
 DECAPx6_ASAP7_75t_R FILLER_174_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_174_1308 ();
 FILLER_ASAP7_75t_R FILLER_174_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_174_1349 ();
 DECAPx2_ASAP7_75t_R FILLER_174_1371 ();
 DECAPx10_ASAP7_75t_R FILLER_175_2 ();
 DECAPx4_ASAP7_75t_R FILLER_175_24 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_40 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_46 ();
 FILLER_ASAP7_75t_R FILLER_175_52 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_62 ();
 FILLER_ASAP7_75t_R FILLER_175_71 ();
 DECAPx4_ASAP7_75t_R FILLER_175_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_89 ();
 DECAPx4_ASAP7_75t_R FILLER_175_96 ();
 DECAPx2_ASAP7_75t_R FILLER_175_132 ();
 FILLER_ASAP7_75t_R FILLER_175_144 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_154 ();
 FILLER_ASAP7_75t_R FILLER_175_163 ();
 DECAPx2_ASAP7_75t_R FILLER_175_171 ();
 FILLER_ASAP7_75t_R FILLER_175_177 ();
 DECAPx2_ASAP7_75t_R FILLER_175_185 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_194 ();
 DECAPx10_ASAP7_75t_R FILLER_175_205 ();
 FILLER_ASAP7_75t_R FILLER_175_233 ();
 FILLER_ASAP7_75t_R FILLER_175_261 ();
 DECAPx2_ASAP7_75t_R FILLER_175_289 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_295 ();
 FILLER_ASAP7_75t_R FILLER_175_304 ();
 DECAPx4_ASAP7_75t_R FILLER_175_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_322 ();
 DECAPx2_ASAP7_75t_R FILLER_175_326 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_332 ();
 DECAPx4_ASAP7_75t_R FILLER_175_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_351 ();
 DECAPx2_ASAP7_75t_R FILLER_175_378 ();
 FILLER_ASAP7_75t_R FILLER_175_384 ();
 DECAPx1_ASAP7_75t_R FILLER_175_392 ();
 DECAPx2_ASAP7_75t_R FILLER_175_399 ();
 DECAPx2_ASAP7_75t_R FILLER_175_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_414 ();
 DECAPx4_ASAP7_75t_R FILLER_175_421 ();
 FILLER_ASAP7_75t_R FILLER_175_457 ();
 DECAPx4_ASAP7_75t_R FILLER_175_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_495 ();
 DECAPx4_ASAP7_75t_R FILLER_175_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_512 ();
 DECAPx1_ASAP7_75t_R FILLER_175_519 ();
 DECAPx2_ASAP7_75t_R FILLER_175_526 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_532 ();
 FILLER_ASAP7_75t_R FILLER_175_541 ();
 FILLER_ASAP7_75t_R FILLER_175_549 ();
 DECAPx4_ASAP7_75t_R FILLER_175_558 ();
 FILLER_ASAP7_75t_R FILLER_175_568 ();
 FILLER_ASAP7_75t_R FILLER_175_573 ();
 DECAPx4_ASAP7_75t_R FILLER_175_581 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_591 ();
 DECAPx2_ASAP7_75t_R FILLER_175_600 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_606 ();
 DECAPx1_ASAP7_75t_R FILLER_175_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_623 ();
 DECAPx2_ASAP7_75t_R FILLER_175_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_637 ();
 DECAPx2_ASAP7_75t_R FILLER_175_645 ();
 FILLER_ASAP7_75t_R FILLER_175_651 ();
 DECAPx4_ASAP7_75t_R FILLER_175_660 ();
 DECAPx2_ASAP7_75t_R FILLER_175_683 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_689 ();
 DECAPx6_ASAP7_75t_R FILLER_175_700 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_714 ();
 FILLER_ASAP7_75t_R FILLER_175_723 ();
 FILLER_ASAP7_75t_R FILLER_175_733 ();
 DECAPx1_ASAP7_75t_R FILLER_175_738 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_748 ();
 FILLER_ASAP7_75t_R FILLER_175_757 ();
 DECAPx1_ASAP7_75t_R FILLER_175_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_769 ();
 FILLER_ASAP7_75t_R FILLER_175_776 ();
 DECAPx1_ASAP7_75t_R FILLER_175_788 ();
 FILLER_ASAP7_75t_R FILLER_175_798 ();
 FILLER_ASAP7_75t_R FILLER_175_808 ();
 DECAPx1_ASAP7_75t_R FILLER_175_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_822 ();
 DECAPx6_ASAP7_75t_R FILLER_175_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_843 ();
 FILLER_ASAP7_75t_R FILLER_175_853 ();
 DECAPx2_ASAP7_75t_R FILLER_175_858 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_864 ();
 DECAPx1_ASAP7_75t_R FILLER_175_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_879 ();
 DECAPx1_ASAP7_75t_R FILLER_175_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_894 ();
 DECAPx4_ASAP7_75t_R FILLER_175_903 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_913 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_922 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_927 ();
 DECAPx2_ASAP7_75t_R FILLER_175_936 ();
 FILLER_ASAP7_75t_R FILLER_175_948 ();
 DECAPx2_ASAP7_75t_R FILLER_175_958 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_964 ();
 FILLER_ASAP7_75t_R FILLER_175_981 ();
 FILLER_ASAP7_75t_R FILLER_175_993 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1010 ();
 FILLER_ASAP7_75t_R FILLER_175_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1044 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1061 ();
 FILLER_ASAP7_75t_R FILLER_175_1067 ();
 DECAPx4_ASAP7_75t_R FILLER_175_1075 ();
 FILLER_ASAP7_75t_R FILLER_175_1085 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1093 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_1107 ();
 FILLER_ASAP7_75t_R FILLER_175_1117 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1139 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1161 ();
 FILLER_ASAP7_75t_R FILLER_175_1175 ();
 DECAPx6_ASAP7_75t_R FILLER_175_1203 ();
 DECAPx1_ASAP7_75t_R FILLER_175_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_1221 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1248 ();
 FILLER_ASAP7_75t_R FILLER_175_1261 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1269 ();
 FILLER_ASAP7_75t_R FILLER_175_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_175_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_175_1369 ();
 FILLER_ASAP7_75t_R FILLER_175_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_176_2 ();
 DECAPx1_ASAP7_75t_R FILLER_176_24 ();
 FILLER_ASAP7_75t_R FILLER_176_54 ();
 DECAPx10_ASAP7_75t_R FILLER_176_62 ();
 DECAPx10_ASAP7_75t_R FILLER_176_84 ();
 DECAPx6_ASAP7_75t_R FILLER_176_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_120 ();
 DECAPx1_ASAP7_75t_R FILLER_176_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_131 ();
 DECAPx1_ASAP7_75t_R FILLER_176_138 ();
 FILLER_ASAP7_75t_R FILLER_176_148 ();
 DECAPx6_ASAP7_75t_R FILLER_176_153 ();
 DECAPx1_ASAP7_75t_R FILLER_176_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_197 ();
 FILLER_ASAP7_75t_R FILLER_176_206 ();
 DECAPx6_ASAP7_75t_R FILLER_176_214 ();
 DECAPx2_ASAP7_75t_R FILLER_176_234 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_240 ();
 DECAPx1_ASAP7_75t_R FILLER_176_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_253 ();
 DECAPx6_ASAP7_75t_R FILLER_176_257 ();
 DECAPx2_ASAP7_75t_R FILLER_176_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_277 ();
 DECAPx1_ASAP7_75t_R FILLER_176_281 ();
 DECAPx4_ASAP7_75t_R FILLER_176_288 ();
 FILLER_ASAP7_75t_R FILLER_176_298 ();
 DECAPx4_ASAP7_75t_R FILLER_176_326 ();
 FILLER_ASAP7_75t_R FILLER_176_344 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_352 ();
 DECAPx1_ASAP7_75t_R FILLER_176_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_365 ();
 FILLER_ASAP7_75t_R FILLER_176_369 ();
 DECAPx6_ASAP7_75t_R FILLER_176_397 ();
 FILLER_ASAP7_75t_R FILLER_176_411 ();
 DECAPx1_ASAP7_75t_R FILLER_176_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_423 ();
 DECAPx6_ASAP7_75t_R FILLER_176_427 ();
 FILLER_ASAP7_75t_R FILLER_176_447 ();
 DECAPx4_ASAP7_75t_R FILLER_176_452 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_464 ();
 FILLER_ASAP7_75t_R FILLER_176_473 ();
 DECAPx4_ASAP7_75t_R FILLER_176_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_488 ();
 DECAPx10_ASAP7_75t_R FILLER_176_497 ();
 DECAPx2_ASAP7_75t_R FILLER_176_519 ();
 DECAPx1_ASAP7_75t_R FILLER_176_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_539 ();
 DECAPx1_ASAP7_75t_R FILLER_176_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_570 ();
 FILLER_ASAP7_75t_R FILLER_176_577 ();
 DECAPx1_ASAP7_75t_R FILLER_176_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_591 ();
 DECAPx6_ASAP7_75t_R FILLER_176_598 ();
 FILLER_ASAP7_75t_R FILLER_176_612 ();
 DECAPx4_ASAP7_75t_R FILLER_176_620 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_630 ();
 FILLER_ASAP7_75t_R FILLER_176_639 ();
 DECAPx4_ASAP7_75t_R FILLER_176_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_658 ();
 DECAPx2_ASAP7_75t_R FILLER_176_665 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_671 ();
 FILLER_ASAP7_75t_R FILLER_176_700 ();
 FILLER_ASAP7_75t_R FILLER_176_709 ();
 DECAPx10_ASAP7_75t_R FILLER_176_714 ();
 DECAPx10_ASAP7_75t_R FILLER_176_736 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_758 ();
 DECAPx2_ASAP7_75t_R FILLER_176_767 ();
 DECAPx10_ASAP7_75t_R FILLER_176_787 ();
 DECAPx2_ASAP7_75t_R FILLER_176_809 ();
 FILLER_ASAP7_75t_R FILLER_176_815 ();
 DECAPx6_ASAP7_75t_R FILLER_176_820 ();
 DECAPx1_ASAP7_75t_R FILLER_176_834 ();
 FILLER_ASAP7_75t_R FILLER_176_846 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_851 ();
 FILLER_ASAP7_75t_R FILLER_176_860 ();
 DECAPx2_ASAP7_75t_R FILLER_176_888 ();
 DECAPx2_ASAP7_75t_R FILLER_176_900 ();
 FILLER_ASAP7_75t_R FILLER_176_906 ();
 DECAPx1_ASAP7_75t_R FILLER_176_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_918 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_927 ();
 DECAPx10_ASAP7_75t_R FILLER_176_938 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_960 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_1001 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_1007 ();
 DECAPx4_ASAP7_75t_R FILLER_176_1017 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_1027 ();
 FILLER_ASAP7_75t_R FILLER_176_1036 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1078 ();
 FILLER_ASAP7_75t_R FILLER_176_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_176_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1120 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_1126 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1139 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_1145 ();
 DECAPx6_ASAP7_75t_R FILLER_176_1174 ();
 DECAPx1_ASAP7_75t_R FILLER_176_1188 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1195 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_1201 ();
 FILLER_ASAP7_75t_R FILLER_176_1210 ();
 DECAPx6_ASAP7_75t_R FILLER_176_1215 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1229 ();
 FILLER_ASAP7_75t_R FILLER_176_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_176_1246 ();
 DECAPx6_ASAP7_75t_R FILLER_176_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_176_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_176_1361 ();
 FILLER_ASAP7_75t_R FILLER_176_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_177_2 ();
 DECAPx1_ASAP7_75t_R FILLER_177_16 ();
 DECAPx1_ASAP7_75t_R FILLER_177_26 ();
 DECAPx10_ASAP7_75t_R FILLER_177_36 ();
 DECAPx6_ASAP7_75t_R FILLER_177_58 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_177_78 ();
 DECAPx1_ASAP7_75t_R FILLER_177_84 ();
 FILLER_ASAP7_75t_R FILLER_177_96 ();
 DECAPx4_ASAP7_75t_R FILLER_177_104 ();
 FILLER_ASAP7_75t_R FILLER_177_114 ();
 DECAPx4_ASAP7_75t_R FILLER_177_142 ();
 FILLER_ASAP7_75t_R FILLER_177_152 ();
 DECAPx4_ASAP7_75t_R FILLER_177_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_172 ();
 FILLER_ASAP7_75t_R FILLER_177_179 ();
 DECAPx6_ASAP7_75t_R FILLER_177_184 ();
 DECAPx6_ASAP7_75t_R FILLER_177_204 ();
 FILLER_ASAP7_75t_R FILLER_177_218 ();
 DECAPx10_ASAP7_75t_R FILLER_177_226 ();
 DECAPx6_ASAP7_75t_R FILLER_177_248 ();
 FILLER_ASAP7_75t_R FILLER_177_262 ();
 DECAPx4_ASAP7_75t_R FILLER_177_270 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_177_280 ();
 FILLER_ASAP7_75t_R FILLER_177_289 ();
 DECAPx4_ASAP7_75t_R FILLER_177_297 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_177_307 ();
 FILLER_ASAP7_75t_R FILLER_177_316 ();
 FILLER_ASAP7_75t_R FILLER_177_321 ();
 DECAPx4_ASAP7_75t_R FILLER_177_326 ();
 FILLER_ASAP7_75t_R FILLER_177_336 ();
 DECAPx10_ASAP7_75t_R FILLER_177_346 ();
 DECAPx2_ASAP7_75t_R FILLER_177_368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_177_374 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_177_383 ();
 DECAPx2_ASAP7_75t_R FILLER_177_389 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_177_403 ();
 FILLER_ASAP7_75t_R FILLER_177_414 ();
 FILLER_ASAP7_75t_R FILLER_177_422 ();
 DECAPx10_ASAP7_75t_R FILLER_177_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_452 ();
 DECAPx4_ASAP7_75t_R FILLER_177_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_487 ();
 FILLER_ASAP7_75t_R FILLER_177_496 ();
 FILLER_ASAP7_75t_R FILLER_177_520 ();
 FILLER_ASAP7_75t_R FILLER_177_525 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_177_537 ();
 FILLER_ASAP7_75t_R FILLER_177_546 ();
 DECAPx1_ASAP7_75t_R FILLER_177_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_578 ();
 DECAPx2_ASAP7_75t_R FILLER_177_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_593 ();
 FILLER_ASAP7_75t_R FILLER_177_602 ();
 DECAPx2_ASAP7_75t_R FILLER_177_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_616 ();
 DECAPx10_ASAP7_75t_R FILLER_177_624 ();
 DECAPx1_ASAP7_75t_R FILLER_177_646 ();
 DECAPx2_ASAP7_75t_R FILLER_177_660 ();
 FILLER_ASAP7_75t_R FILLER_177_666 ();
 DECAPx1_ASAP7_75t_R FILLER_177_674 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_177_686 ();
 DECAPx4_ASAP7_75t_R FILLER_177_692 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_177_710 ();
 FILLER_ASAP7_75t_R FILLER_177_719 ();
 DECAPx1_ASAP7_75t_R FILLER_177_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_731 ();
 DECAPx2_ASAP7_75t_R FILLER_177_742 ();
 FILLER_ASAP7_75t_R FILLER_177_748 ();
 FILLER_ASAP7_75t_R FILLER_177_764 ();
 DECAPx2_ASAP7_75t_R FILLER_177_773 ();
 FILLER_ASAP7_75t_R FILLER_177_779 ();
 DECAPx4_ASAP7_75t_R FILLER_177_791 ();
 DECAPx1_ASAP7_75t_R FILLER_177_804 ();
 DECAPx6_ASAP7_75t_R FILLER_177_814 ();
 DECAPx1_ASAP7_75t_R FILLER_177_828 ();
 DECAPx4_ASAP7_75t_R FILLER_177_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_868 ();
 FILLER_ASAP7_75t_R FILLER_177_877 ();
 DECAPx10_ASAP7_75t_R FILLER_177_882 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_177_904 ();
 DECAPx4_ASAP7_75t_R FILLER_177_915 ();
 DECAPx1_ASAP7_75t_R FILLER_177_927 ();
 DECAPx4_ASAP7_75t_R FILLER_177_939 ();
 FILLER_ASAP7_75t_R FILLER_177_949 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_177_965 ();
 DECAPx4_ASAP7_75t_R FILLER_177_978 ();
 FILLER_ASAP7_75t_R FILLER_177_988 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1038 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_177_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1054 ();
 FILLER_ASAP7_75t_R FILLER_177_1060 ();
 FILLER_ASAP7_75t_R FILLER_177_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1076 ();
 DECAPx4_ASAP7_75t_R FILLER_177_1098 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1128 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_177_1137 ();
 FILLER_ASAP7_75t_R FILLER_177_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_177_1176 ();
 DECAPx4_ASAP7_75t_R FILLER_177_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1243 ();
 FILLER_ASAP7_75t_R FILLER_177_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_177_1336 ();
 DECAPx6_ASAP7_75t_R FILLER_177_1358 ();
 DECAPx1_ASAP7_75t_R FILLER_177_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_178_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_8 ();
 DECAPx4_ASAP7_75t_R FILLER_178_37 ();
 FILLER_ASAP7_75t_R FILLER_178_47 ();
 DECAPx2_ASAP7_75t_R FILLER_178_55 ();
 FILLER_ASAP7_75t_R FILLER_178_61 ();
 FILLER_ASAP7_75t_R FILLER_178_71 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_81 ();
 FILLER_ASAP7_75t_R FILLER_178_90 ();
 DECAPx2_ASAP7_75t_R FILLER_178_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_104 ();
 DECAPx1_ASAP7_75t_R FILLER_178_111 ();
 DECAPx4_ASAP7_75t_R FILLER_178_118 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_128 ();
 DECAPx6_ASAP7_75t_R FILLER_178_134 ();
 DECAPx2_ASAP7_75t_R FILLER_178_148 ();
 DECAPx10_ASAP7_75t_R FILLER_178_162 ();
 DECAPx10_ASAP7_75t_R FILLER_178_184 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_206 ();
 DECAPx2_ASAP7_75t_R FILLER_178_235 ();
 DECAPx2_ASAP7_75t_R FILLER_178_247 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_253 ();
 DECAPx1_ASAP7_75t_R FILLER_178_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_286 ();
 DECAPx10_ASAP7_75t_R FILLER_178_295 ();
 DECAPx4_ASAP7_75t_R FILLER_178_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_327 ();
 DECAPx1_ASAP7_75t_R FILLER_178_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_340 ();
 DECAPx2_ASAP7_75t_R FILLER_178_347 ();
 FILLER_ASAP7_75t_R FILLER_178_353 ();
 DECAPx2_ASAP7_75t_R FILLER_178_361 ();
 FILLER_ASAP7_75t_R FILLER_178_367 ();
 DECAPx10_ASAP7_75t_R FILLER_178_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_397 ();
 DECAPx2_ASAP7_75t_R FILLER_178_407 ();
 DECAPx2_ASAP7_75t_R FILLER_178_421 ();
 DECAPx1_ASAP7_75t_R FILLER_178_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_438 ();
 DECAPx4_ASAP7_75t_R FILLER_178_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_461 ();
 FILLER_ASAP7_75t_R FILLER_178_464 ();
 FILLER_ASAP7_75t_R FILLER_178_472 ();
 DECAPx1_ASAP7_75t_R FILLER_178_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_481 ();
 DECAPx2_ASAP7_75t_R FILLER_178_485 ();
 DECAPx1_ASAP7_75t_R FILLER_178_497 ();
 FILLER_ASAP7_75t_R FILLER_178_527 ();
 DECAPx6_ASAP7_75t_R FILLER_178_535 ();
 DECAPx1_ASAP7_75t_R FILLER_178_549 ();
 DECAPx1_ASAP7_75t_R FILLER_178_559 ();
 DECAPx10_ASAP7_75t_R FILLER_178_566 ();
 DECAPx2_ASAP7_75t_R FILLER_178_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_594 ();
 DECAPx2_ASAP7_75t_R FILLER_178_603 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_609 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_622 ();
 DECAPx4_ASAP7_75t_R FILLER_178_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_645 ();
 DECAPx1_ASAP7_75t_R FILLER_178_654 ();
 DECAPx1_ASAP7_75t_R FILLER_178_670 ();
 DECAPx10_ASAP7_75t_R FILLER_178_682 ();
 FILLER_ASAP7_75t_R FILLER_178_704 ();
 FILLER_ASAP7_75t_R FILLER_178_709 ();
 FILLER_ASAP7_75t_R FILLER_178_718 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_728 ();
 FILLER_ASAP7_75t_R FILLER_178_757 ();
 FILLER_ASAP7_75t_R FILLER_178_773 ();
 DECAPx4_ASAP7_75t_R FILLER_178_785 ();
 FILLER_ASAP7_75t_R FILLER_178_795 ();
 DECAPx1_ASAP7_75t_R FILLER_178_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_807 ();
 FILLER_ASAP7_75t_R FILLER_178_834 ();
 DECAPx10_ASAP7_75t_R FILLER_178_846 ();
 FILLER_ASAP7_75t_R FILLER_178_868 ();
 DECAPx4_ASAP7_75t_R FILLER_178_874 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_884 ();
 DECAPx1_ASAP7_75t_R FILLER_178_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_897 ();
 DECAPx2_ASAP7_75t_R FILLER_178_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_930 ();
 DECAPx10_ASAP7_75t_R FILLER_178_937 ();
 DECAPx2_ASAP7_75t_R FILLER_178_959 ();
 FILLER_ASAP7_75t_R FILLER_178_965 ();
 DECAPx2_ASAP7_75t_R FILLER_178_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_985 ();
 FILLER_ASAP7_75t_R FILLER_178_993 ();
 FILLER_ASAP7_75t_R FILLER_178_1001 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_1009 ();
 FILLER_ASAP7_75t_R FILLER_178_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1028 ();
 FILLER_ASAP7_75t_R FILLER_178_1034 ();
 FILLER_ASAP7_75t_R FILLER_178_1043 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_1048 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1072 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_178_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1098 ();
 DECAPx1_ASAP7_75t_R FILLER_178_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1117 ();
 DECAPx4_ASAP7_75t_R FILLER_178_1139 ();
 DECAPx1_ASAP7_75t_R FILLER_178_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1161 ();
 FILLER_ASAP7_75t_R FILLER_178_1165 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1193 ();
 FILLER_ASAP7_75t_R FILLER_178_1207 ();
 DECAPx6_ASAP7_75t_R FILLER_178_1212 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_178_1349 ();
 DECAPx2_ASAP7_75t_R FILLER_178_1371 ();
 DECAPx6_ASAP7_75t_R FILLER_179_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_16 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_23 ();
 DECAPx1_ASAP7_75t_R FILLER_179_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_33 ();
 DECAPx2_ASAP7_75t_R FILLER_179_60 ();
 DECAPx4_ASAP7_75t_R FILLER_179_72 ();
 FILLER_ASAP7_75t_R FILLER_179_85 ();
 DECAPx1_ASAP7_75t_R FILLER_179_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_99 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_126 ();
 DECAPx2_ASAP7_75t_R FILLER_179_135 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_141 ();
 DECAPx2_ASAP7_75t_R FILLER_179_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_153 ();
 FILLER_ASAP7_75t_R FILLER_179_160 ();
 DECAPx10_ASAP7_75t_R FILLER_179_168 ();
 DECAPx2_ASAP7_75t_R FILLER_179_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_196 ();
 DECAPx4_ASAP7_75t_R FILLER_179_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_213 ();
 DECAPx1_ASAP7_75t_R FILLER_179_220 ();
 DECAPx2_ASAP7_75t_R FILLER_179_227 ();
 FILLER_ASAP7_75t_R FILLER_179_259 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_267 ();
 DECAPx4_ASAP7_75t_R FILLER_179_273 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_283 ();
 FILLER_ASAP7_75t_R FILLER_179_294 ();
 DECAPx2_ASAP7_75t_R FILLER_179_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_308 ();
 DECAPx2_ASAP7_75t_R FILLER_179_315 ();
 FILLER_ASAP7_75t_R FILLER_179_327 ();
 DECAPx2_ASAP7_75t_R FILLER_179_337 ();
 FILLER_ASAP7_75t_R FILLER_179_343 ();
 FILLER_ASAP7_75t_R FILLER_179_351 ();
 DECAPx6_ASAP7_75t_R FILLER_179_359 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_379 ();
 DECAPx10_ASAP7_75t_R FILLER_179_388 ();
 DECAPx2_ASAP7_75t_R FILLER_179_410 ();
 FILLER_ASAP7_75t_R FILLER_179_416 ();
 DECAPx2_ASAP7_75t_R FILLER_179_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_432 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_443 ();
 FILLER_ASAP7_75t_R FILLER_179_453 ();
 DECAPx2_ASAP7_75t_R FILLER_179_481 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_487 ();
 DECAPx2_ASAP7_75t_R FILLER_179_496 ();
 FILLER_ASAP7_75t_R FILLER_179_508 ();
 DECAPx1_ASAP7_75t_R FILLER_179_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_520 ();
 FILLER_ASAP7_75t_R FILLER_179_527 ();
 DECAPx6_ASAP7_75t_R FILLER_179_535 ();
 DECAPx1_ASAP7_75t_R FILLER_179_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_553 ();
 DECAPx10_ASAP7_75t_R FILLER_179_557 ();
 DECAPx10_ASAP7_75t_R FILLER_179_579 ();
 DECAPx6_ASAP7_75t_R FILLER_179_601 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_615 ();
 FILLER_ASAP7_75t_R FILLER_179_632 ();
 DECAPx1_ASAP7_75t_R FILLER_179_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_646 ();
 DECAPx2_ASAP7_75t_R FILLER_179_655 ();
 FILLER_ASAP7_75t_R FILLER_179_664 ();
 DECAPx1_ASAP7_75t_R FILLER_179_684 ();
 DECAPx6_ASAP7_75t_R FILLER_179_714 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_728 ();
 DECAPx2_ASAP7_75t_R FILLER_179_737 ();
 FILLER_ASAP7_75t_R FILLER_179_743 ();
 DECAPx6_ASAP7_75t_R FILLER_179_748 ();
 DECAPx2_ASAP7_75t_R FILLER_179_762 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_774 ();
 DECAPx1_ASAP7_75t_R FILLER_179_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_788 ();
 FILLER_ASAP7_75t_R FILLER_179_795 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_805 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_814 ();
 FILLER_ASAP7_75t_R FILLER_179_820 ();
 DECAPx2_ASAP7_75t_R FILLER_179_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_842 ();
 DECAPx10_ASAP7_75t_R FILLER_179_851 ();
 DECAPx10_ASAP7_75t_R FILLER_179_873 ();
 DECAPx2_ASAP7_75t_R FILLER_179_905 ();
 FILLER_ASAP7_75t_R FILLER_179_911 ();
 DECAPx2_ASAP7_75t_R FILLER_179_916 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_922 ();
 FILLER_ASAP7_75t_R FILLER_179_927 ();
 DECAPx4_ASAP7_75t_R FILLER_179_937 ();
 DECAPx2_ASAP7_75t_R FILLER_179_954 ();
 FILLER_ASAP7_75t_R FILLER_179_960 ();
 FILLER_ASAP7_75t_R FILLER_179_965 ();
 FILLER_ASAP7_75t_R FILLER_179_981 ();
 FILLER_ASAP7_75t_R FILLER_179_993 ();
 FILLER_ASAP7_75t_R FILLER_179_1003 ();
 FILLER_ASAP7_75t_R FILLER_179_1011 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_1020 ();
 FILLER_ASAP7_75t_R FILLER_179_1031 ();
 FILLER_ASAP7_75t_R FILLER_179_1043 ();
 FILLER_ASAP7_75t_R FILLER_179_1052 ();
 FILLER_ASAP7_75t_R FILLER_179_1062 ();
 DECAPx1_ASAP7_75t_R FILLER_179_1070 ();
 FILLER_ASAP7_75t_R FILLER_179_1082 ();
 FILLER_ASAP7_75t_R FILLER_179_1091 ();
 FILLER_ASAP7_75t_R FILLER_179_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_179_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1120 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_179_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1143 ();
 FILLER_ASAP7_75t_R FILLER_179_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_179_1157 ();
 FILLER_ASAP7_75t_R FILLER_179_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_179_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_179_1337 ();
 DECAPx6_ASAP7_75t_R FILLER_179_1359 ();
 DECAPx1_ASAP7_75t_R FILLER_179_1373 ();
 DECAPx10_ASAP7_75t_R FILLER_180_2 ();
 FILLER_ASAP7_75t_R FILLER_180_24 ();
 DECAPx4_ASAP7_75t_R FILLER_180_32 ();
 FILLER_ASAP7_75t_R FILLER_180_48 ();
 DECAPx2_ASAP7_75t_R FILLER_180_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_59 ();
 DECAPx10_ASAP7_75t_R FILLER_180_63 ();
 DECAPx6_ASAP7_75t_R FILLER_180_85 ();
 DECAPx1_ASAP7_75t_R FILLER_180_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_103 ();
 DECAPx2_ASAP7_75t_R FILLER_180_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_116 ();
 DECAPx2_ASAP7_75t_R FILLER_180_143 ();
 FILLER_ASAP7_75t_R FILLER_180_149 ();
 DECAPx4_ASAP7_75t_R FILLER_180_157 ();
 FILLER_ASAP7_75t_R FILLER_180_173 ();
 FILLER_ASAP7_75t_R FILLER_180_181 ();
 DECAPx4_ASAP7_75t_R FILLER_180_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_219 ();
 DECAPx4_ASAP7_75t_R FILLER_180_226 ();
 DECAPx1_ASAP7_75t_R FILLER_180_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_246 ();
 DECAPx6_ASAP7_75t_R FILLER_180_250 ();
 DECAPx10_ASAP7_75t_R FILLER_180_270 ();
 DECAPx2_ASAP7_75t_R FILLER_180_292 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_180_298 ();
 FILLER_ASAP7_75t_R FILLER_180_327 ();
 DECAPx6_ASAP7_75t_R FILLER_180_335 ();
 DECAPx2_ASAP7_75t_R FILLER_180_349 ();
 DECAPx2_ASAP7_75t_R FILLER_180_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_370 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_180_379 ();
 FILLER_ASAP7_75t_R FILLER_180_390 ();
 FILLER_ASAP7_75t_R FILLER_180_398 ();
 DECAPx4_ASAP7_75t_R FILLER_180_409 ();
 FILLER_ASAP7_75t_R FILLER_180_419 ();
 DECAPx2_ASAP7_75t_R FILLER_180_431 ();
 FILLER_ASAP7_75t_R FILLER_180_443 ();
 DECAPx4_ASAP7_75t_R FILLER_180_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_461 ();
 FILLER_ASAP7_75t_R FILLER_180_464 ();
 DECAPx2_ASAP7_75t_R FILLER_180_472 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_180_478 ();
 FILLER_ASAP7_75t_R FILLER_180_487 ();
 DECAPx10_ASAP7_75t_R FILLER_180_495 ();
 DECAPx2_ASAP7_75t_R FILLER_180_539 ();
 DECAPx2_ASAP7_75t_R FILLER_180_551 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_180_557 ();
 DECAPx1_ASAP7_75t_R FILLER_180_563 ();
 FILLER_ASAP7_75t_R FILLER_180_573 ();
 FILLER_ASAP7_75t_R FILLER_180_578 ();
 DECAPx2_ASAP7_75t_R FILLER_180_588 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_180_594 ();
 FILLER_ASAP7_75t_R FILLER_180_603 ();
 FILLER_ASAP7_75t_R FILLER_180_611 ();
 DECAPx2_ASAP7_75t_R FILLER_180_616 ();
 FILLER_ASAP7_75t_R FILLER_180_622 ();
 FILLER_ASAP7_75t_R FILLER_180_634 ();
 DECAPx4_ASAP7_75t_R FILLER_180_643 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_180_653 ();
 DECAPx4_ASAP7_75t_R FILLER_180_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_670 ();
 FILLER_ASAP7_75t_R FILLER_180_677 ();
 DECAPx2_ASAP7_75t_R FILLER_180_683 ();
 DECAPx1_ASAP7_75t_R FILLER_180_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_701 ();
 DECAPx10_ASAP7_75t_R FILLER_180_705 ();
 FILLER_ASAP7_75t_R FILLER_180_727 ();
 DECAPx10_ASAP7_75t_R FILLER_180_735 ();
 DECAPx4_ASAP7_75t_R FILLER_180_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_770 ();
 DECAPx1_ASAP7_75t_R FILLER_180_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_779 ();
 FILLER_ASAP7_75t_R FILLER_180_790 ();
 DECAPx6_ASAP7_75t_R FILLER_180_798 ();
 DECAPx2_ASAP7_75t_R FILLER_180_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_818 ();
 DECAPx6_ASAP7_75t_R FILLER_180_827 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_180_841 ();
 FILLER_ASAP7_75t_R FILLER_180_870 ();
 FILLER_ASAP7_75t_R FILLER_180_880 ();
 DECAPx2_ASAP7_75t_R FILLER_180_888 ();
 DECAPx1_ASAP7_75t_R FILLER_180_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_905 ();
 DECAPx1_ASAP7_75t_R FILLER_180_912 ();
 FILLER_ASAP7_75t_R FILLER_180_922 ();
 FILLER_ASAP7_75t_R FILLER_180_950 ();
 FILLER_ASAP7_75t_R FILLER_180_978 ();
 FILLER_ASAP7_75t_R FILLER_180_990 ();
 DECAPx6_ASAP7_75t_R FILLER_180_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_180_1020 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_180_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_180_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_180_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_180_1058 ();
 DECAPx6_ASAP7_75t_R FILLER_180_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_180_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_180_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1103 ();
 FILLER_ASAP7_75t_R FILLER_180_1110 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1119 ();
 DECAPx4_ASAP7_75t_R FILLER_180_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_180_1346 ();
 DECAPx2_ASAP7_75t_R FILLER_180_1368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_180_1374 ();
 DECAPx6_ASAP7_75t_R FILLER_181_2 ();
 DECAPx1_ASAP7_75t_R FILLER_181_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_20 ();
 DECAPx4_ASAP7_75t_R FILLER_181_47 ();
 FILLER_ASAP7_75t_R FILLER_181_57 ();
 FILLER_ASAP7_75t_R FILLER_181_65 ();
 DECAPx6_ASAP7_75t_R FILLER_181_73 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_87 ();
 FILLER_ASAP7_75t_R FILLER_181_96 ();
 DECAPx6_ASAP7_75t_R FILLER_181_104 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_118 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_127 ();
 FILLER_ASAP7_75t_R FILLER_181_133 ();
 DECAPx2_ASAP7_75t_R FILLER_181_161 ();
 FILLER_ASAP7_75t_R FILLER_181_193 ();
 FILLER_ASAP7_75t_R FILLER_181_201 ();
 DECAPx1_ASAP7_75t_R FILLER_181_206 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_236 ();
 DECAPx2_ASAP7_75t_R FILLER_181_245 ();
 FILLER_ASAP7_75t_R FILLER_181_251 ();
 DECAPx6_ASAP7_75t_R FILLER_181_279 ();
 DECAPx1_ASAP7_75t_R FILLER_181_293 ();
 FILLER_ASAP7_75t_R FILLER_181_303 ();
 DECAPx1_ASAP7_75t_R FILLER_181_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_315 ();
 DECAPx10_ASAP7_75t_R FILLER_181_319 ();
 DECAPx4_ASAP7_75t_R FILLER_181_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_351 ();
 DECAPx4_ASAP7_75t_R FILLER_181_358 ();
 FILLER_ASAP7_75t_R FILLER_181_371 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_395 ();
 DECAPx2_ASAP7_75t_R FILLER_181_408 ();
 FILLER_ASAP7_75t_R FILLER_181_424 ();
 DECAPx2_ASAP7_75t_R FILLER_181_432 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_438 ();
 DECAPx2_ASAP7_75t_R FILLER_181_467 ();
 FILLER_ASAP7_75t_R FILLER_181_473 ();
 DECAPx2_ASAP7_75t_R FILLER_181_501 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_507 ();
 DECAPx2_ASAP7_75t_R FILLER_181_516 ();
 FILLER_ASAP7_75t_R FILLER_181_528 ();
 FILLER_ASAP7_75t_R FILLER_181_556 ();
 FILLER_ASAP7_75t_R FILLER_181_584 ();
 DECAPx1_ASAP7_75t_R FILLER_181_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_598 ();
 DECAPx2_ASAP7_75t_R FILLER_181_625 ();
 DECAPx10_ASAP7_75t_R FILLER_181_639 ();
 DECAPx2_ASAP7_75t_R FILLER_181_661 ();
 FILLER_ASAP7_75t_R FILLER_181_676 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_685 ();
 DECAPx4_ASAP7_75t_R FILLER_181_694 ();
 FILLER_ASAP7_75t_R FILLER_181_704 ();
 DECAPx10_ASAP7_75t_R FILLER_181_709 ();
 FILLER_ASAP7_75t_R FILLER_181_731 ();
 FILLER_ASAP7_75t_R FILLER_181_740 ();
 DECAPx10_ASAP7_75t_R FILLER_181_768 ();
 DECAPx4_ASAP7_75t_R FILLER_181_790 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_800 ();
 DECAPx10_ASAP7_75t_R FILLER_181_809 ();
 DECAPx2_ASAP7_75t_R FILLER_181_831 ();
 DECAPx2_ASAP7_75t_R FILLER_181_840 ();
 FILLER_ASAP7_75t_R FILLER_181_846 ();
 DECAPx1_ASAP7_75t_R FILLER_181_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_858 ();
 FILLER_ASAP7_75t_R FILLER_181_862 ();
 DECAPx2_ASAP7_75t_R FILLER_181_867 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_873 ();
 FILLER_ASAP7_75t_R FILLER_181_884 ();
 DECAPx4_ASAP7_75t_R FILLER_181_894 ();
 FILLER_ASAP7_75t_R FILLER_181_904 ();
 DECAPx4_ASAP7_75t_R FILLER_181_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_924 ();
 DECAPx1_ASAP7_75t_R FILLER_181_927 ();
 FILLER_ASAP7_75t_R FILLER_181_939 ();
 DECAPx1_ASAP7_75t_R FILLER_181_944 ();
 DECAPx10_ASAP7_75t_R FILLER_181_954 ();
 DECAPx10_ASAP7_75t_R FILLER_181_976 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1026 ();
 DECAPx6_ASAP7_75t_R FILLER_181_1048 ();
 FILLER_ASAP7_75t_R FILLER_181_1062 ();
 DECAPx6_ASAP7_75t_R FILLER_181_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_181_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1090 ();
 DECAPx6_ASAP7_75t_R FILLER_181_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_1112 ();
 DECAPx4_ASAP7_75t_R FILLER_181_1119 ();
 DECAPx4_ASAP7_75t_R FILLER_181_1137 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1158 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1208 ();
 FILLER_ASAP7_75t_R FILLER_181_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_181_1349 ();
 DECAPx2_ASAP7_75t_R FILLER_181_1371 ();
 DECAPx6_ASAP7_75t_R FILLER_182_2 ();
 DECAPx1_ASAP7_75t_R FILLER_182_16 ();
 DECAPx1_ASAP7_75t_R FILLER_182_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_30 ();
 FILLER_ASAP7_75t_R FILLER_182_37 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_42 ();
 DECAPx1_ASAP7_75t_R FILLER_182_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_55 ();
 FILLER_ASAP7_75t_R FILLER_182_82 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_110 ();
 DECAPx2_ASAP7_75t_R FILLER_182_119 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_125 ();
 DECAPx1_ASAP7_75t_R FILLER_182_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_138 ();
 DECAPx1_ASAP7_75t_R FILLER_182_145 ();
 DECAPx4_ASAP7_75t_R FILLER_182_152 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_162 ();
 DECAPx4_ASAP7_75t_R FILLER_182_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_181 ();
 DECAPx6_ASAP7_75t_R FILLER_182_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_199 ();
 DECAPx2_ASAP7_75t_R FILLER_182_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_212 ();
 DECAPx2_ASAP7_75t_R FILLER_182_219 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_228 ();
 FILLER_ASAP7_75t_R FILLER_182_234 ();
 FILLER_ASAP7_75t_R FILLER_182_244 ();
 DECAPx2_ASAP7_75t_R FILLER_182_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_258 ();
 FILLER_ASAP7_75t_R FILLER_182_265 ();
 DECAPx2_ASAP7_75t_R FILLER_182_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_276 ();
 DECAPx6_ASAP7_75t_R FILLER_182_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_294 ();
 DECAPx10_ASAP7_75t_R FILLER_182_301 ();
 DECAPx6_ASAP7_75t_R FILLER_182_323 ();
 DECAPx1_ASAP7_75t_R FILLER_182_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_341 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_368 ();
 DECAPx6_ASAP7_75t_R FILLER_182_377 ();
 DECAPx1_ASAP7_75t_R FILLER_182_391 ();
 DECAPx10_ASAP7_75t_R FILLER_182_401 ();
 DECAPx10_ASAP7_75t_R FILLER_182_423 ();
 DECAPx4_ASAP7_75t_R FILLER_182_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_461 ();
 DECAPx2_ASAP7_75t_R FILLER_182_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_470 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_477 ();
 DECAPx2_ASAP7_75t_R FILLER_182_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_489 ();
 DECAPx2_ASAP7_75t_R FILLER_182_493 ();
 FILLER_ASAP7_75t_R FILLER_182_499 ();
 DECAPx4_ASAP7_75t_R FILLER_182_527 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_537 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_546 ();
 DECAPx4_ASAP7_75t_R FILLER_182_552 ();
 DECAPx2_ASAP7_75t_R FILLER_182_568 ();
 FILLER_ASAP7_75t_R FILLER_182_580 ();
 DECAPx10_ASAP7_75t_R FILLER_182_588 ();
 FILLER_ASAP7_75t_R FILLER_182_610 ();
 DECAPx4_ASAP7_75t_R FILLER_182_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_625 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_636 ();
 DECAPx1_ASAP7_75t_R FILLER_182_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_651 ();
 DECAPx6_ASAP7_75t_R FILLER_182_664 ();
 DECAPx1_ASAP7_75t_R FILLER_182_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_682 ();
 FILLER_ASAP7_75t_R FILLER_182_689 ();
 FILLER_ASAP7_75t_R FILLER_182_717 ();
 DECAPx1_ASAP7_75t_R FILLER_182_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_726 ();
 FILLER_ASAP7_75t_R FILLER_182_734 ();
 DECAPx6_ASAP7_75t_R FILLER_182_742 ();
 DECAPx4_ASAP7_75t_R FILLER_182_764 ();
 FILLER_ASAP7_75t_R FILLER_182_774 ();
 FILLER_ASAP7_75t_R FILLER_182_782 ();
 DECAPx1_ASAP7_75t_R FILLER_182_793 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_800 ();
 FILLER_ASAP7_75t_R FILLER_182_829 ();
 FILLER_ASAP7_75t_R FILLER_182_837 ();
 FILLER_ASAP7_75t_R FILLER_182_844 ();
 DECAPx2_ASAP7_75t_R FILLER_182_852 ();
 DECAPx6_ASAP7_75t_R FILLER_182_884 ();
 DECAPx2_ASAP7_75t_R FILLER_182_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_904 ();
 DECAPx10_ASAP7_75t_R FILLER_182_913 ();
 DECAPx10_ASAP7_75t_R FILLER_182_935 ();
 DECAPx1_ASAP7_75t_R FILLER_182_957 ();
 DECAPx2_ASAP7_75t_R FILLER_182_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_981 ();
 FILLER_ASAP7_75t_R FILLER_182_992 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1001 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_182_1018 ();
 DECAPx6_ASAP7_75t_R FILLER_182_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_182_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1074 ();
 FILLER_ASAP7_75t_R FILLER_182_1106 ();
 FILLER_ASAP7_75t_R FILLER_182_1114 ();
 DECAPx1_ASAP7_75t_R FILLER_182_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1136 ();
 DECAPx4_ASAP7_75t_R FILLER_182_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_182_1348 ();
 DECAPx2_ASAP7_75t_R FILLER_182_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_183_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_8 ();
 DECAPx2_ASAP7_75t_R FILLER_183_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_41 ();
 FILLER_ASAP7_75t_R FILLER_183_45 ();
 DECAPx6_ASAP7_75t_R FILLER_183_55 ();
 DECAPx1_ASAP7_75t_R FILLER_183_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_73 ();
 DECAPx10_ASAP7_75t_R FILLER_183_77 ();
 DECAPx1_ASAP7_75t_R FILLER_183_102 ();
 DECAPx1_ASAP7_75t_R FILLER_183_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_113 ();
 DECAPx6_ASAP7_75t_R FILLER_183_136 ();
 DECAPx2_ASAP7_75t_R FILLER_183_150 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_183_182 ();
 DECAPx2_ASAP7_75t_R FILLER_183_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_197 ();
 DECAPx6_ASAP7_75t_R FILLER_183_224 ();
 FILLER_ASAP7_75t_R FILLER_183_238 ();
 DECAPx6_ASAP7_75t_R FILLER_183_248 ();
 DECAPx1_ASAP7_75t_R FILLER_183_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_272 ();
 FILLER_ASAP7_75t_R FILLER_183_279 ();
 FILLER_ASAP7_75t_R FILLER_183_289 ();
 DECAPx2_ASAP7_75t_R FILLER_183_299 ();
 FILLER_ASAP7_75t_R FILLER_183_305 ();
 DECAPx2_ASAP7_75t_R FILLER_183_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_319 ();
 FILLER_ASAP7_75t_R FILLER_183_328 ();
 DECAPx2_ASAP7_75t_R FILLER_183_338 ();
 FILLER_ASAP7_75t_R FILLER_183_344 ();
 DECAPx1_ASAP7_75t_R FILLER_183_352 ();
 DECAPx6_ASAP7_75t_R FILLER_183_359 ();
 DECAPx2_ASAP7_75t_R FILLER_183_379 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_183_385 ();
 FILLER_ASAP7_75t_R FILLER_183_394 ();
 DECAPx2_ASAP7_75t_R FILLER_183_402 ();
 DECAPx2_ASAP7_75t_R FILLER_183_414 ();
 FILLER_ASAP7_75t_R FILLER_183_428 ();
 DECAPx2_ASAP7_75t_R FILLER_183_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_442 ();
 DECAPx2_ASAP7_75t_R FILLER_183_449 ();
 DECAPx2_ASAP7_75t_R FILLER_183_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_464 ();
 DECAPx6_ASAP7_75t_R FILLER_183_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_505 ();
 DECAPx1_ASAP7_75t_R FILLER_183_512 ();
 DECAPx1_ASAP7_75t_R FILLER_183_519 ();
 FILLER_ASAP7_75t_R FILLER_183_529 ();
 FILLER_ASAP7_75t_R FILLER_183_537 ();
 DECAPx10_ASAP7_75t_R FILLER_183_542 ();
 DECAPx6_ASAP7_75t_R FILLER_183_564 ();
 DECAPx2_ASAP7_75t_R FILLER_183_578 ();
 DECAPx1_ASAP7_75t_R FILLER_183_590 ();
 FILLER_ASAP7_75t_R FILLER_183_600 ();
 DECAPx6_ASAP7_75t_R FILLER_183_609 ();
 FILLER_ASAP7_75t_R FILLER_183_623 ();
 FILLER_ASAP7_75t_R FILLER_183_637 ();
 DECAPx2_ASAP7_75t_R FILLER_183_646 ();
 FILLER_ASAP7_75t_R FILLER_183_652 ();
 DECAPx6_ASAP7_75t_R FILLER_183_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_680 ();
 DECAPx2_ASAP7_75t_R FILLER_183_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_693 ();
 DECAPx1_ASAP7_75t_R FILLER_183_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_704 ();
 FILLER_ASAP7_75t_R FILLER_183_731 ();
 DECAPx6_ASAP7_75t_R FILLER_183_739 ();
 FILLER_ASAP7_75t_R FILLER_183_753 ();
 FILLER_ASAP7_75t_R FILLER_183_761 ();
 DECAPx1_ASAP7_75t_R FILLER_183_769 ();
 DECAPx6_ASAP7_75t_R FILLER_183_779 ();
 DECAPx1_ASAP7_75t_R FILLER_183_793 ();
 FILLER_ASAP7_75t_R FILLER_183_805 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_183_813 ();
 DECAPx1_ASAP7_75t_R FILLER_183_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_846 ();
 DECAPx6_ASAP7_75t_R FILLER_183_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_868 ();
 FILLER_ASAP7_75t_R FILLER_183_875 ();
 FILLER_ASAP7_75t_R FILLER_183_880 ();
 FILLER_ASAP7_75t_R FILLER_183_890 ();
 DECAPx2_ASAP7_75t_R FILLER_183_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_924 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_183_927 ();
 DECAPx1_ASAP7_75t_R FILLER_183_938 ();
 DECAPx2_ASAP7_75t_R FILLER_183_945 ();
 FILLER_ASAP7_75t_R FILLER_183_951 ();
 DECAPx2_ASAP7_75t_R FILLER_183_959 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_183_991 ();
 DECAPx2_ASAP7_75t_R FILLER_183_1001 ();
 FILLER_ASAP7_75t_R FILLER_183_1007 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_183_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_183_1026 ();
 FILLER_ASAP7_75t_R FILLER_183_1040 ();
 FILLER_ASAP7_75t_R FILLER_183_1048 ();
 DECAPx4_ASAP7_75t_R FILLER_183_1056 ();
 FILLER_ASAP7_75t_R FILLER_183_1066 ();
 FILLER_ASAP7_75t_R FILLER_183_1075 ();
 FILLER_ASAP7_75t_R FILLER_183_1085 ();
 FILLER_ASAP7_75t_R FILLER_183_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1098 ();
 DECAPx1_ASAP7_75t_R FILLER_183_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_183_1349 ();
 DECAPx2_ASAP7_75t_R FILLER_183_1371 ();
 DECAPx4_ASAP7_75t_R FILLER_184_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_12 ();
 DECAPx1_ASAP7_75t_R FILLER_184_19 ();
 DECAPx10_ASAP7_75t_R FILLER_184_26 ();
 DECAPx4_ASAP7_75t_R FILLER_184_56 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_66 ();
 DECAPx10_ASAP7_75t_R FILLER_184_75 ();
 DECAPx4_ASAP7_75t_R FILLER_184_97 ();
 FILLER_ASAP7_75t_R FILLER_184_107 ();
 DECAPx2_ASAP7_75t_R FILLER_184_117 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_123 ();
 FILLER_ASAP7_75t_R FILLER_184_152 ();
 FILLER_ASAP7_75t_R FILLER_184_164 ();
 DECAPx2_ASAP7_75t_R FILLER_184_172 ();
 FILLER_ASAP7_75t_R FILLER_184_184 ();
 DECAPx4_ASAP7_75t_R FILLER_184_194 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_210 ();
 DECAPx2_ASAP7_75t_R FILLER_184_216 ();
 DECAPx10_ASAP7_75t_R FILLER_184_225 ();
 DECAPx1_ASAP7_75t_R FILLER_184_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_251 ();
 FILLER_ASAP7_75t_R FILLER_184_278 ();
 DECAPx1_ASAP7_75t_R FILLER_184_286 ();
 FILLER_ASAP7_75t_R FILLER_184_296 ();
 FILLER_ASAP7_75t_R FILLER_184_324 ();
 FILLER_ASAP7_75t_R FILLER_184_332 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_340 ();
 FILLER_ASAP7_75t_R FILLER_184_349 ();
 FILLER_ASAP7_75t_R FILLER_184_357 ();
 FILLER_ASAP7_75t_R FILLER_184_365 ();
 FILLER_ASAP7_75t_R FILLER_184_375 ();
 DECAPx4_ASAP7_75t_R FILLER_184_385 ();
 DECAPx2_ASAP7_75t_R FILLER_184_401 ();
 DECAPx2_ASAP7_75t_R FILLER_184_413 ();
 FILLER_ASAP7_75t_R FILLER_184_427 ();
 DECAPx2_ASAP7_75t_R FILLER_184_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_461 ();
 FILLER_ASAP7_75t_R FILLER_184_464 ();
 DECAPx4_ASAP7_75t_R FILLER_184_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_482 ();
 DECAPx6_ASAP7_75t_R FILLER_184_489 ();
 DECAPx1_ASAP7_75t_R FILLER_184_503 ();
 FILLER_ASAP7_75t_R FILLER_184_513 ();
 DECAPx2_ASAP7_75t_R FILLER_184_518 ();
 DECAPx2_ASAP7_75t_R FILLER_184_550 ();
 DECAPx2_ASAP7_75t_R FILLER_184_559 ();
 FILLER_ASAP7_75t_R FILLER_184_565 ();
 FILLER_ASAP7_75t_R FILLER_184_570 ();
 DECAPx6_ASAP7_75t_R FILLER_184_580 ();
 DECAPx4_ASAP7_75t_R FILLER_184_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_610 ();
 DECAPx4_ASAP7_75t_R FILLER_184_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_629 ();
 DECAPx6_ASAP7_75t_R FILLER_184_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_650 ();
 DECAPx2_ASAP7_75t_R FILLER_184_663 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_669 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_681 ();
 DECAPx6_ASAP7_75t_R FILLER_184_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_704 ();
 DECAPx10_ASAP7_75t_R FILLER_184_708 ();
 DECAPx4_ASAP7_75t_R FILLER_184_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_740 ();
 DECAPx2_ASAP7_75t_R FILLER_184_751 ();
 FILLER_ASAP7_75t_R FILLER_184_757 ();
 FILLER_ASAP7_75t_R FILLER_184_785 ();
 DECAPx10_ASAP7_75t_R FILLER_184_790 ();
 DECAPx2_ASAP7_75t_R FILLER_184_812 ();
 DECAPx2_ASAP7_75t_R FILLER_184_821 ();
 FILLER_ASAP7_75t_R FILLER_184_827 ();
 FILLER_ASAP7_75t_R FILLER_184_832 ();
 DECAPx2_ASAP7_75t_R FILLER_184_837 ();
 FILLER_ASAP7_75t_R FILLER_184_843 ();
 DECAPx1_ASAP7_75t_R FILLER_184_855 ();
 DECAPx6_ASAP7_75t_R FILLER_184_865 ();
 DECAPx1_ASAP7_75t_R FILLER_184_879 ();
 DECAPx6_ASAP7_75t_R FILLER_184_889 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_903 ();
 DECAPx4_ASAP7_75t_R FILLER_184_909 ();
 FILLER_ASAP7_75t_R FILLER_184_925 ();
 DECAPx6_ASAP7_75t_R FILLER_184_953 ();
 FILLER_ASAP7_75t_R FILLER_184_967 ();
 DECAPx1_ASAP7_75t_R FILLER_184_975 ();
 DECAPx6_ASAP7_75t_R FILLER_184_982 ();
 FILLER_ASAP7_75t_R FILLER_184_996 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_1004 ();
 DECAPx6_ASAP7_75t_R FILLER_184_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1038 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_1044 ();
 DECAPx4_ASAP7_75t_R FILLER_184_1055 ();
 FILLER_ASAP7_75t_R FILLER_184_1072 ();
 DECAPx4_ASAP7_75t_R FILLER_184_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1091 ();
 DECAPx2_ASAP7_75t_R FILLER_184_1118 ();
 FILLER_ASAP7_75t_R FILLER_184_1124 ();
 FILLER_ASAP7_75t_R FILLER_184_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1148 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1157 ();
 FILLER_ASAP7_75t_R FILLER_184_1164 ();
 DECAPx1_ASAP7_75t_R FILLER_184_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_184_1338 ();
 DECAPx6_ASAP7_75t_R FILLER_184_1360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_1374 ();
 DECAPx6_ASAP7_75t_R FILLER_185_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_16 ();
 DECAPx10_ASAP7_75t_R FILLER_185_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_45 ();
 DECAPx2_ASAP7_75t_R FILLER_185_52 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_58 ();
 FILLER_ASAP7_75t_R FILLER_185_87 ();
 DECAPx2_ASAP7_75t_R FILLER_185_95 ();
 FILLER_ASAP7_75t_R FILLER_185_107 ();
 FILLER_ASAP7_75t_R FILLER_185_117 ();
 DECAPx1_ASAP7_75t_R FILLER_185_125 ();
 DECAPx2_ASAP7_75t_R FILLER_185_135 ();
 FILLER_ASAP7_75t_R FILLER_185_151 ();
 DECAPx6_ASAP7_75t_R FILLER_185_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_170 ();
 DECAPx2_ASAP7_75t_R FILLER_185_174 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_183 ();
 DECAPx10_ASAP7_75t_R FILLER_185_194 ();
 DECAPx4_ASAP7_75t_R FILLER_185_216 ();
 FILLER_ASAP7_75t_R FILLER_185_226 ();
 DECAPx2_ASAP7_75t_R FILLER_185_234 ();
 FILLER_ASAP7_75t_R FILLER_185_262 ();
 FILLER_ASAP7_75t_R FILLER_185_270 ();
 DECAPx10_ASAP7_75t_R FILLER_185_275 ();
 DECAPx1_ASAP7_75t_R FILLER_185_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_301 ();
 DECAPx1_ASAP7_75t_R FILLER_185_308 ();
 DECAPx2_ASAP7_75t_R FILLER_185_315 ();
 FILLER_ASAP7_75t_R FILLER_185_321 ();
 DECAPx4_ASAP7_75t_R FILLER_185_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_336 ();
 DECAPx1_ASAP7_75t_R FILLER_185_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_347 ();
 DECAPx6_ASAP7_75t_R FILLER_185_374 ();
 DECAPx1_ASAP7_75t_R FILLER_185_388 ();
 FILLER_ASAP7_75t_R FILLER_185_398 ();
 DECAPx6_ASAP7_75t_R FILLER_185_403 ();
 DECAPx2_ASAP7_75t_R FILLER_185_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_423 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_430 ();
 FILLER_ASAP7_75t_R FILLER_185_439 ();
 DECAPx1_ASAP7_75t_R FILLER_185_447 ();
 DECAPx2_ASAP7_75t_R FILLER_185_477 ();
 FILLER_ASAP7_75t_R FILLER_185_491 ();
 FILLER_ASAP7_75t_R FILLER_185_499 ();
 DECAPx2_ASAP7_75t_R FILLER_185_527 ();
 FILLER_ASAP7_75t_R FILLER_185_533 ();
 FILLER_ASAP7_75t_R FILLER_185_541 ();
 FILLER_ASAP7_75t_R FILLER_185_569 ();
 FILLER_ASAP7_75t_R FILLER_185_579 ();
 DECAPx2_ASAP7_75t_R FILLER_185_589 ();
 DECAPx4_ASAP7_75t_R FILLER_185_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_611 ();
 FILLER_ASAP7_75t_R FILLER_185_620 ();
 DECAPx10_ASAP7_75t_R FILLER_185_628 ();
 DECAPx4_ASAP7_75t_R FILLER_185_650 ();
 DECAPx4_ASAP7_75t_R FILLER_185_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_678 ();
 FILLER_ASAP7_75t_R FILLER_185_705 ();
 FILLER_ASAP7_75t_R FILLER_185_714 ();
 FILLER_ASAP7_75t_R FILLER_185_722 ();
 FILLER_ASAP7_75t_R FILLER_185_727 ();
 FILLER_ASAP7_75t_R FILLER_185_751 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_759 ();
 DECAPx2_ASAP7_75t_R FILLER_185_768 ();
 DECAPx4_ASAP7_75t_R FILLER_185_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_787 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_796 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_805 ();
 DECAPx6_ASAP7_75t_R FILLER_185_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_827 ();
 DECAPx4_ASAP7_75t_R FILLER_185_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_844 ();
 DECAPx4_ASAP7_75t_R FILLER_185_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_861 ();
 DECAPx4_ASAP7_75t_R FILLER_185_870 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_880 ();
 FILLER_ASAP7_75t_R FILLER_185_889 ();
 FILLER_ASAP7_75t_R FILLER_185_899 ();
 DECAPx1_ASAP7_75t_R FILLER_185_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_908 ();
 DECAPx1_ASAP7_75t_R FILLER_185_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_916 ();
 FILLER_ASAP7_75t_R FILLER_185_923 ();
 FILLER_ASAP7_75t_R FILLER_185_927 ();
 DECAPx10_ASAP7_75t_R FILLER_185_955 ();
 DECAPx4_ASAP7_75t_R FILLER_185_977 ();
 FILLER_ASAP7_75t_R FILLER_185_987 ();
 DECAPx10_ASAP7_75t_R FILLER_185_995 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1017 ();
 DECAPx6_ASAP7_75t_R FILLER_185_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1057 ();
 FILLER_ASAP7_75t_R FILLER_185_1064 ();
 DECAPx4_ASAP7_75t_R FILLER_185_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1082 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_1091 ();
 DECAPx1_ASAP7_75t_R FILLER_185_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1110 ();
 DECAPx2_ASAP7_75t_R FILLER_185_1132 ();
 FILLER_ASAP7_75t_R FILLER_185_1138 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_1143 ();
 FILLER_ASAP7_75t_R FILLER_185_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_185_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_186_2 ();
 FILLER_ASAP7_75t_R FILLER_186_34 ();
 DECAPx4_ASAP7_75t_R FILLER_186_42 ();
 DECAPx2_ASAP7_75t_R FILLER_186_58 ();
 FILLER_ASAP7_75t_R FILLER_186_64 ();
 DECAPx1_ASAP7_75t_R FILLER_186_72 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_186_79 ();
 FILLER_ASAP7_75t_R FILLER_186_88 ();
 FILLER_ASAP7_75t_R FILLER_186_98 ();
 DECAPx1_ASAP7_75t_R FILLER_186_107 ();
 DECAPx2_ASAP7_75t_R FILLER_186_118 ();
 FILLER_ASAP7_75t_R FILLER_186_124 ();
 DECAPx6_ASAP7_75t_R FILLER_186_148 ();
 FILLER_ASAP7_75t_R FILLER_186_162 ();
 DECAPx10_ASAP7_75t_R FILLER_186_170 ();
 DECAPx6_ASAP7_75t_R FILLER_186_192 ();
 DECAPx2_ASAP7_75t_R FILLER_186_206 ();
 FILLER_ASAP7_75t_R FILLER_186_218 ();
 FILLER_ASAP7_75t_R FILLER_186_228 ();
 FILLER_ASAP7_75t_R FILLER_186_238 ();
 FILLER_ASAP7_75t_R FILLER_186_246 ();
 FILLER_ASAP7_75t_R FILLER_186_286 ();
 DECAPx6_ASAP7_75t_R FILLER_186_296 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_186_310 ();
 FILLER_ASAP7_75t_R FILLER_186_319 ();
 DECAPx10_ASAP7_75t_R FILLER_186_324 ();
 DECAPx4_ASAP7_75t_R FILLER_186_346 ();
 FILLER_ASAP7_75t_R FILLER_186_356 ();
 FILLER_ASAP7_75t_R FILLER_186_364 ();
 DECAPx6_ASAP7_75t_R FILLER_186_369 ();
 FILLER_ASAP7_75t_R FILLER_186_383 ();
 DECAPx1_ASAP7_75t_R FILLER_186_411 ();
 DECAPx10_ASAP7_75t_R FILLER_186_421 ();
 DECAPx2_ASAP7_75t_R FILLER_186_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_452 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_186_459 ();
 FILLER_ASAP7_75t_R FILLER_186_464 ();
 DECAPx1_ASAP7_75t_R FILLER_186_472 ();
 DECAPx2_ASAP7_75t_R FILLER_186_479 ();
 DECAPx4_ASAP7_75t_R FILLER_186_493 ();
 DECAPx6_ASAP7_75t_R FILLER_186_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_523 ();
 DECAPx6_ASAP7_75t_R FILLER_186_527 ();
 DECAPx2_ASAP7_75t_R FILLER_186_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_547 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_186_554 ();
 DECAPx2_ASAP7_75t_R FILLER_186_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_566 ();
 FILLER_ASAP7_75t_R FILLER_186_573 ();
 DECAPx4_ASAP7_75t_R FILLER_186_581 ();
 FILLER_ASAP7_75t_R FILLER_186_591 ();
 FILLER_ASAP7_75t_R FILLER_186_599 ();
 DECAPx2_ASAP7_75t_R FILLER_186_608 ();
 DECAPx4_ASAP7_75t_R FILLER_186_620 ();
 DECAPx4_ASAP7_75t_R FILLER_186_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_646 ();
 DECAPx2_ASAP7_75t_R FILLER_186_653 ();
 FILLER_ASAP7_75t_R FILLER_186_665 ();
 DECAPx4_ASAP7_75t_R FILLER_186_673 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_186_690 ();
 FILLER_ASAP7_75t_R FILLER_186_696 ();
 FILLER_ASAP7_75t_R FILLER_186_724 ();
 DECAPx2_ASAP7_75t_R FILLER_186_732 ();
 FILLER_ASAP7_75t_R FILLER_186_738 ();
 FILLER_ASAP7_75t_R FILLER_186_748 ();
 DECAPx2_ASAP7_75t_R FILLER_186_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_760 ();
 DECAPx2_ASAP7_75t_R FILLER_186_769 ();
 FILLER_ASAP7_75t_R FILLER_186_781 ();
 DECAPx2_ASAP7_75t_R FILLER_186_809 ();
 DECAPx6_ASAP7_75t_R FILLER_186_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_837 ();
 DECAPx2_ASAP7_75t_R FILLER_186_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_850 ();
 DECAPx2_ASAP7_75t_R FILLER_186_877 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_186_883 ();
 FILLER_ASAP7_75t_R FILLER_186_912 ();
 FILLER_ASAP7_75t_R FILLER_186_920 ();
 DECAPx2_ASAP7_75t_R FILLER_186_930 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_186_936 ();
 DECAPx1_ASAP7_75t_R FILLER_186_942 ();
 DECAPx1_ASAP7_75t_R FILLER_186_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_953 ();
 DECAPx6_ASAP7_75t_R FILLER_186_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_975 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_186_983 ();
 FILLER_ASAP7_75t_R FILLER_186_1000 ();
 FILLER_ASAP7_75t_R FILLER_186_1010 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_186_1015 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1025 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_186_1031 ();
 FILLER_ASAP7_75t_R FILLER_186_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1060 ();
 DECAPx6_ASAP7_75t_R FILLER_186_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_186_1130 ();
 FILLER_ASAP7_75t_R FILLER_186_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_186_1353 ();
 FILLER_ASAP7_75t_R FILLER_186_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_187_2 ();
 DECAPx2_ASAP7_75t_R FILLER_187_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_22 ();
 DECAPx4_ASAP7_75t_R FILLER_187_26 ();
 DECAPx2_ASAP7_75t_R FILLER_187_39 ();
 FILLER_ASAP7_75t_R FILLER_187_51 ();
 DECAPx4_ASAP7_75t_R FILLER_187_59 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_69 ();
 DECAPx2_ASAP7_75t_R FILLER_187_78 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_84 ();
 DECAPx6_ASAP7_75t_R FILLER_187_95 ();
 FILLER_ASAP7_75t_R FILLER_187_117 ();
 DECAPx6_ASAP7_75t_R FILLER_187_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_140 ();
 DECAPx2_ASAP7_75t_R FILLER_187_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_153 ();
 FILLER_ASAP7_75t_R FILLER_187_180 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_185 ();
 FILLER_ASAP7_75t_R FILLER_187_194 ();
 FILLER_ASAP7_75t_R FILLER_187_202 ();
 FILLER_ASAP7_75t_R FILLER_187_230 ();
 DECAPx4_ASAP7_75t_R FILLER_187_238 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_248 ();
 DECAPx4_ASAP7_75t_R FILLER_187_257 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_267 ();
 DECAPx1_ASAP7_75t_R FILLER_187_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_280 ();
 FILLER_ASAP7_75t_R FILLER_187_287 ();
 DECAPx2_ASAP7_75t_R FILLER_187_297 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_303 ();
 DECAPx4_ASAP7_75t_R FILLER_187_332 ();
 FILLER_ASAP7_75t_R FILLER_187_342 ();
 DECAPx10_ASAP7_75t_R FILLER_187_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_372 ();
 FILLER_ASAP7_75t_R FILLER_187_379 ();
 DECAPx1_ASAP7_75t_R FILLER_187_384 ();
 DECAPx1_ASAP7_75t_R FILLER_187_394 ();
 FILLER_ASAP7_75t_R FILLER_187_424 ();
 DECAPx10_ASAP7_75t_R FILLER_187_429 ();
 DECAPx6_ASAP7_75t_R FILLER_187_451 ();
 DECAPx10_ASAP7_75t_R FILLER_187_468 ();
 DECAPx6_ASAP7_75t_R FILLER_187_490 ();
 DECAPx1_ASAP7_75t_R FILLER_187_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_508 ();
 FILLER_ASAP7_75t_R FILLER_187_515 ();
 DECAPx6_ASAP7_75t_R FILLER_187_520 ();
 DECAPx2_ASAP7_75t_R FILLER_187_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_540 ();
 DECAPx1_ASAP7_75t_R FILLER_187_547 ();
 DECAPx10_ASAP7_75t_R FILLER_187_554 ();
 DECAPx1_ASAP7_75t_R FILLER_187_576 ();
 DECAPx1_ASAP7_75t_R FILLER_187_586 ();
 DECAPx6_ASAP7_75t_R FILLER_187_596 ();
 DECAPx1_ASAP7_75t_R FILLER_187_610 ();
 DECAPx1_ASAP7_75t_R FILLER_187_620 ();
 DECAPx4_ASAP7_75t_R FILLER_187_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_637 ();
 FILLER_ASAP7_75t_R FILLER_187_648 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_657 ();
 FILLER_ASAP7_75t_R FILLER_187_666 ();
 DECAPx6_ASAP7_75t_R FILLER_187_674 ();
 DECAPx1_ASAP7_75t_R FILLER_187_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_692 ();
 DECAPx4_ASAP7_75t_R FILLER_187_696 ();
 FILLER_ASAP7_75t_R FILLER_187_709 ();
 FILLER_ASAP7_75t_R FILLER_187_733 ();
 DECAPx6_ASAP7_75t_R FILLER_187_761 ();
 DECAPx2_ASAP7_75t_R FILLER_187_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_781 ();
 FILLER_ASAP7_75t_R FILLER_187_790 ();
 FILLER_ASAP7_75t_R FILLER_187_795 ();
 DECAPx2_ASAP7_75t_R FILLER_187_805 ();
 FILLER_ASAP7_75t_R FILLER_187_817 ();
 FILLER_ASAP7_75t_R FILLER_187_845 ();
 DECAPx2_ASAP7_75t_R FILLER_187_850 ();
 FILLER_ASAP7_75t_R FILLER_187_862 ();
 FILLER_ASAP7_75t_R FILLER_187_872 ();
 DECAPx10_ASAP7_75t_R FILLER_187_877 ();
 DECAPx2_ASAP7_75t_R FILLER_187_899 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_905 ();
 DECAPx2_ASAP7_75t_R FILLER_187_916 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_922 ();
 DECAPx1_ASAP7_75t_R FILLER_187_927 ();
 DECAPx6_ASAP7_75t_R FILLER_187_937 ();
 DECAPx1_ASAP7_75t_R FILLER_187_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_955 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_964 ();
 FILLER_ASAP7_75t_R FILLER_187_973 ();
 DECAPx2_ASAP7_75t_R FILLER_187_983 ();
 FILLER_ASAP7_75t_R FILLER_187_989 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_1017 ();
 FILLER_ASAP7_75t_R FILLER_187_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1041 ();
 DECAPx6_ASAP7_75t_R FILLER_187_1068 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_1082 ();
 FILLER_ASAP7_75t_R FILLER_187_1091 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1099 ();
 FILLER_ASAP7_75t_R FILLER_187_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1118 ();
 FILLER_ASAP7_75t_R FILLER_187_1124 ();
 FILLER_ASAP7_75t_R FILLER_187_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_187_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_187_1342 ();
 DECAPx4_ASAP7_75t_R FILLER_187_1364 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_1374 ();
 DECAPx6_ASAP7_75t_R FILLER_188_2 ();
 DECAPx1_ASAP7_75t_R FILLER_188_16 ();
 DECAPx4_ASAP7_75t_R FILLER_188_26 ();
 FILLER_ASAP7_75t_R FILLER_188_36 ();
 FILLER_ASAP7_75t_R FILLER_188_44 ();
 DECAPx6_ASAP7_75t_R FILLER_188_52 ();
 DECAPx1_ASAP7_75t_R FILLER_188_66 ();
 FILLER_ASAP7_75t_R FILLER_188_76 ();
 FILLER_ASAP7_75t_R FILLER_188_84 ();
 DECAPx4_ASAP7_75t_R FILLER_188_89 ();
 FILLER_ASAP7_75t_R FILLER_188_99 ();
 DECAPx10_ASAP7_75t_R FILLER_188_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_131 ();
 FILLER_ASAP7_75t_R FILLER_188_158 ();
 FILLER_ASAP7_75t_R FILLER_188_166 ();
 DECAPx6_ASAP7_75t_R FILLER_188_171 ();
 DECAPx6_ASAP7_75t_R FILLER_188_193 ();
 FILLER_ASAP7_75t_R FILLER_188_207 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_188_215 ();
 DECAPx6_ASAP7_75t_R FILLER_188_221 ();
 DECAPx2_ASAP7_75t_R FILLER_188_235 ();
 DECAPx2_ASAP7_75t_R FILLER_188_247 ();
 DECAPx1_ASAP7_75t_R FILLER_188_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_264 ();
 FILLER_ASAP7_75t_R FILLER_188_291 ();
 FILLER_ASAP7_75t_R FILLER_188_299 ();
 FILLER_ASAP7_75t_R FILLER_188_307 ();
 DECAPx4_ASAP7_75t_R FILLER_188_315 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_188_325 ();
 FILLER_ASAP7_75t_R FILLER_188_334 ();
 DECAPx6_ASAP7_75t_R FILLER_188_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_358 ();
 FILLER_ASAP7_75t_R FILLER_188_385 ();
 DECAPx2_ASAP7_75t_R FILLER_188_425 ();
 FILLER_ASAP7_75t_R FILLER_188_431 ();
 DECAPx6_ASAP7_75t_R FILLER_188_439 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_188_459 ();
 FILLER_ASAP7_75t_R FILLER_188_464 ();
 DECAPx6_ASAP7_75t_R FILLER_188_472 ();
 FILLER_ASAP7_75t_R FILLER_188_492 ();
 FILLER_ASAP7_75t_R FILLER_188_500 ();
 DECAPx2_ASAP7_75t_R FILLER_188_528 ();
 FILLER_ASAP7_75t_R FILLER_188_534 ();
 DECAPx2_ASAP7_75t_R FILLER_188_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_568 ();
 DECAPx1_ASAP7_75t_R FILLER_188_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_576 ();
 FILLER_ASAP7_75t_R FILLER_188_583 ();
 DECAPx6_ASAP7_75t_R FILLER_188_593 ();
 FILLER_ASAP7_75t_R FILLER_188_607 ();
 FILLER_ASAP7_75t_R FILLER_188_635 ();
 DECAPx2_ASAP7_75t_R FILLER_188_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_650 ();
 FILLER_ASAP7_75t_R FILLER_188_659 ();
 FILLER_ASAP7_75t_R FILLER_188_669 ();
 DECAPx1_ASAP7_75t_R FILLER_188_678 ();
 DECAPx10_ASAP7_75t_R FILLER_188_690 ();
 FILLER_ASAP7_75t_R FILLER_188_718 ();
 DECAPx4_ASAP7_75t_R FILLER_188_728 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_188_738 ();
 FILLER_ASAP7_75t_R FILLER_188_749 ();
 DECAPx2_ASAP7_75t_R FILLER_188_754 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_188_760 ();
 FILLER_ASAP7_75t_R FILLER_188_769 ();
 DECAPx10_ASAP7_75t_R FILLER_188_777 ();
 DECAPx10_ASAP7_75t_R FILLER_188_799 ();
 DECAPx2_ASAP7_75t_R FILLER_188_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_833 ();
 DECAPx10_ASAP7_75t_R FILLER_188_837 ();
 DECAPx4_ASAP7_75t_R FILLER_188_859 ();
 FILLER_ASAP7_75t_R FILLER_188_869 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_188_874 ();
 DECAPx1_ASAP7_75t_R FILLER_188_883 ();
 DECAPx10_ASAP7_75t_R FILLER_188_895 ();
 DECAPx6_ASAP7_75t_R FILLER_188_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_931 ();
 FILLER_ASAP7_75t_R FILLER_188_940 ();
 FILLER_ASAP7_75t_R FILLER_188_948 ();
 FILLER_ASAP7_75t_R FILLER_188_957 ();
 FILLER_ASAP7_75t_R FILLER_188_966 ();
 FILLER_ASAP7_75t_R FILLER_188_975 ();
 DECAPx10_ASAP7_75t_R FILLER_188_984 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_188_1006 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1015 ();
 FILLER_ASAP7_75t_R FILLER_188_1031 ();
 FILLER_ASAP7_75t_R FILLER_188_1041 ();
 DECAPx4_ASAP7_75t_R FILLER_188_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1059 ();
 FILLER_ASAP7_75t_R FILLER_188_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_188_1126 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_188_1141 ();
 FILLER_ASAP7_75t_R FILLER_188_1154 ();
 DECAPx2_ASAP7_75t_R FILLER_188_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_188_1351 ();
 DECAPx1_ASAP7_75t_R FILLER_188_1373 ();
 DECAPx2_ASAP7_75t_R FILLER_189_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_8 ();
 DECAPx2_ASAP7_75t_R FILLER_189_37 ();
 DECAPx6_ASAP7_75t_R FILLER_189_49 ();
 FILLER_ASAP7_75t_R FILLER_189_63 ();
 DECAPx10_ASAP7_75t_R FILLER_189_91 ();
 DECAPx2_ASAP7_75t_R FILLER_189_113 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_119 ();
 FILLER_ASAP7_75t_R FILLER_189_128 ();
 FILLER_ASAP7_75t_R FILLER_189_136 ();
 FILLER_ASAP7_75t_R FILLER_189_144 ();
 DECAPx6_ASAP7_75t_R FILLER_189_149 ();
 FILLER_ASAP7_75t_R FILLER_189_169 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_174 ();
 FILLER_ASAP7_75t_R FILLER_189_183 ();
 FILLER_ASAP7_75t_R FILLER_189_193 ();
 DECAPx4_ASAP7_75t_R FILLER_189_201 ();
 DECAPx6_ASAP7_75t_R FILLER_189_217 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_231 ();
 DECAPx10_ASAP7_75t_R FILLER_189_240 ();
 DECAPx1_ASAP7_75t_R FILLER_189_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_266 ();
 DECAPx2_ASAP7_75t_R FILLER_189_273 ();
 DECAPx6_ASAP7_75t_R FILLER_189_282 ();
 DECAPx2_ASAP7_75t_R FILLER_189_296 ();
 FILLER_ASAP7_75t_R FILLER_189_328 ();
 FILLER_ASAP7_75t_R FILLER_189_336 ();
 DECAPx2_ASAP7_75t_R FILLER_189_360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_372 ();
 DECAPx10_ASAP7_75t_R FILLER_189_378 ();
 FILLER_ASAP7_75t_R FILLER_189_406 ();
 DECAPx1_ASAP7_75t_R FILLER_189_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_422 ();
 FILLER_ASAP7_75t_R FILLER_189_449 ();
 DECAPx2_ASAP7_75t_R FILLER_189_477 ();
 FILLER_ASAP7_75t_R FILLER_189_483 ();
 DECAPx1_ASAP7_75t_R FILLER_189_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_515 ();
 FILLER_ASAP7_75t_R FILLER_189_522 ();
 DECAPx2_ASAP7_75t_R FILLER_189_532 ();
 FILLER_ASAP7_75t_R FILLER_189_544 ();
 FILLER_ASAP7_75t_R FILLER_189_552 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_580 ();
 DECAPx6_ASAP7_75t_R FILLER_189_586 ();
 FILLER_ASAP7_75t_R FILLER_189_600 ();
 DECAPx1_ASAP7_75t_R FILLER_189_608 ();
 DECAPx6_ASAP7_75t_R FILLER_189_618 ();
 DECAPx2_ASAP7_75t_R FILLER_189_632 ();
 DECAPx6_ASAP7_75t_R FILLER_189_644 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_658 ();
 DECAPx2_ASAP7_75t_R FILLER_189_669 ();
 FILLER_ASAP7_75t_R FILLER_189_675 ();
 FILLER_ASAP7_75t_R FILLER_189_683 ();
 DECAPx10_ASAP7_75t_R FILLER_189_693 ();
 DECAPx1_ASAP7_75t_R FILLER_189_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_719 ();
 DECAPx4_ASAP7_75t_R FILLER_189_728 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_738 ();
 DECAPx1_ASAP7_75t_R FILLER_189_767 ();
 DECAPx2_ASAP7_75t_R FILLER_189_779 ();
 FILLER_ASAP7_75t_R FILLER_189_785 ();
 DECAPx6_ASAP7_75t_R FILLER_189_791 ();
 DECAPx1_ASAP7_75t_R FILLER_189_805 ();
 DECAPx6_ASAP7_75t_R FILLER_189_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_826 ();
 DECAPx2_ASAP7_75t_R FILLER_189_835 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_841 ();
 FILLER_ASAP7_75t_R FILLER_189_847 ();
 DECAPx6_ASAP7_75t_R FILLER_189_857 ();
 DECAPx1_ASAP7_75t_R FILLER_189_879 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_909 ();
 DECAPx2_ASAP7_75t_R FILLER_189_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_924 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_927 ();
 FILLER_ASAP7_75t_R FILLER_189_956 ();
 DECAPx4_ASAP7_75t_R FILLER_189_961 ();
 DECAPx4_ASAP7_75t_R FILLER_189_977 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_987 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1002 ();
 DECAPx6_ASAP7_75t_R FILLER_189_1024 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1042 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1059 ();
 FILLER_ASAP7_75t_R FILLER_189_1065 ();
 FILLER_ASAP7_75t_R FILLER_189_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1096 ();
 FILLER_ASAP7_75t_R FILLER_189_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1118 ();
 FILLER_ASAP7_75t_R FILLER_189_1125 ();
 DECAPx2_ASAP7_75t_R FILLER_189_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1139 ();
 FILLER_ASAP7_75t_R FILLER_189_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_189_1350 ();
 DECAPx1_ASAP7_75t_R FILLER_189_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_1376 ();
 DECAPx4_ASAP7_75t_R FILLER_190_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_12 ();
 DECAPx1_ASAP7_75t_R FILLER_190_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_25 ();
 DECAPx10_ASAP7_75t_R FILLER_190_29 ();
 DECAPx2_ASAP7_75t_R FILLER_190_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_57 ();
 DECAPx6_ASAP7_75t_R FILLER_190_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_78 ();
 DECAPx10_ASAP7_75t_R FILLER_190_82 ();
 FILLER_ASAP7_75t_R FILLER_190_110 ();
 FILLER_ASAP7_75t_R FILLER_190_118 ();
 DECAPx4_ASAP7_75t_R FILLER_190_128 ();
 DECAPx6_ASAP7_75t_R FILLER_190_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_155 ();
 FILLER_ASAP7_75t_R FILLER_190_182 ();
 DECAPx4_ASAP7_75t_R FILLER_190_190 ();
 FILLER_ASAP7_75t_R FILLER_190_200 ();
 FILLER_ASAP7_75t_R FILLER_190_228 ();
 DECAPx1_ASAP7_75t_R FILLER_190_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_260 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_267 ();
 DECAPx6_ASAP7_75t_R FILLER_190_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_287 ();
 DECAPx6_ASAP7_75t_R FILLER_190_291 ();
 DECAPx1_ASAP7_75t_R FILLER_190_305 ();
 FILLER_ASAP7_75t_R FILLER_190_315 ();
 DECAPx6_ASAP7_75t_R FILLER_190_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_334 ();
 DECAPx2_ASAP7_75t_R FILLER_190_343 ();
 FILLER_ASAP7_75t_R FILLER_190_349 ();
 FILLER_ASAP7_75t_R FILLER_190_359 ();
 DECAPx10_ASAP7_75t_R FILLER_190_367 ();
 FILLER_ASAP7_75t_R FILLER_190_389 ();
 DECAPx4_ASAP7_75t_R FILLER_190_397 ();
 FILLER_ASAP7_75t_R FILLER_190_407 ();
 FILLER_ASAP7_75t_R FILLER_190_415 ();
 DECAPx2_ASAP7_75t_R FILLER_190_420 ();
 FILLER_ASAP7_75t_R FILLER_190_426 ();
 DECAPx1_ASAP7_75t_R FILLER_190_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_438 ();
 FILLER_ASAP7_75t_R FILLER_190_442 ();
 DECAPx6_ASAP7_75t_R FILLER_190_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_461 ();
 FILLER_ASAP7_75t_R FILLER_190_464 ();
 DECAPx1_ASAP7_75t_R FILLER_190_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_473 ();
 FILLER_ASAP7_75t_R FILLER_190_480 ();
 DECAPx1_ASAP7_75t_R FILLER_190_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_489 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_496 ();
 DECAPx6_ASAP7_75t_R FILLER_190_502 ();
 DECAPx1_ASAP7_75t_R FILLER_190_516 ();
 FILLER_ASAP7_75t_R FILLER_190_526 ();
 DECAPx6_ASAP7_75t_R FILLER_190_536 ();
 DECAPx2_ASAP7_75t_R FILLER_190_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_556 ();
 DECAPx10_ASAP7_75t_R FILLER_190_563 ();
 DECAPx6_ASAP7_75t_R FILLER_190_585 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_599 ();
 DECAPx2_ASAP7_75t_R FILLER_190_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_614 ();
 DECAPx2_ASAP7_75t_R FILLER_190_621 ();
 FILLER_ASAP7_75t_R FILLER_190_627 ();
 DECAPx4_ASAP7_75t_R FILLER_190_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_642 ();
 FILLER_ASAP7_75t_R FILLER_190_650 ();
 DECAPx6_ASAP7_75t_R FILLER_190_659 ();
 DECAPx1_ASAP7_75t_R FILLER_190_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_677 ();
 FILLER_ASAP7_75t_R FILLER_190_704 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_709 ();
 DECAPx1_ASAP7_75t_R FILLER_190_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_719 ();
 DECAPx1_ASAP7_75t_R FILLER_190_723 ();
 FILLER_ASAP7_75t_R FILLER_190_733 ();
 DECAPx6_ASAP7_75t_R FILLER_190_738 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_752 ();
 DECAPx2_ASAP7_75t_R FILLER_190_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_764 ();
 DECAPx1_ASAP7_75t_R FILLER_190_768 ();
 FILLER_ASAP7_75t_R FILLER_190_780 ();
 FILLER_ASAP7_75t_R FILLER_190_788 ();
 FILLER_ASAP7_75t_R FILLER_190_796 ();
 FILLER_ASAP7_75t_R FILLER_190_804 ();
 FILLER_ASAP7_75t_R FILLER_190_812 ();
 FILLER_ASAP7_75t_R FILLER_190_817 ();
 FILLER_ASAP7_75t_R FILLER_190_825 ();
 FILLER_ASAP7_75t_R FILLER_190_853 ();
 FILLER_ASAP7_75t_R FILLER_190_869 ();
 DECAPx2_ASAP7_75t_R FILLER_190_879 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_885 ();
 FILLER_ASAP7_75t_R FILLER_190_896 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_901 ();
 DECAPx4_ASAP7_75t_R FILLER_190_910 ();
 DECAPx6_ASAP7_75t_R FILLER_190_926 ();
 DECAPx1_ASAP7_75t_R FILLER_190_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_944 ();
 DECAPx2_ASAP7_75t_R FILLER_190_948 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_954 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_963 ();
 FILLER_ASAP7_75t_R FILLER_190_972 ();
 FILLER_ASAP7_75t_R FILLER_190_982 ();
 FILLER_ASAP7_75t_R FILLER_190_990 ();
 DECAPx6_ASAP7_75t_R FILLER_190_1018 ();
 FILLER_ASAP7_75t_R FILLER_190_1032 ();
 FILLER_ASAP7_75t_R FILLER_190_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1068 ();
 FILLER_ASAP7_75t_R FILLER_190_1074 ();
 FILLER_ASAP7_75t_R FILLER_190_1084 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1102 ();
 DECAPx6_ASAP7_75t_R FILLER_190_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_1152 ();
 FILLER_ASAP7_75t_R FILLER_190_1161 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_190_1349 ();
 DECAPx2_ASAP7_75t_R FILLER_190_1371 ();
 DECAPx10_ASAP7_75t_R FILLER_191_2 ();
 DECAPx6_ASAP7_75t_R FILLER_191_24 ();
 FILLER_ASAP7_75t_R FILLER_191_44 ();
 FILLER_ASAP7_75t_R FILLER_191_49 ();
 DECAPx4_ASAP7_75t_R FILLER_191_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_87 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_114 ();
 DECAPx10_ASAP7_75t_R FILLER_191_123 ();
 DECAPx6_ASAP7_75t_R FILLER_191_145 ();
 FILLER_ASAP7_75t_R FILLER_191_165 ();
 DECAPx6_ASAP7_75t_R FILLER_191_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_187 ();
 DECAPx4_ASAP7_75t_R FILLER_191_194 ();
 DECAPx2_ASAP7_75t_R FILLER_191_210 ();
 DECAPx4_ASAP7_75t_R FILLER_191_219 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_229 ();
 FILLER_ASAP7_75t_R FILLER_191_238 ();
 FILLER_ASAP7_75t_R FILLER_191_243 ();
 DECAPx2_ASAP7_75t_R FILLER_191_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_254 ();
 DECAPx1_ASAP7_75t_R FILLER_191_281 ();
 DECAPx2_ASAP7_75t_R FILLER_191_291 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_297 ();
 DECAPx6_ASAP7_75t_R FILLER_191_306 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_320 ();
 FILLER_ASAP7_75t_R FILLER_191_326 ();
 DECAPx2_ASAP7_75t_R FILLER_191_334 ();
 FILLER_ASAP7_75t_R FILLER_191_340 ();
 FILLER_ASAP7_75t_R FILLER_191_345 ();
 FILLER_ASAP7_75t_R FILLER_191_355 ();
 DECAPx1_ASAP7_75t_R FILLER_191_363 ();
 DECAPx4_ASAP7_75t_R FILLER_191_373 ();
 DECAPx4_ASAP7_75t_R FILLER_191_409 ();
 FILLER_ASAP7_75t_R FILLER_191_419 ();
 DECAPx6_ASAP7_75t_R FILLER_191_427 ();
 DECAPx2_ASAP7_75t_R FILLER_191_441 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_473 ();
 FILLER_ASAP7_75t_R FILLER_191_484 ();
 DECAPx1_ASAP7_75t_R FILLER_191_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_500 ();
 DECAPx6_ASAP7_75t_R FILLER_191_511 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_525 ();
 DECAPx1_ASAP7_75t_R FILLER_191_534 ();
 DECAPx4_ASAP7_75t_R FILLER_191_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_554 ();
 DECAPx4_ASAP7_75t_R FILLER_191_562 ();
 DECAPx2_ASAP7_75t_R FILLER_191_578 ();
 FILLER_ASAP7_75t_R FILLER_191_584 ();
 DECAPx2_ASAP7_75t_R FILLER_191_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_598 ();
 DECAPx2_ASAP7_75t_R FILLER_191_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_613 ();
 FILLER_ASAP7_75t_R FILLER_191_640 ();
 DECAPx10_ASAP7_75t_R FILLER_191_652 ();
 DECAPx6_ASAP7_75t_R FILLER_191_674 ();
 DECAPx1_ASAP7_75t_R FILLER_191_688 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_695 ();
 FILLER_ASAP7_75t_R FILLER_191_724 ();
 DECAPx1_ASAP7_75t_R FILLER_191_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_738 ();
 DECAPx2_ASAP7_75t_R FILLER_191_747 ();
 FILLER_ASAP7_75t_R FILLER_191_753 ();
 DECAPx2_ASAP7_75t_R FILLER_191_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_764 ();
 DECAPx10_ASAP7_75t_R FILLER_191_771 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_793 ();
 FILLER_ASAP7_75t_R FILLER_191_802 ();
 DECAPx4_ASAP7_75t_R FILLER_191_812 ();
 FILLER_ASAP7_75t_R FILLER_191_822 ();
 DECAPx2_ASAP7_75t_R FILLER_191_832 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_838 ();
 DECAPx1_ASAP7_75t_R FILLER_191_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_848 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_855 ();
 DECAPx1_ASAP7_75t_R FILLER_191_864 ();
 DECAPx4_ASAP7_75t_R FILLER_191_876 ();
 FILLER_ASAP7_75t_R FILLER_191_886 ();
 DECAPx6_ASAP7_75t_R FILLER_191_894 ();
 DECAPx2_ASAP7_75t_R FILLER_191_916 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_922 ();
 FILLER_ASAP7_75t_R FILLER_191_927 ();
 DECAPx2_ASAP7_75t_R FILLER_191_937 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_943 ();
 DECAPx2_ASAP7_75t_R FILLER_191_949 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_955 ();
 DECAPx10_ASAP7_75t_R FILLER_191_966 ();
 DECAPx6_ASAP7_75t_R FILLER_191_988 ();
 FILLER_ASAP7_75t_R FILLER_191_1002 ();
 FILLER_ASAP7_75t_R FILLER_191_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_191_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_191_1028 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1094 ();
 FILLER_ASAP7_75t_R FILLER_191_1098 ();
 FILLER_ASAP7_75t_R FILLER_191_1106 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_191_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1144 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_191_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_191_1341 ();
 DECAPx6_ASAP7_75t_R FILLER_191_1363 ();
 DECAPx6_ASAP7_75t_R FILLER_192_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_16 ();
 DECAPx1_ASAP7_75t_R FILLER_192_25 ();
 FILLER_ASAP7_75t_R FILLER_192_55 ();
 FILLER_ASAP7_75t_R FILLER_192_63 ();
 DECAPx6_ASAP7_75t_R FILLER_192_68 ();
 FILLER_ASAP7_75t_R FILLER_192_82 ();
 DECAPx4_ASAP7_75t_R FILLER_192_90 ();
 FILLER_ASAP7_75t_R FILLER_192_106 ();
 DECAPx2_ASAP7_75t_R FILLER_192_111 ();
 FILLER_ASAP7_75t_R FILLER_192_125 ();
 FILLER_ASAP7_75t_R FILLER_192_142 ();
 DECAPx4_ASAP7_75t_R FILLER_192_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_160 ();
 DECAPx2_ASAP7_75t_R FILLER_192_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_193 ();
 FILLER_ASAP7_75t_R FILLER_192_200 ();
 DECAPx2_ASAP7_75t_R FILLER_192_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_211 ();
 FILLER_ASAP7_75t_R FILLER_192_218 ();
 DECAPx10_ASAP7_75t_R FILLER_192_226 ();
 DECAPx2_ASAP7_75t_R FILLER_192_248 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_254 ();
 FILLER_ASAP7_75t_R FILLER_192_263 ();
 DECAPx2_ASAP7_75t_R FILLER_192_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_274 ();
 DECAPx1_ASAP7_75t_R FILLER_192_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_305 ();
 DECAPx2_ASAP7_75t_R FILLER_192_312 ();
 DECAPx2_ASAP7_75t_R FILLER_192_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_350 ();
 DECAPx1_ASAP7_75t_R FILLER_192_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_361 ();
 FILLER_ASAP7_75t_R FILLER_192_388 ();
 FILLER_ASAP7_75t_R FILLER_192_396 ();
 DECAPx4_ASAP7_75t_R FILLER_192_401 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_411 ();
 DECAPx4_ASAP7_75t_R FILLER_192_440 ();
 FILLER_ASAP7_75t_R FILLER_192_450 ();
 DECAPx1_ASAP7_75t_R FILLER_192_458 ();
 FILLER_ASAP7_75t_R FILLER_192_464 ();
 FILLER_ASAP7_75t_R FILLER_192_473 ();
 FILLER_ASAP7_75t_R FILLER_192_478 ();
 DECAPx2_ASAP7_75t_R FILLER_192_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_492 ();
 DECAPx10_ASAP7_75t_R FILLER_192_499 ();
 DECAPx6_ASAP7_75t_R FILLER_192_521 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_535 ();
 DECAPx4_ASAP7_75t_R FILLER_192_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_554 ();
 FILLER_ASAP7_75t_R FILLER_192_581 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_586 ();
 DECAPx1_ASAP7_75t_R FILLER_192_595 ();
 DECAPx2_ASAP7_75t_R FILLER_192_607 ();
 FILLER_ASAP7_75t_R FILLER_192_613 ();
 DECAPx2_ASAP7_75t_R FILLER_192_621 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_627 ();
 DECAPx1_ASAP7_75t_R FILLER_192_637 ();
 DECAPx4_ASAP7_75t_R FILLER_192_647 ();
 FILLER_ASAP7_75t_R FILLER_192_664 ();
 DECAPx2_ASAP7_75t_R FILLER_192_672 ();
 DECAPx1_ASAP7_75t_R FILLER_192_684 ();
 DECAPx10_ASAP7_75t_R FILLER_192_696 ();
 FILLER_ASAP7_75t_R FILLER_192_718 ();
 DECAPx6_ASAP7_75t_R FILLER_192_726 ();
 FILLER_ASAP7_75t_R FILLER_192_766 ();
 DECAPx10_ASAP7_75t_R FILLER_192_776 ();
 DECAPx6_ASAP7_75t_R FILLER_192_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_812 ();
 DECAPx1_ASAP7_75t_R FILLER_192_819 ();
 DECAPx10_ASAP7_75t_R FILLER_192_829 ();
 DECAPx6_ASAP7_75t_R FILLER_192_851 ();
 FILLER_ASAP7_75t_R FILLER_192_865 ();
 DECAPx10_ASAP7_75t_R FILLER_192_873 ();
 DECAPx2_ASAP7_75t_R FILLER_192_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_901 ();
 DECAPx1_ASAP7_75t_R FILLER_192_928 ();
 DECAPx1_ASAP7_75t_R FILLER_192_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_962 ();
 DECAPx6_ASAP7_75t_R FILLER_192_989 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_192_1010 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_1016 ();
 FILLER_ASAP7_75t_R FILLER_192_1026 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_1035 ();
 DECAPx4_ASAP7_75t_R FILLER_192_1049 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1077 ();
 DECAPx4_ASAP7_75t_R FILLER_192_1084 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_1094 ();
 FILLER_ASAP7_75t_R FILLER_192_1105 ();
 FILLER_ASAP7_75t_R FILLER_192_1133 ();
 DECAPx1_ASAP7_75t_R FILLER_192_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_192_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_192_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_192_1341 ();
 DECAPx6_ASAP7_75t_R FILLER_192_1363 ();
 DECAPx2_ASAP7_75t_R FILLER_193_2 ();
 FILLER_ASAP7_75t_R FILLER_193_8 ();
 FILLER_ASAP7_75t_R FILLER_193_36 ();
 DECAPx4_ASAP7_75t_R FILLER_193_44 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_54 ();
 DECAPx2_ASAP7_75t_R FILLER_193_60 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_72 ();
 DECAPx6_ASAP7_75t_R FILLER_193_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_115 ();
 FILLER_ASAP7_75t_R FILLER_193_122 ();
 DECAPx2_ASAP7_75t_R FILLER_193_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_133 ();
 DECAPx4_ASAP7_75t_R FILLER_193_160 ();
 FILLER_ASAP7_75t_R FILLER_193_176 ();
 DECAPx1_ASAP7_75t_R FILLER_193_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_185 ();
 FILLER_ASAP7_75t_R FILLER_193_212 ();
 DECAPx1_ASAP7_75t_R FILLER_193_217 ();
 DECAPx2_ASAP7_75t_R FILLER_193_229 ();
 DECAPx4_ASAP7_75t_R FILLER_193_241 ();
 FILLER_ASAP7_75t_R FILLER_193_251 ();
 DECAPx6_ASAP7_75t_R FILLER_193_263 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_277 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_286 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_292 ();
 FILLER_ASAP7_75t_R FILLER_193_321 ();
 DECAPx1_ASAP7_75t_R FILLER_193_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_333 ();
 FILLER_ASAP7_75t_R FILLER_193_340 ();
 DECAPx1_ASAP7_75t_R FILLER_193_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_349 ();
 DECAPx4_ASAP7_75t_R FILLER_193_356 ();
 DECAPx1_ASAP7_75t_R FILLER_193_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_376 ();
 DECAPx6_ASAP7_75t_R FILLER_193_380 ();
 DECAPx2_ASAP7_75t_R FILLER_193_394 ();
 DECAPx4_ASAP7_75t_R FILLER_193_406 ();
 DECAPx1_ASAP7_75t_R FILLER_193_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_426 ();
 FILLER_ASAP7_75t_R FILLER_193_430 ();
 DECAPx4_ASAP7_75t_R FILLER_193_440 ();
 DECAPx2_ASAP7_75t_R FILLER_193_456 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_462 ();
 FILLER_ASAP7_75t_R FILLER_193_472 ();
 FILLER_ASAP7_75t_R FILLER_193_481 ();
 FILLER_ASAP7_75t_R FILLER_193_489 ();
 DECAPx2_ASAP7_75t_R FILLER_193_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_503 ();
 DECAPx4_ASAP7_75t_R FILLER_193_510 ();
 FILLER_ASAP7_75t_R FILLER_193_520 ();
 DECAPx1_ASAP7_75t_R FILLER_193_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_534 ();
 FILLER_ASAP7_75t_R FILLER_193_543 ();
 DECAPx1_ASAP7_75t_R FILLER_193_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_556 ();
 DECAPx2_ASAP7_75t_R FILLER_193_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_569 ();
 FILLER_ASAP7_75t_R FILLER_193_576 ();
 DECAPx6_ASAP7_75t_R FILLER_193_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_600 ();
 DECAPx6_ASAP7_75t_R FILLER_193_604 ();
 DECAPx2_ASAP7_75t_R FILLER_193_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_624 ();
 DECAPx10_ASAP7_75t_R FILLER_193_631 ();
 DECAPx2_ASAP7_75t_R FILLER_193_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_659 ();
 DECAPx2_ASAP7_75t_R FILLER_193_667 ();
 FILLER_ASAP7_75t_R FILLER_193_673 ();
 FILLER_ASAP7_75t_R FILLER_193_683 ();
 FILLER_ASAP7_75t_R FILLER_193_711 ();
 DECAPx6_ASAP7_75t_R FILLER_193_719 ();
 DECAPx10_ASAP7_75t_R FILLER_193_736 ();
 DECAPx2_ASAP7_75t_R FILLER_193_758 ();
 FILLER_ASAP7_75t_R FILLER_193_764 ();
 DECAPx2_ASAP7_75t_R FILLER_193_774 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_780 ();
 DECAPx2_ASAP7_75t_R FILLER_193_791 ();
 FILLER_ASAP7_75t_R FILLER_193_797 ();
 FILLER_ASAP7_75t_R FILLER_193_805 ();
 DECAPx6_ASAP7_75t_R FILLER_193_813 ();
 DECAPx4_ASAP7_75t_R FILLER_193_833 ();
 FILLER_ASAP7_75t_R FILLER_193_843 ();
 DECAPx6_ASAP7_75t_R FILLER_193_851 ();
 DECAPx2_ASAP7_75t_R FILLER_193_865 ();
 DECAPx2_ASAP7_75t_R FILLER_193_878 ();
 FILLER_ASAP7_75t_R FILLER_193_884 ();
 DECAPx10_ASAP7_75t_R FILLER_193_892 ();
 FILLER_ASAP7_75t_R FILLER_193_914 ();
 DECAPx2_ASAP7_75t_R FILLER_193_919 ();
 FILLER_ASAP7_75t_R FILLER_193_927 ();
 FILLER_ASAP7_75t_R FILLER_193_935 ();
 DECAPx2_ASAP7_75t_R FILLER_193_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_949 ();
 DECAPx10_ASAP7_75t_R FILLER_193_953 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_975 ();
 FILLER_ASAP7_75t_R FILLER_193_981 ();
 DECAPx4_ASAP7_75t_R FILLER_193_989 ();
 FILLER_ASAP7_75t_R FILLER_193_999 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1042 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1060 ();
 FILLER_ASAP7_75t_R FILLER_193_1067 ();
 FILLER_ASAP7_75t_R FILLER_193_1076 ();
 FILLER_ASAP7_75t_R FILLER_193_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1114 ();
 FILLER_ASAP7_75t_R FILLER_193_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1125 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_1131 ();
 FILLER_ASAP7_75t_R FILLER_193_1143 ();
 DECAPx2_ASAP7_75t_R FILLER_193_1155 ();
 FILLER_ASAP7_75t_R FILLER_193_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_193_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_193_1350 ();
 DECAPx1_ASAP7_75t_R FILLER_193_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_1376 ();
 DECAPx4_ASAP7_75t_R FILLER_194_2 ();
 FILLER_ASAP7_75t_R FILLER_194_12 ();
 DECAPx1_ASAP7_75t_R FILLER_194_20 ();
 DECAPx4_ASAP7_75t_R FILLER_194_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_37 ();
 DECAPx4_ASAP7_75t_R FILLER_194_44 ();
 FILLER_ASAP7_75t_R FILLER_194_54 ();
 FILLER_ASAP7_75t_R FILLER_194_62 ();
 DECAPx2_ASAP7_75t_R FILLER_194_72 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_78 ();
 FILLER_ASAP7_75t_R FILLER_194_87 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_96 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_102 ();
 DECAPx4_ASAP7_75t_R FILLER_194_131 ();
 FILLER_ASAP7_75t_R FILLER_194_147 ();
 DECAPx6_ASAP7_75t_R FILLER_194_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_166 ();
 DECAPx6_ASAP7_75t_R FILLER_194_173 ();
 FILLER_ASAP7_75t_R FILLER_194_187 ();
 DECAPx4_ASAP7_75t_R FILLER_194_192 ();
 DECAPx4_ASAP7_75t_R FILLER_194_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_234 ();
 DECAPx2_ASAP7_75t_R FILLER_194_243 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_249 ();
 FILLER_ASAP7_75t_R FILLER_194_259 ();
 DECAPx2_ASAP7_75t_R FILLER_194_267 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_273 ();
 DECAPx2_ASAP7_75t_R FILLER_194_282 ();
 DECAPx6_ASAP7_75t_R FILLER_194_291 ();
 DECAPx1_ASAP7_75t_R FILLER_194_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_309 ();
 DECAPx6_ASAP7_75t_R FILLER_194_313 ();
 DECAPx1_ASAP7_75t_R FILLER_194_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_331 ();
 DECAPx10_ASAP7_75t_R FILLER_194_358 ();
 DECAPx4_ASAP7_75t_R FILLER_194_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_390 ();
 DECAPx2_ASAP7_75t_R FILLER_194_417 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_423 ();
 FILLER_ASAP7_75t_R FILLER_194_432 ();
 DECAPx1_ASAP7_75t_R FILLER_194_442 ();
 FILLER_ASAP7_75t_R FILLER_194_452 ();
 FILLER_ASAP7_75t_R FILLER_194_460 ();
 FILLER_ASAP7_75t_R FILLER_194_464 ();
 DECAPx2_ASAP7_75t_R FILLER_194_473 ();
 FILLER_ASAP7_75t_R FILLER_194_479 ();
 DECAPx2_ASAP7_75t_R FILLER_194_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_495 ();
 FILLER_ASAP7_75t_R FILLER_194_522 ();
 DECAPx2_ASAP7_75t_R FILLER_194_532 ();
 DECAPx4_ASAP7_75t_R FILLER_194_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_570 ();
 FILLER_ASAP7_75t_R FILLER_194_579 ();
 DECAPx4_ASAP7_75t_R FILLER_194_587 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_597 ();
 FILLER_ASAP7_75t_R FILLER_194_606 ();
 DECAPx4_ASAP7_75t_R FILLER_194_611 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_621 ();
 DECAPx4_ASAP7_75t_R FILLER_194_650 ();
 DECAPx4_ASAP7_75t_R FILLER_194_666 ();
 FILLER_ASAP7_75t_R FILLER_194_676 ();
 DECAPx6_ASAP7_75t_R FILLER_194_686 ();
 DECAPx1_ASAP7_75t_R FILLER_194_703 ();
 FILLER_ASAP7_75t_R FILLER_194_713 ();
 DECAPx1_ASAP7_75t_R FILLER_194_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_724 ();
 FILLER_ASAP7_75t_R FILLER_194_728 ();
 FILLER_ASAP7_75t_R FILLER_194_738 ();
 DECAPx2_ASAP7_75t_R FILLER_194_746 ();
 DECAPx2_ASAP7_75t_R FILLER_194_758 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_764 ();
 DECAPx4_ASAP7_75t_R FILLER_194_773 ();
 FILLER_ASAP7_75t_R FILLER_194_783 ();
 FILLER_ASAP7_75t_R FILLER_194_811 ();
 DECAPx1_ASAP7_75t_R FILLER_194_821 ();
 FILLER_ASAP7_75t_R FILLER_194_831 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_859 ();
 FILLER_ASAP7_75t_R FILLER_194_868 ();
 DECAPx2_ASAP7_75t_R FILLER_194_878 ();
 FILLER_ASAP7_75t_R FILLER_194_884 ();
 FILLER_ASAP7_75t_R FILLER_194_896 ();
 DECAPx10_ASAP7_75t_R FILLER_194_908 ();
 DECAPx4_ASAP7_75t_R FILLER_194_930 ();
 FILLER_ASAP7_75t_R FILLER_194_946 ();
 DECAPx2_ASAP7_75t_R FILLER_194_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_960 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_975 ();
 FILLER_ASAP7_75t_R FILLER_194_985 ();
 FILLER_ASAP7_75t_R FILLER_194_993 ();
 FILLER_ASAP7_75t_R FILLER_194_1001 ();
 DECAPx4_ASAP7_75t_R FILLER_194_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1020 ();
 FILLER_ASAP7_75t_R FILLER_194_1027 ();
 DECAPx4_ASAP7_75t_R FILLER_194_1035 ();
 DECAPx4_ASAP7_75t_R FILLER_194_1051 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_1061 ();
 FILLER_ASAP7_75t_R FILLER_194_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_194_1080 ();
 FILLER_ASAP7_75t_R FILLER_194_1086 ();
 FILLER_ASAP7_75t_R FILLER_194_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1123 ();
 FILLER_ASAP7_75t_R FILLER_194_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_194_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_194_1350 ();
 DECAPx1_ASAP7_75t_R FILLER_194_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_195_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_8 ();
 DECAPx10_ASAP7_75t_R FILLER_195_17 ();
 FILLER_ASAP7_75t_R FILLER_195_47 ();
 FILLER_ASAP7_75t_R FILLER_195_55 ();
 DECAPx6_ASAP7_75t_R FILLER_195_63 ();
 FILLER_ASAP7_75t_R FILLER_195_77 ();
 DECAPx2_ASAP7_75t_R FILLER_195_85 ();
 FILLER_ASAP7_75t_R FILLER_195_113 ();
 FILLER_ASAP7_75t_R FILLER_195_121 ();
 DECAPx10_ASAP7_75t_R FILLER_195_126 ();
 DECAPx4_ASAP7_75t_R FILLER_195_148 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_158 ();
 FILLER_ASAP7_75t_R FILLER_195_187 ();
 FILLER_ASAP7_75t_R FILLER_195_195 ();
 DECAPx2_ASAP7_75t_R FILLER_195_205 ();
 FILLER_ASAP7_75t_R FILLER_195_211 ();
 FILLER_ASAP7_75t_R FILLER_195_221 ();
 DECAPx2_ASAP7_75t_R FILLER_195_245 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_251 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_262 ();
 FILLER_ASAP7_75t_R FILLER_195_271 ();
 DECAPx2_ASAP7_75t_R FILLER_195_299 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_305 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_314 ();
 DECAPx10_ASAP7_75t_R FILLER_195_320 ();
 DECAPx1_ASAP7_75t_R FILLER_195_342 ();
 DECAPx1_ASAP7_75t_R FILLER_195_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_353 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_357 ();
 FILLER_ASAP7_75t_R FILLER_195_366 ();
 FILLER_ASAP7_75t_R FILLER_195_374 ();
 DECAPx1_ASAP7_75t_R FILLER_195_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_386 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_390 ();
 DECAPx2_ASAP7_75t_R FILLER_195_399 ();
 DECAPx2_ASAP7_75t_R FILLER_195_408 ();
 FILLER_ASAP7_75t_R FILLER_195_414 ();
 DECAPx6_ASAP7_75t_R FILLER_195_419 ();
 DECAPx4_ASAP7_75t_R FILLER_195_439 ();
 FILLER_ASAP7_75t_R FILLER_195_475 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_480 ();
 DECAPx2_ASAP7_75t_R FILLER_195_491 ();
 FILLER_ASAP7_75t_R FILLER_195_497 ();
 DECAPx2_ASAP7_75t_R FILLER_195_505 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_514 ();
 FILLER_ASAP7_75t_R FILLER_195_523 ();
 FILLER_ASAP7_75t_R FILLER_195_531 ();
 DECAPx1_ASAP7_75t_R FILLER_195_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_543 ();
 FILLER_ASAP7_75t_R FILLER_195_570 ();
 DECAPx6_ASAP7_75t_R FILLER_195_575 ();
 DECAPx1_ASAP7_75t_R FILLER_195_589 ();
 DECAPx1_ASAP7_75t_R FILLER_195_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_623 ();
 DECAPx2_ASAP7_75t_R FILLER_195_630 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_636 ();
 DECAPx1_ASAP7_75t_R FILLER_195_642 ();
 DECAPx4_ASAP7_75t_R FILLER_195_649 ();
 DECAPx2_ASAP7_75t_R FILLER_195_666 ();
 FILLER_ASAP7_75t_R FILLER_195_678 ();
 DECAPx4_ASAP7_75t_R FILLER_195_688 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_698 ();
 FILLER_ASAP7_75t_R FILLER_195_711 ();
 FILLER_ASAP7_75t_R FILLER_195_739 ();
 FILLER_ASAP7_75t_R FILLER_195_747 ();
 FILLER_ASAP7_75t_R FILLER_195_757 ();
 FILLER_ASAP7_75t_R FILLER_195_762 ();
 FILLER_ASAP7_75t_R FILLER_195_790 ();
 DECAPx1_ASAP7_75t_R FILLER_195_795 ();
 DECAPx2_ASAP7_75t_R FILLER_195_802 ();
 DECAPx2_ASAP7_75t_R FILLER_195_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_822 ();
 FILLER_ASAP7_75t_R FILLER_195_831 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_839 ();
 FILLER_ASAP7_75t_R FILLER_195_850 ();
 FILLER_ASAP7_75t_R FILLER_195_855 ();
 FILLER_ASAP7_75t_R FILLER_195_860 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_868 ();
 DECAPx2_ASAP7_75t_R FILLER_195_878 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_884 ();
 DECAPx1_ASAP7_75t_R FILLER_195_893 ();
 FILLER_ASAP7_75t_R FILLER_195_905 ();
 FILLER_ASAP7_75t_R FILLER_195_913 ();
 DECAPx1_ASAP7_75t_R FILLER_195_921 ();
 FILLER_ASAP7_75t_R FILLER_195_927 ();
 FILLER_ASAP7_75t_R FILLER_195_935 ();
 DECAPx2_ASAP7_75t_R FILLER_195_943 ();
 DECAPx1_ASAP7_75t_R FILLER_195_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_961 ();
 DECAPx6_ASAP7_75t_R FILLER_195_965 ();
 FILLER_ASAP7_75t_R FILLER_195_986 ();
 DECAPx2_ASAP7_75t_R FILLER_195_996 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_1002 ();
 FILLER_ASAP7_75t_R FILLER_195_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1020 ();
 DECAPx4_ASAP7_75t_R FILLER_195_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1050 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1068 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1088 ();
 DECAPx1_ASAP7_75t_R FILLER_195_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1102 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1112 ();
 FILLER_ASAP7_75t_R FILLER_195_1126 ();
 DECAPx4_ASAP7_75t_R FILLER_195_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1143 ();
 DECAPx6_ASAP7_75t_R FILLER_195_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_195_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_195_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_195_1343 ();
 DECAPx4_ASAP7_75t_R FILLER_195_1365 ();
 FILLER_ASAP7_75t_R FILLER_195_1375 ();
 FILLER_ASAP7_75t_R FILLER_196_2 ();
 FILLER_ASAP7_75t_R FILLER_196_30 ();
 DECAPx1_ASAP7_75t_R FILLER_196_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_39 ();
 DECAPx4_ASAP7_75t_R FILLER_196_48 ();
 FILLER_ASAP7_75t_R FILLER_196_58 ();
 DECAPx2_ASAP7_75t_R FILLER_196_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_74 ();
 FILLER_ASAP7_75t_R FILLER_196_81 ();
 FILLER_ASAP7_75t_R FILLER_196_90 ();
 FILLER_ASAP7_75t_R FILLER_196_100 ();
 FILLER_ASAP7_75t_R FILLER_196_109 ();
 DECAPx1_ASAP7_75t_R FILLER_196_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_121 ();
 FILLER_ASAP7_75t_R FILLER_196_128 ();
 DECAPx4_ASAP7_75t_R FILLER_196_136 ();
 DECAPx4_ASAP7_75t_R FILLER_196_152 ();
 DECAPx2_ASAP7_75t_R FILLER_196_168 ();
 FILLER_ASAP7_75t_R FILLER_196_174 ();
 DECAPx1_ASAP7_75t_R FILLER_196_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_183 ();
 DECAPx2_ASAP7_75t_R FILLER_196_191 ();
 FILLER_ASAP7_75t_R FILLER_196_205 ();
 DECAPx1_ASAP7_75t_R FILLER_196_213 ();
 FILLER_ASAP7_75t_R FILLER_196_223 ();
 FILLER_ASAP7_75t_R FILLER_196_231 ();
 DECAPx2_ASAP7_75t_R FILLER_196_241 ();
 FILLER_ASAP7_75t_R FILLER_196_253 ();
 DECAPx2_ASAP7_75t_R FILLER_196_270 ();
 DECAPx2_ASAP7_75t_R FILLER_196_288 ();
 FILLER_ASAP7_75t_R FILLER_196_300 ();
 FILLER_ASAP7_75t_R FILLER_196_328 ();
 DECAPx10_ASAP7_75t_R FILLER_196_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_355 ();
 DECAPx2_ASAP7_75t_R FILLER_196_364 ();
 FILLER_ASAP7_75t_R FILLER_196_370 ();
 DECAPx1_ASAP7_75t_R FILLER_196_398 ();
 DECAPx4_ASAP7_75t_R FILLER_196_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_418 ();
 FILLER_ASAP7_75t_R FILLER_196_425 ();
 DECAPx10_ASAP7_75t_R FILLER_196_433 ();
 DECAPx2_ASAP7_75t_R FILLER_196_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_461 ();
 FILLER_ASAP7_75t_R FILLER_196_464 ();
 FILLER_ASAP7_75t_R FILLER_196_473 ();
 DECAPx1_ASAP7_75t_R FILLER_196_478 ();
 DECAPx10_ASAP7_75t_R FILLER_196_488 ();
 DECAPx10_ASAP7_75t_R FILLER_196_510 ();
 DECAPx4_ASAP7_75t_R FILLER_196_532 ();
 FILLER_ASAP7_75t_R FILLER_196_542 ();
 FILLER_ASAP7_75t_R FILLER_196_550 ();
 FILLER_ASAP7_75t_R FILLER_196_558 ();
 DECAPx6_ASAP7_75t_R FILLER_196_563 ();
 DECAPx1_ASAP7_75t_R FILLER_196_577 ();
 DECAPx1_ASAP7_75t_R FILLER_196_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_595 ();
 DECAPx10_ASAP7_75t_R FILLER_196_602 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_196_624 ();
 DECAPx2_ASAP7_75t_R FILLER_196_653 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_196_659 ();
 DECAPx1_ASAP7_75t_R FILLER_196_688 ();
 DECAPx10_ASAP7_75t_R FILLER_196_698 ();
 DECAPx2_ASAP7_75t_R FILLER_196_720 ();
 FILLER_ASAP7_75t_R FILLER_196_726 ();
 FILLER_ASAP7_75t_R FILLER_196_734 ();
 DECAPx2_ASAP7_75t_R FILLER_196_742 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_196_748 ();
 DECAPx1_ASAP7_75t_R FILLER_196_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_781 ();
 DECAPx6_ASAP7_75t_R FILLER_196_788 ();
 DECAPx2_ASAP7_75t_R FILLER_196_802 ();
 DECAPx10_ASAP7_75t_R FILLER_196_814 ();
 DECAPx1_ASAP7_75t_R FILLER_196_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_840 ();
 DECAPx6_ASAP7_75t_R FILLER_196_847 ();
 DECAPx2_ASAP7_75t_R FILLER_196_861 ();
 DECAPx10_ASAP7_75t_R FILLER_196_873 ();
 DECAPx6_ASAP7_75t_R FILLER_196_895 ();
 DECAPx1_ASAP7_75t_R FILLER_196_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_913 ();
 FILLER_ASAP7_75t_R FILLER_196_921 ();
 DECAPx2_ASAP7_75t_R FILLER_196_930 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_196_936 ();
 FILLER_ASAP7_75t_R FILLER_196_946 ();
 DECAPx10_ASAP7_75t_R FILLER_196_974 ();
 DECAPx4_ASAP7_75t_R FILLER_196_996 ();
 FILLER_ASAP7_75t_R FILLER_196_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_196_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_196_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1033 ();
 FILLER_ASAP7_75t_R FILLER_196_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1051 ();
 FILLER_ASAP7_75t_R FILLER_196_1065 ();
 DECAPx6_ASAP7_75t_R FILLER_196_1073 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_196_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_196_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_1100 ();
 FILLER_ASAP7_75t_R FILLER_196_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_196_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_196_1146 ();
 DECAPx4_ASAP7_75t_R FILLER_196_1158 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_196_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_196_1351 ();
 DECAPx1_ASAP7_75t_R FILLER_196_1373 ();
 DECAPx2_ASAP7_75t_R FILLER_197_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_197_14 ();
 DECAPx10_ASAP7_75t_R FILLER_197_20 ();
 DECAPx2_ASAP7_75t_R FILLER_197_42 ();
 DECAPx2_ASAP7_75t_R FILLER_197_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_60 ();
 FILLER_ASAP7_75t_R FILLER_197_68 ();
 DECAPx4_ASAP7_75t_R FILLER_197_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_86 ();
 FILLER_ASAP7_75t_R FILLER_197_95 ();
 DECAPx6_ASAP7_75t_R FILLER_197_104 ();
 DECAPx1_ASAP7_75t_R FILLER_197_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_122 ();
 FILLER_ASAP7_75t_R FILLER_197_149 ();
 DECAPx2_ASAP7_75t_R FILLER_197_157 ();
 FILLER_ASAP7_75t_R FILLER_197_163 ();
 FILLER_ASAP7_75t_R FILLER_197_171 ();
 DECAPx6_ASAP7_75t_R FILLER_197_176 ();
 DECAPx2_ASAP7_75t_R FILLER_197_190 ();
 DECAPx1_ASAP7_75t_R FILLER_197_218 ();
 DECAPx2_ASAP7_75t_R FILLER_197_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_235 ();
 DECAPx2_ASAP7_75t_R FILLER_197_242 ();
 FILLER_ASAP7_75t_R FILLER_197_248 ();
 FILLER_ASAP7_75t_R FILLER_197_256 ();
 FILLER_ASAP7_75t_R FILLER_197_265 ();
 FILLER_ASAP7_75t_R FILLER_197_274 ();
 FILLER_ASAP7_75t_R FILLER_197_283 ();
 FILLER_ASAP7_75t_R FILLER_197_291 ();
 FILLER_ASAP7_75t_R FILLER_197_315 ();
 DECAPx4_ASAP7_75t_R FILLER_197_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_333 ();
 DECAPx2_ASAP7_75t_R FILLER_197_340 ();
 FILLER_ASAP7_75t_R FILLER_197_354 ();
 FILLER_ASAP7_75t_R FILLER_197_378 ();
 DECAPx1_ASAP7_75t_R FILLER_197_386 ();
 FILLER_ASAP7_75t_R FILLER_197_393 ();
 FILLER_ASAP7_75t_R FILLER_197_421 ();
 DECAPx1_ASAP7_75t_R FILLER_197_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_435 ();
 DECAPx10_ASAP7_75t_R FILLER_197_442 ();
 DECAPx2_ASAP7_75t_R FILLER_197_464 ();
 FILLER_ASAP7_75t_R FILLER_197_470 ();
 FILLER_ASAP7_75t_R FILLER_197_478 ();
 DECAPx6_ASAP7_75t_R FILLER_197_486 ();
 DECAPx1_ASAP7_75t_R FILLER_197_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_504 ();
 DECAPx2_ASAP7_75t_R FILLER_197_511 ();
 FILLER_ASAP7_75t_R FILLER_197_517 ();
 DECAPx6_ASAP7_75t_R FILLER_197_522 ();
 FILLER_ASAP7_75t_R FILLER_197_536 ();
 DECAPx10_ASAP7_75t_R FILLER_197_544 ();
 DECAPx1_ASAP7_75t_R FILLER_197_566 ();
 DECAPx10_ASAP7_75t_R FILLER_197_596 ();
 DECAPx2_ASAP7_75t_R FILLER_197_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_624 ();
 FILLER_ASAP7_75t_R FILLER_197_631 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_197_639 ();
 DECAPx4_ASAP7_75t_R FILLER_197_645 ();
 FILLER_ASAP7_75t_R FILLER_197_655 ();
 DECAPx6_ASAP7_75t_R FILLER_197_663 ();
 DECAPx4_ASAP7_75t_R FILLER_197_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_690 ();
 FILLER_ASAP7_75t_R FILLER_197_698 ();
 DECAPx10_ASAP7_75t_R FILLER_197_710 ();
 DECAPx10_ASAP7_75t_R FILLER_197_732 ();
 DECAPx4_ASAP7_75t_R FILLER_197_754 ();
 FILLER_ASAP7_75t_R FILLER_197_778 ();
 DECAPx6_ASAP7_75t_R FILLER_197_783 ();
 DECAPx2_ASAP7_75t_R FILLER_197_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_803 ();
 DECAPx6_ASAP7_75t_R FILLER_197_812 ();
 DECAPx10_ASAP7_75t_R FILLER_197_834 ();
 DECAPx2_ASAP7_75t_R FILLER_197_856 ();
 DECAPx1_ASAP7_75t_R FILLER_197_869 ();
 DECAPx10_ASAP7_75t_R FILLER_197_880 ();
 DECAPx4_ASAP7_75t_R FILLER_197_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_912 ();
 DECAPx2_ASAP7_75t_R FILLER_197_919 ();
 FILLER_ASAP7_75t_R FILLER_197_927 ();
 DECAPx10_ASAP7_75t_R FILLER_197_935 ();
 DECAPx6_ASAP7_75t_R FILLER_197_957 ();
 FILLER_ASAP7_75t_R FILLER_197_977 ();
 DECAPx10_ASAP7_75t_R FILLER_197_985 ();
 DECAPx1_ASAP7_75t_R FILLER_197_1007 ();
 DECAPx4_ASAP7_75t_R FILLER_197_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_197_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1057 ();
 DECAPx6_ASAP7_75t_R FILLER_197_1084 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1104 ();
 FILLER_ASAP7_75t_R FILLER_197_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_197_1119 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_197_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_197_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_197_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_197_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_197_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_197_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_197_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_197_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_197_1343 ();
 DECAPx4_ASAP7_75t_R FILLER_197_1365 ();
 FILLER_ASAP7_75t_R FILLER_197_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_198_2 ();
 DECAPx2_ASAP7_75t_R FILLER_198_16 ();
 DECAPx2_ASAP7_75t_R FILLER_198_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_34 ();
 FILLER_ASAP7_75t_R FILLER_198_41 ();
 DECAPx6_ASAP7_75t_R FILLER_198_51 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_65 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_74 ();
 DECAPx1_ASAP7_75t_R FILLER_198_85 ();
 DECAPx2_ASAP7_75t_R FILLER_198_96 ();
 FILLER_ASAP7_75t_R FILLER_198_110 ();
 DECAPx2_ASAP7_75t_R FILLER_198_118 ();
 FILLER_ASAP7_75t_R FILLER_198_124 ();
 FILLER_ASAP7_75t_R FILLER_198_136 ();
 FILLER_ASAP7_75t_R FILLER_198_141 ();
 FILLER_ASAP7_75t_R FILLER_198_149 ();
 FILLER_ASAP7_75t_R FILLER_198_157 ();
 DECAPx2_ASAP7_75t_R FILLER_198_185 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_191 ();
 FILLER_ASAP7_75t_R FILLER_198_202 ();
 DECAPx2_ASAP7_75t_R FILLER_198_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_216 ();
 DECAPx6_ASAP7_75t_R FILLER_198_233 ();
 DECAPx2_ASAP7_75t_R FILLER_198_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_253 ();
 DECAPx6_ASAP7_75t_R FILLER_198_257 ();
 FILLER_ASAP7_75t_R FILLER_198_278 ();
 DECAPx1_ASAP7_75t_R FILLER_198_306 ();
 FILLER_ASAP7_75t_R FILLER_198_336 ();
 DECAPx1_ASAP7_75t_R FILLER_198_346 ();
 FILLER_ASAP7_75t_R FILLER_198_356 ();
 DECAPx2_ASAP7_75t_R FILLER_198_380 ();
 FILLER_ASAP7_75t_R FILLER_198_386 ();
 FILLER_ASAP7_75t_R FILLER_198_395 ();
 FILLER_ASAP7_75t_R FILLER_198_403 ();
 FILLER_ASAP7_75t_R FILLER_198_411 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_416 ();
 FILLER_ASAP7_75t_R FILLER_198_427 ();
 DECAPx4_ASAP7_75t_R FILLER_198_439 ();
 FILLER_ASAP7_75t_R FILLER_198_455 ();
 FILLER_ASAP7_75t_R FILLER_198_460 ();
 DECAPx1_ASAP7_75t_R FILLER_198_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_468 ();
 FILLER_ASAP7_75t_R FILLER_198_495 ();
 DECAPx2_ASAP7_75t_R FILLER_198_523 ();
 DECAPx6_ASAP7_75t_R FILLER_198_555 ();
 FILLER_ASAP7_75t_R FILLER_198_569 ();
 DECAPx1_ASAP7_75t_R FILLER_198_577 ();
 FILLER_ASAP7_75t_R FILLER_198_587 ();
 DECAPx1_ASAP7_75t_R FILLER_198_615 ();
 DECAPx10_ASAP7_75t_R FILLER_198_625 ();
 DECAPx6_ASAP7_75t_R FILLER_198_653 ();
 DECAPx6_ASAP7_75t_R FILLER_198_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_687 ();
 DECAPx4_ASAP7_75t_R FILLER_198_698 ();
 FILLER_ASAP7_75t_R FILLER_198_714 ();
 FILLER_ASAP7_75t_R FILLER_198_730 ();
 FILLER_ASAP7_75t_R FILLER_198_740 ();
 FILLER_ASAP7_75t_R FILLER_198_750 ();
 DECAPx2_ASAP7_75t_R FILLER_198_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_764 ();
 DECAPx6_ASAP7_75t_R FILLER_198_768 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_782 ();
 FILLER_ASAP7_75t_R FILLER_198_791 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_799 ();
 FILLER_ASAP7_75t_R FILLER_198_828 ();
 DECAPx2_ASAP7_75t_R FILLER_198_839 ();
 FILLER_ASAP7_75t_R FILLER_198_845 ();
 FILLER_ASAP7_75t_R FILLER_198_853 ();
 DECAPx4_ASAP7_75t_R FILLER_198_861 ();
 FILLER_ASAP7_75t_R FILLER_198_871 ();
 DECAPx6_ASAP7_75t_R FILLER_198_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_895 ();
 FILLER_ASAP7_75t_R FILLER_198_903 ();
 DECAPx2_ASAP7_75t_R FILLER_198_911 ();
 DECAPx2_ASAP7_75t_R FILLER_198_923 ();
 FILLER_ASAP7_75t_R FILLER_198_929 ();
 DECAPx6_ASAP7_75t_R FILLER_198_938 ();
 FILLER_ASAP7_75t_R FILLER_198_952 ();
 DECAPx6_ASAP7_75t_R FILLER_198_960 ();
 DECAPx2_ASAP7_75t_R FILLER_198_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_987 ();
 FILLER_ASAP7_75t_R FILLER_198_994 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1003 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_1013 ();
 FILLER_ASAP7_75t_R FILLER_198_1042 ();
 DECAPx6_ASAP7_75t_R FILLER_198_1047 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_1061 ();
 FILLER_ASAP7_75t_R FILLER_198_1067 ();
 FILLER_ASAP7_75t_R FILLER_198_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1103 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1125 ();
 FILLER_ASAP7_75t_R FILLER_198_1139 ();
 DECAPx4_ASAP7_75t_R FILLER_198_1150 ();
 FILLER_ASAP7_75t_R FILLER_198_1160 ();
 DECAPx1_ASAP7_75t_R FILLER_198_1172 ();
 FILLER_ASAP7_75t_R FILLER_198_1182 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_198_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_198_1369 ();
 FILLER_ASAP7_75t_R FILLER_198_1375 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_2 ();
 FILLER_ASAP7_75t_R FILLER_199_31 ();
 DECAPx2_ASAP7_75t_R FILLER_199_39 ();
 FILLER_ASAP7_75t_R FILLER_199_45 ();
 FILLER_ASAP7_75t_R FILLER_199_53 ();
 DECAPx1_ASAP7_75t_R FILLER_199_58 ();
 DECAPx2_ASAP7_75t_R FILLER_199_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_76 ();
 DECAPx1_ASAP7_75t_R FILLER_199_88 ();
 FILLER_ASAP7_75t_R FILLER_199_98 ();
 DECAPx2_ASAP7_75t_R FILLER_199_108 ();
 FILLER_ASAP7_75t_R FILLER_199_120 ();
 DECAPx6_ASAP7_75t_R FILLER_199_128 ();
 FILLER_ASAP7_75t_R FILLER_199_142 ();
 FILLER_ASAP7_75t_R FILLER_199_150 ();
 FILLER_ASAP7_75t_R FILLER_199_170 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_178 ();
 FILLER_ASAP7_75t_R FILLER_199_184 ();
 FILLER_ASAP7_75t_R FILLER_199_192 ();
 FILLER_ASAP7_75t_R FILLER_199_202 ();
 DECAPx2_ASAP7_75t_R FILLER_199_210 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_224 ();
 DECAPx2_ASAP7_75t_R FILLER_199_253 ();
 DECAPx6_ASAP7_75t_R FILLER_199_262 ();
 DECAPx2_ASAP7_75t_R FILLER_199_283 ();
 FILLER_ASAP7_75t_R FILLER_199_289 ();
 FILLER_ASAP7_75t_R FILLER_199_297 ();
 DECAPx4_ASAP7_75t_R FILLER_199_302 ();
 DECAPx2_ASAP7_75t_R FILLER_199_318 ();
 FILLER_ASAP7_75t_R FILLER_199_327 ();
 FILLER_ASAP7_75t_R FILLER_199_335 ();
 DECAPx4_ASAP7_75t_R FILLER_199_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_355 ();
 DECAPx2_ASAP7_75t_R FILLER_199_362 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_368 ();
 DECAPx2_ASAP7_75t_R FILLER_199_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_403 ();
 DECAPx6_ASAP7_75t_R FILLER_199_410 ();
 DECAPx2_ASAP7_75t_R FILLER_199_424 ();
 FILLER_ASAP7_75t_R FILLER_199_436 ();
 FILLER_ASAP7_75t_R FILLER_199_444 ();
 DECAPx2_ASAP7_75t_R FILLER_199_472 ();
 FILLER_ASAP7_75t_R FILLER_199_484 ();
 DECAPx4_ASAP7_75t_R FILLER_199_489 ();
 DECAPx2_ASAP7_75t_R FILLER_199_505 ();
 DECAPx1_ASAP7_75t_R FILLER_199_514 ();
 FILLER_ASAP7_75t_R FILLER_199_524 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_529 ();
 DECAPx1_ASAP7_75t_R FILLER_199_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_542 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_546 ();
 FILLER_ASAP7_75t_R FILLER_199_552 ();
 FILLER_ASAP7_75t_R FILLER_199_560 ();
 DECAPx1_ASAP7_75t_R FILLER_199_568 ();
 DECAPx2_ASAP7_75t_R FILLER_199_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_584 ();
 DECAPx1_ASAP7_75t_R FILLER_199_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_592 ();
 DECAPx1_ASAP7_75t_R FILLER_199_599 ();
 DECAPx1_ASAP7_75t_R FILLER_199_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_610 ();
 FILLER_ASAP7_75t_R FILLER_199_614 ();
 DECAPx10_ASAP7_75t_R FILLER_199_624 ();
 DECAPx6_ASAP7_75t_R FILLER_199_654 ();
 DECAPx4_ASAP7_75t_R FILLER_199_675 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_685 ();
 DECAPx2_ASAP7_75t_R FILLER_199_700 ();
 FILLER_ASAP7_75t_R FILLER_199_718 ();
 DECAPx6_ASAP7_75t_R FILLER_199_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_740 ();
 FILLER_ASAP7_75t_R FILLER_199_751 ();
 DECAPx6_ASAP7_75t_R FILLER_199_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_773 ();
 FILLER_ASAP7_75t_R FILLER_199_780 ();
 DECAPx6_ASAP7_75t_R FILLER_199_788 ();
 FILLER_ASAP7_75t_R FILLER_199_802 ();
 DECAPx2_ASAP7_75t_R FILLER_199_810 ();
 DECAPx1_ASAP7_75t_R FILLER_199_819 ();
 DECAPx1_ASAP7_75t_R FILLER_199_826 ();
 DECAPx2_ASAP7_75t_R FILLER_199_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_862 ();
 FILLER_ASAP7_75t_R FILLER_199_871 ();
 DECAPx2_ASAP7_75t_R FILLER_199_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_886 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_895 ();
 DECAPx2_ASAP7_75t_R FILLER_199_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_910 ();
 DECAPx2_ASAP7_75t_R FILLER_199_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_924 ();
 DECAPx2_ASAP7_75t_R FILLER_199_927 ();
 FILLER_ASAP7_75t_R FILLER_199_933 ();
 DECAPx2_ASAP7_75t_R FILLER_199_943 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_949 ();
 FILLER_ASAP7_75t_R FILLER_199_959 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_971 ();
 DECAPx6_ASAP7_75t_R FILLER_199_980 ();
 FILLER_ASAP7_75t_R FILLER_199_1000 ();
 DECAPx4_ASAP7_75t_R FILLER_199_1008 ();
 DECAPx1_ASAP7_75t_R FILLER_199_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1056 ();
 FILLER_ASAP7_75t_R FILLER_199_1062 ();
 FILLER_ASAP7_75t_R FILLER_199_1071 ();
 DECAPx4_ASAP7_75t_R FILLER_199_1081 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1094 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1114 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1124 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1133 ();
 FILLER_ASAP7_75t_R FILLER_199_1155 ();
 FILLER_ASAP7_75t_R FILLER_199_1165 ();
 FILLER_ASAP7_75t_R FILLER_199_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_199_1334 ();
 DECAPx6_ASAP7_75t_R FILLER_199_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_199_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_200_2 ();
 FILLER_ASAP7_75t_R FILLER_200_8 ();
 DECAPx1_ASAP7_75t_R FILLER_200_16 ();
 DECAPx2_ASAP7_75t_R FILLER_200_23 ();
 FILLER_ASAP7_75t_R FILLER_200_29 ();
 DECAPx2_ASAP7_75t_R FILLER_200_34 ();
 FILLER_ASAP7_75t_R FILLER_200_40 ();
 DECAPx10_ASAP7_75t_R FILLER_200_50 ();
 DECAPx1_ASAP7_75t_R FILLER_200_78 ();
 DECAPx10_ASAP7_75t_R FILLER_200_88 ();
 DECAPx4_ASAP7_75t_R FILLER_200_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_146 ();
 DECAPx2_ASAP7_75t_R FILLER_200_157 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_200_163 ();
 FILLER_ASAP7_75t_R FILLER_200_192 ();
 DECAPx4_ASAP7_75t_R FILLER_200_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_210 ();
 DECAPx4_ASAP7_75t_R FILLER_200_219 ();
 FILLER_ASAP7_75t_R FILLER_200_235 ();
 FILLER_ASAP7_75t_R FILLER_200_243 ();
 DECAPx1_ASAP7_75t_R FILLER_200_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_275 ();
 DECAPx2_ASAP7_75t_R FILLER_200_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_288 ();
 FILLER_ASAP7_75t_R FILLER_200_295 ();
 DECAPx10_ASAP7_75t_R FILLER_200_303 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_200_325 ();
 DECAPx10_ASAP7_75t_R FILLER_200_334 ();
 DECAPx1_ASAP7_75t_R FILLER_200_356 ();
 DECAPx2_ASAP7_75t_R FILLER_200_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_372 ();
 DECAPx2_ASAP7_75t_R FILLER_200_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_385 ();
 FILLER_ASAP7_75t_R FILLER_200_394 ();
 FILLER_ASAP7_75t_R FILLER_200_402 ();
 DECAPx10_ASAP7_75t_R FILLER_200_416 ();
 DECAPx2_ASAP7_75t_R FILLER_200_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_444 ();
 DECAPx4_ASAP7_75t_R FILLER_200_452 ();
 FILLER_ASAP7_75t_R FILLER_200_464 ();
 DECAPx6_ASAP7_75t_R FILLER_200_472 ();
 FILLER_ASAP7_75t_R FILLER_200_486 ();
 DECAPx6_ASAP7_75t_R FILLER_200_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_508 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_200_535 ();
 DECAPx2_ASAP7_75t_R FILLER_200_544 ();
 FILLER_ASAP7_75t_R FILLER_200_558 ();
 DECAPx10_ASAP7_75t_R FILLER_200_568 ();
 DECAPx10_ASAP7_75t_R FILLER_200_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_612 ();
 DECAPx2_ASAP7_75t_R FILLER_200_621 ();
 DECAPx1_ASAP7_75t_R FILLER_200_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_637 ();
 FILLER_ASAP7_75t_R FILLER_200_645 ();
 DECAPx4_ASAP7_75t_R FILLER_200_655 ();
 FILLER_ASAP7_75t_R FILLER_200_672 ();
 DECAPx2_ASAP7_75t_R FILLER_200_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_686 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_200_695 ();
 DECAPx2_ASAP7_75t_R FILLER_200_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_707 ();
 DECAPx4_ASAP7_75t_R FILLER_200_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_728 ();
 FILLER_ASAP7_75t_R FILLER_200_736 ();
 FILLER_ASAP7_75t_R FILLER_200_744 ();
 DECAPx6_ASAP7_75t_R FILLER_200_752 ();
 DECAPx2_ASAP7_75t_R FILLER_200_766 ();
 DECAPx1_ASAP7_75t_R FILLER_200_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_782 ();
 DECAPx10_ASAP7_75t_R FILLER_200_789 ();
 DECAPx10_ASAP7_75t_R FILLER_200_811 ();
 DECAPx4_ASAP7_75t_R FILLER_200_833 ();
 FILLER_ASAP7_75t_R FILLER_200_843 ();
 FILLER_ASAP7_75t_R FILLER_200_848 ();
 FILLER_ASAP7_75t_R FILLER_200_856 ();
 DECAPx1_ASAP7_75t_R FILLER_200_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_868 ();
 DECAPx1_ASAP7_75t_R FILLER_200_875 ();
 FILLER_ASAP7_75t_R FILLER_200_885 ();
 DECAPx1_ASAP7_75t_R FILLER_200_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_897 ();
 DECAPx2_ASAP7_75t_R FILLER_200_905 ();
 DECAPx6_ASAP7_75t_R FILLER_200_918 ();
 FILLER_ASAP7_75t_R FILLER_200_932 ();
 FILLER_ASAP7_75t_R FILLER_200_940 ();
 FILLER_ASAP7_75t_R FILLER_200_948 ();
 FILLER_ASAP7_75t_R FILLER_200_958 ();
 DECAPx2_ASAP7_75t_R FILLER_200_972 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_200_978 ();
 FILLER_ASAP7_75t_R FILLER_200_988 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_200_996 ();
 DECAPx4_ASAP7_75t_R FILLER_200_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_200_1021 ();
 FILLER_ASAP7_75t_R FILLER_200_1035 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1044 ();
 DECAPx4_ASAP7_75t_R FILLER_200_1056 ();
 FILLER_ASAP7_75t_R FILLER_200_1066 ();
 DECAPx6_ASAP7_75t_R FILLER_200_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_200_1090 ();
 FILLER_ASAP7_75t_R FILLER_200_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_200_1109 ();
 FILLER_ASAP7_75t_R FILLER_200_1119 ();
 DECAPx4_ASAP7_75t_R FILLER_200_1131 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_200_1141 ();
 DECAPx1_ASAP7_75t_R FILLER_200_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_200_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_200_1369 ();
 FILLER_ASAP7_75t_R FILLER_200_1375 ();
 FILLER_ASAP7_75t_R FILLER_201_2 ();
 DECAPx4_ASAP7_75t_R FILLER_201_30 ();
 FILLER_ASAP7_75t_R FILLER_201_40 ();
 DECAPx6_ASAP7_75t_R FILLER_201_48 ();
 DECAPx6_ASAP7_75t_R FILLER_201_68 ();
 DECAPx2_ASAP7_75t_R FILLER_201_82 ();
 FILLER_ASAP7_75t_R FILLER_201_94 ();
 FILLER_ASAP7_75t_R FILLER_201_102 ();
 DECAPx2_ASAP7_75t_R FILLER_201_107 ();
 DECAPx1_ASAP7_75t_R FILLER_201_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_123 ();
 FILLER_ASAP7_75t_R FILLER_201_127 ();
 FILLER_ASAP7_75t_R FILLER_201_155 ();
 DECAPx1_ASAP7_75t_R FILLER_201_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_167 ();
 DECAPx2_ASAP7_75t_R FILLER_201_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_180 ();
 DECAPx10_ASAP7_75t_R FILLER_201_184 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_206 ();
 FILLER_ASAP7_75t_R FILLER_201_215 ();
 DECAPx1_ASAP7_75t_R FILLER_201_226 ();
 DECAPx2_ASAP7_75t_R FILLER_201_236 ();
 DECAPx2_ASAP7_75t_R FILLER_201_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_251 ();
 DECAPx2_ASAP7_75t_R FILLER_201_258 ();
 FILLER_ASAP7_75t_R FILLER_201_264 ();
 DECAPx1_ASAP7_75t_R FILLER_201_292 ();
 FILLER_ASAP7_75t_R FILLER_201_302 ();
 DECAPx2_ASAP7_75t_R FILLER_201_314 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_320 ();
 FILLER_ASAP7_75t_R FILLER_201_349 ();
 DECAPx4_ASAP7_75t_R FILLER_201_357 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_367 ();
 DECAPx4_ASAP7_75t_R FILLER_201_376 ();
 DECAPx6_ASAP7_75t_R FILLER_201_396 ();
 DECAPx4_ASAP7_75t_R FILLER_201_416 ();
 DECAPx1_ASAP7_75t_R FILLER_201_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_433 ();
 FILLER_ASAP7_75t_R FILLER_201_444 ();
 DECAPx2_ASAP7_75t_R FILLER_201_454 ();
 FILLER_ASAP7_75t_R FILLER_201_460 ();
 DECAPx2_ASAP7_75t_R FILLER_201_472 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_478 ();
 DECAPx1_ASAP7_75t_R FILLER_201_507 ();
 DECAPx2_ASAP7_75t_R FILLER_201_517 ();
 FILLER_ASAP7_75t_R FILLER_201_523 ();
 FILLER_ASAP7_75t_R FILLER_201_528 ();
 DECAPx1_ASAP7_75t_R FILLER_201_548 ();
 DECAPx2_ASAP7_75t_R FILLER_201_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_564 ();
 DECAPx2_ASAP7_75t_R FILLER_201_571 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_577 ();
 DECAPx2_ASAP7_75t_R FILLER_201_586 ();
 DECAPx2_ASAP7_75t_R FILLER_201_598 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_604 ();
 FILLER_ASAP7_75t_R FILLER_201_613 ();
 DECAPx2_ASAP7_75t_R FILLER_201_618 ();
 FILLER_ASAP7_75t_R FILLER_201_630 ();
 DECAPx1_ASAP7_75t_R FILLER_201_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_642 ();
 FILLER_ASAP7_75t_R FILLER_201_649 ();
 DECAPx4_ASAP7_75t_R FILLER_201_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_667 ();
 DECAPx2_ASAP7_75t_R FILLER_201_675 ();
 FILLER_ASAP7_75t_R FILLER_201_681 ();
 DECAPx1_ASAP7_75t_R FILLER_201_709 ();
 DECAPx4_ASAP7_75t_R FILLER_201_716 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_726 ();
 DECAPx4_ASAP7_75t_R FILLER_201_741 ();
 FILLER_ASAP7_75t_R FILLER_201_751 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_763 ();
 DECAPx4_ASAP7_75t_R FILLER_201_772 ();
 DECAPx2_ASAP7_75t_R FILLER_201_788 ();
 DECAPx4_ASAP7_75t_R FILLER_201_802 ();
 DECAPx1_ASAP7_75t_R FILLER_201_819 ();
 DECAPx1_ASAP7_75t_R FILLER_201_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_833 ();
 DECAPx10_ASAP7_75t_R FILLER_201_840 ();
 DECAPx4_ASAP7_75t_R FILLER_201_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_872 ();
 DECAPx4_ASAP7_75t_R FILLER_201_880 ();
 DECAPx6_ASAP7_75t_R FILLER_201_896 ();
 DECAPx1_ASAP7_75t_R FILLER_201_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_914 ();
 FILLER_ASAP7_75t_R FILLER_201_923 ();
 FILLER_ASAP7_75t_R FILLER_201_927 ();
 FILLER_ASAP7_75t_R FILLER_201_941 ();
 FILLER_ASAP7_75t_R FILLER_201_951 ();
 DECAPx10_ASAP7_75t_R FILLER_201_959 ();
 DECAPx4_ASAP7_75t_R FILLER_201_988 ();
 FILLER_ASAP7_75t_R FILLER_201_998 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_201_1020 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_1026 ();
 FILLER_ASAP7_75t_R FILLER_201_1055 ();
 DECAPx6_ASAP7_75t_R FILLER_201_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1079 ();
 DECAPx4_ASAP7_75t_R FILLER_201_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_201_1102 ();
 FILLER_ASAP7_75t_R FILLER_201_1132 ();
 FILLER_ASAP7_75t_R FILLER_201_1142 ();
 DECAPx4_ASAP7_75t_R FILLER_201_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_201_1342 ();
 DECAPx4_ASAP7_75t_R FILLER_201_1364 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_1374 ();
 DECAPx1_ASAP7_75t_R FILLER_202_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_6 ();
 DECAPx1_ASAP7_75t_R FILLER_202_13 ();
 DECAPx4_ASAP7_75t_R FILLER_202_20 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_30 ();
 DECAPx4_ASAP7_75t_R FILLER_202_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_49 ();
 FILLER_ASAP7_75t_R FILLER_202_53 ();
 DECAPx2_ASAP7_75t_R FILLER_202_63 ();
 DECAPx2_ASAP7_75t_R FILLER_202_75 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_81 ();
 DECAPx10_ASAP7_75t_R FILLER_202_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_132 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_139 ();
 FILLER_ASAP7_75t_R FILLER_202_145 ();
 DECAPx2_ASAP7_75t_R FILLER_202_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_163 ();
 DECAPx10_ASAP7_75t_R FILLER_202_170 ();
 DECAPx6_ASAP7_75t_R FILLER_202_192 ();
 DECAPx1_ASAP7_75t_R FILLER_202_206 ();
 DECAPx10_ASAP7_75t_R FILLER_202_216 ();
 DECAPx10_ASAP7_75t_R FILLER_202_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_260 ();
 FILLER_ASAP7_75t_R FILLER_202_267 ();
 DECAPx2_ASAP7_75t_R FILLER_202_275 ();
 DECAPx2_ASAP7_75t_R FILLER_202_284 ();
 FILLER_ASAP7_75t_R FILLER_202_290 ();
 DECAPx2_ASAP7_75t_R FILLER_202_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_304 ();
 DECAPx2_ASAP7_75t_R FILLER_202_315 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_321 ();
 DECAPx2_ASAP7_75t_R FILLER_202_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_336 ();
 FILLER_ASAP7_75t_R FILLER_202_340 ();
 FILLER_ASAP7_75t_R FILLER_202_348 ();
 FILLER_ASAP7_75t_R FILLER_202_358 ();
 DECAPx10_ASAP7_75t_R FILLER_202_366 ();
 DECAPx6_ASAP7_75t_R FILLER_202_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_402 ();
 FILLER_ASAP7_75t_R FILLER_202_429 ();
 DECAPx6_ASAP7_75t_R FILLER_202_439 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_459 ();
 FILLER_ASAP7_75t_R FILLER_202_464 ();
 DECAPx4_ASAP7_75t_R FILLER_202_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_482 ();
 DECAPx2_ASAP7_75t_R FILLER_202_489 ();
 DECAPx1_ASAP7_75t_R FILLER_202_498 ();
 DECAPx6_ASAP7_75t_R FILLER_202_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_522 ();
 FILLER_ASAP7_75t_R FILLER_202_545 ();
 FILLER_ASAP7_75t_R FILLER_202_555 ();
 DECAPx2_ASAP7_75t_R FILLER_202_563 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_569 ();
 DECAPx2_ASAP7_75t_R FILLER_202_578 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_610 ();
 DECAPx2_ASAP7_75t_R FILLER_202_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_627 ();
 DECAPx2_ASAP7_75t_R FILLER_202_634 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_640 ();
 DECAPx4_ASAP7_75t_R FILLER_202_649 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_659 ();
 DECAPx6_ASAP7_75t_R FILLER_202_668 ();
 DECAPx2_ASAP7_75t_R FILLER_202_682 ();
 DECAPx6_ASAP7_75t_R FILLER_202_694 ();
 DECAPx2_ASAP7_75t_R FILLER_202_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_714 ();
 DECAPx10_ASAP7_75t_R FILLER_202_725 ();
 DECAPx1_ASAP7_75t_R FILLER_202_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_751 ();
 FILLER_ASAP7_75t_R FILLER_202_758 ();
 FILLER_ASAP7_75t_R FILLER_202_766 ();
 DECAPx1_ASAP7_75t_R FILLER_202_776 ();
 DECAPx1_ASAP7_75t_R FILLER_202_786 ();
 DECAPx2_ASAP7_75t_R FILLER_202_796 ();
 FILLER_ASAP7_75t_R FILLER_202_812 ();
 FILLER_ASAP7_75t_R FILLER_202_820 ();
 DECAPx2_ASAP7_75t_R FILLER_202_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_834 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_843 ();
 FILLER_ASAP7_75t_R FILLER_202_855 ();
 DECAPx1_ASAP7_75t_R FILLER_202_869 ();
 DECAPx2_ASAP7_75t_R FILLER_202_885 ();
 FILLER_ASAP7_75t_R FILLER_202_891 ();
 DECAPx1_ASAP7_75t_R FILLER_202_900 ();
 DECAPx2_ASAP7_75t_R FILLER_202_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_916 ();
 FILLER_ASAP7_75t_R FILLER_202_943 ();
 DECAPx1_ASAP7_75t_R FILLER_202_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_956 ();
 DECAPx4_ASAP7_75t_R FILLER_202_968 ();
 FILLER_ASAP7_75t_R FILLER_202_978 ();
 DECAPx6_ASAP7_75t_R FILLER_202_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1000 ();
 DECAPx4_ASAP7_75t_R FILLER_202_1008 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1033 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1046 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1062 ();
 FILLER_ASAP7_75t_R FILLER_202_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1104 ();
 FILLER_ASAP7_75t_R FILLER_202_1126 ();
 DECAPx4_ASAP7_75t_R FILLER_202_1131 ();
 FILLER_ASAP7_75t_R FILLER_202_1153 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_202_1334 ();
 DECAPx6_ASAP7_75t_R FILLER_202_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_202_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_203_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_24 ();
 DECAPx2_ASAP7_75t_R FILLER_203_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_57 ();
 FILLER_ASAP7_75t_R FILLER_203_64 ();
 DECAPx1_ASAP7_75t_R FILLER_203_92 ();
 DECAPx10_ASAP7_75t_R FILLER_203_118 ();
 DECAPx10_ASAP7_75t_R FILLER_203_140 ();
 DECAPx1_ASAP7_75t_R FILLER_203_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_192 ();
 DECAPx2_ASAP7_75t_R FILLER_203_201 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_203_207 ();
 FILLER_ASAP7_75t_R FILLER_203_218 ();
 DECAPx6_ASAP7_75t_R FILLER_203_226 ();
 FILLER_ASAP7_75t_R FILLER_203_240 ();
 DECAPx4_ASAP7_75t_R FILLER_203_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_258 ();
 DECAPx1_ASAP7_75t_R FILLER_203_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_289 ();
 DECAPx1_ASAP7_75t_R FILLER_203_296 ();
 DECAPx10_ASAP7_75t_R FILLER_203_306 ();
 DECAPx4_ASAP7_75t_R FILLER_203_334 ();
 FILLER_ASAP7_75t_R FILLER_203_344 ();
 DECAPx1_ASAP7_75t_R FILLER_203_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_353 ();
 DECAPx4_ASAP7_75t_R FILLER_203_362 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_203_372 ();
 DECAPx2_ASAP7_75t_R FILLER_203_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_387 ();
 DECAPx4_ASAP7_75t_R FILLER_203_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_404 ();
 DECAPx1_ASAP7_75t_R FILLER_203_411 ();
 FILLER_ASAP7_75t_R FILLER_203_418 ();
 FILLER_ASAP7_75t_R FILLER_203_426 ();
 DECAPx6_ASAP7_75t_R FILLER_203_434 ();
 DECAPx2_ASAP7_75t_R FILLER_203_474 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_203_486 ();
 FILLER_ASAP7_75t_R FILLER_203_492 ();
 FILLER_ASAP7_75t_R FILLER_203_500 ();
 DECAPx2_ASAP7_75t_R FILLER_203_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_516 ();
 FILLER_ASAP7_75t_R FILLER_203_543 ();
 DECAPx10_ASAP7_75t_R FILLER_203_553 ();
 DECAPx4_ASAP7_75t_R FILLER_203_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_585 ();
 DECAPx2_ASAP7_75t_R FILLER_203_592 ();
 DECAPx4_ASAP7_75t_R FILLER_203_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_611 ();
 DECAPx4_ASAP7_75t_R FILLER_203_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_628 ();
 DECAPx2_ASAP7_75t_R FILLER_203_655 ();
 FILLER_ASAP7_75t_R FILLER_203_661 ();
 DECAPx4_ASAP7_75t_R FILLER_203_670 ();
 DECAPx1_ASAP7_75t_R FILLER_203_683 ();
 FILLER_ASAP7_75t_R FILLER_203_697 ();
 DECAPx1_ASAP7_75t_R FILLER_203_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_709 ();
 DECAPx2_ASAP7_75t_R FILLER_203_716 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_203_722 ();
 DECAPx1_ASAP7_75t_R FILLER_203_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_738 ();
 DECAPx1_ASAP7_75t_R FILLER_203_749 ();
 FILLER_ASAP7_75t_R FILLER_203_759 ();
 DECAPx10_ASAP7_75t_R FILLER_203_767 ();
 FILLER_ASAP7_75t_R FILLER_203_789 ();
 DECAPx6_ASAP7_75t_R FILLER_203_797 ();
 DECAPx1_ASAP7_75t_R FILLER_203_811 ();
 DECAPx2_ASAP7_75t_R FILLER_203_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_832 ();
 FILLER_ASAP7_75t_R FILLER_203_859 ();
 DECAPx10_ASAP7_75t_R FILLER_203_869 ();
 DECAPx6_ASAP7_75t_R FILLER_203_891 ();
 DECAPx1_ASAP7_75t_R FILLER_203_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_909 ();
 DECAPx2_ASAP7_75t_R FILLER_203_917 ();
 FILLER_ASAP7_75t_R FILLER_203_923 ();
 DECAPx1_ASAP7_75t_R FILLER_203_927 ();
 DECAPx6_ASAP7_75t_R FILLER_203_934 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_203_948 ();
 DECAPx4_ASAP7_75t_R FILLER_203_960 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_203_970 ();
 DECAPx2_ASAP7_75t_R FILLER_203_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_985 ();
 FILLER_ASAP7_75t_R FILLER_203_998 ();
 DECAPx6_ASAP7_75t_R FILLER_203_1006 ();
 FILLER_ASAP7_75t_R FILLER_203_1020 ();
 FILLER_ASAP7_75t_R FILLER_203_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_203_1033 ();
 DECAPx6_ASAP7_75t_R FILLER_203_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1054 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_203_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1132 ();
 DECAPx2_ASAP7_75t_R FILLER_203_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1160 ();
 DECAPx1_ASAP7_75t_R FILLER_203_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_203_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_1376 ();
 FILLER_ASAP7_75t_R FILLER_204_2 ();
 FILLER_ASAP7_75t_R FILLER_204_10 ();
 DECAPx4_ASAP7_75t_R FILLER_204_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_28 ();
 DECAPx1_ASAP7_75t_R FILLER_204_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_39 ();
 DECAPx4_ASAP7_75t_R FILLER_204_43 ();
 DECAPx2_ASAP7_75t_R FILLER_204_59 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_65 ();
 DECAPx2_ASAP7_75t_R FILLER_204_74 ();
 DECAPx6_ASAP7_75t_R FILLER_204_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_97 ();
 DECAPx2_ASAP7_75t_R FILLER_204_101 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_107 ();
 DECAPx10_ASAP7_75t_R FILLER_204_136 ();
 DECAPx4_ASAP7_75t_R FILLER_204_158 ();
 FILLER_ASAP7_75t_R FILLER_204_168 ();
 DECAPx1_ASAP7_75t_R FILLER_204_176 ();
 FILLER_ASAP7_75t_R FILLER_204_183 ();
 FILLER_ASAP7_75t_R FILLER_204_191 ();
 DECAPx2_ASAP7_75t_R FILLER_204_201 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_207 ();
 DECAPx4_ASAP7_75t_R FILLER_204_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_228 ();
 DECAPx4_ASAP7_75t_R FILLER_204_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_265 ();
 FILLER_ASAP7_75t_R FILLER_204_272 ();
 DECAPx4_ASAP7_75t_R FILLER_204_277 ();
 DECAPx2_ASAP7_75t_R FILLER_204_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_319 ();
 DECAPx10_ASAP7_75t_R FILLER_204_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_368 ();
 DECAPx6_ASAP7_75t_R FILLER_204_395 ();
 DECAPx4_ASAP7_75t_R FILLER_204_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_425 ();
 DECAPx10_ASAP7_75t_R FILLER_204_432 ();
 DECAPx2_ASAP7_75t_R FILLER_204_454 ();
 FILLER_ASAP7_75t_R FILLER_204_460 ();
 DECAPx1_ASAP7_75t_R FILLER_204_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_468 ();
 FILLER_ASAP7_75t_R FILLER_204_472 ();
 DECAPx1_ASAP7_75t_R FILLER_204_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_504 ();
 DECAPx1_ASAP7_75t_R FILLER_204_513 ();
 FILLER_ASAP7_75t_R FILLER_204_523 ();
 DECAPx2_ASAP7_75t_R FILLER_204_531 ();
 DECAPx4_ASAP7_75t_R FILLER_204_543 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_553 ();
 DECAPx2_ASAP7_75t_R FILLER_204_562 ();
 FILLER_ASAP7_75t_R FILLER_204_568 ();
 DECAPx10_ASAP7_75t_R FILLER_204_578 ();
 DECAPx10_ASAP7_75t_R FILLER_204_600 ();
 DECAPx1_ASAP7_75t_R FILLER_204_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_626 ();
 DECAPx2_ASAP7_75t_R FILLER_204_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_639 ();
 FILLER_ASAP7_75t_R FILLER_204_643 ();
 DECAPx6_ASAP7_75t_R FILLER_204_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_665 ();
 FILLER_ASAP7_75t_R FILLER_204_692 ();
 DECAPx1_ASAP7_75t_R FILLER_204_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_710 ();
 DECAPx1_ASAP7_75t_R FILLER_204_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_721 ();
 FILLER_ASAP7_75t_R FILLER_204_742 ();
 DECAPx10_ASAP7_75t_R FILLER_204_753 ();
 DECAPx6_ASAP7_75t_R FILLER_204_781 ();
 DECAPx6_ASAP7_75t_R FILLER_204_801 ();
 DECAPx2_ASAP7_75t_R FILLER_204_815 ();
 DECAPx6_ASAP7_75t_R FILLER_204_827 ();
 DECAPx2_ASAP7_75t_R FILLER_204_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_847 ();
 DECAPx1_ASAP7_75t_R FILLER_204_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_855 ();
 DECAPx6_ASAP7_75t_R FILLER_204_862 ();
 FILLER_ASAP7_75t_R FILLER_204_886 ();
 FILLER_ASAP7_75t_R FILLER_204_899 ();
 DECAPx10_ASAP7_75t_R FILLER_204_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_934 ();
 DECAPx4_ASAP7_75t_R FILLER_204_943 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_953 ();
 FILLER_ASAP7_75t_R FILLER_204_964 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_972 ();
 DECAPx4_ASAP7_75t_R FILLER_204_983 ();
 DECAPx6_ASAP7_75t_R FILLER_204_1003 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1048 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1063 ();
 DECAPx4_ASAP7_75t_R FILLER_204_1072 ();
 DECAPx4_ASAP7_75t_R FILLER_204_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1098 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_204_1113 ();
 FILLER_ASAP7_75t_R FILLER_204_1125 ();
 FILLER_ASAP7_75t_R FILLER_204_1134 ();
 FILLER_ASAP7_75t_R FILLER_204_1143 ();
 DECAPx2_ASAP7_75t_R FILLER_204_1152 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_204_1341 ();
 DECAPx6_ASAP7_75t_R FILLER_204_1363 ();
 FILLER_ASAP7_75t_R FILLER_205_2 ();
 FILLER_ASAP7_75t_R FILLER_205_30 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_35 ();
 DECAPx2_ASAP7_75t_R FILLER_205_44 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_50 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_59 ();
 DECAPx6_ASAP7_75t_R FILLER_205_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_82 ();
 DECAPx6_ASAP7_75t_R FILLER_205_91 ();
 DECAPx2_ASAP7_75t_R FILLER_205_105 ();
 FILLER_ASAP7_75t_R FILLER_205_117 ();
 FILLER_ASAP7_75t_R FILLER_205_125 ();
 FILLER_ASAP7_75t_R FILLER_205_133 ();
 DECAPx2_ASAP7_75t_R FILLER_205_143 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_149 ();
 DECAPx4_ASAP7_75t_R FILLER_205_159 ();
 FILLER_ASAP7_75t_R FILLER_205_175 ();
 DECAPx4_ASAP7_75t_R FILLER_205_180 ();
 DECAPx6_ASAP7_75t_R FILLER_205_196 ();
 FILLER_ASAP7_75t_R FILLER_205_210 ();
 DECAPx2_ASAP7_75t_R FILLER_205_218 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_224 ();
 FILLER_ASAP7_75t_R FILLER_205_233 ();
 FILLER_ASAP7_75t_R FILLER_205_241 ();
 DECAPx2_ASAP7_75t_R FILLER_205_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_252 ();
 DECAPx2_ASAP7_75t_R FILLER_205_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_262 ();
 DECAPx10_ASAP7_75t_R FILLER_205_269 ();
 DECAPx4_ASAP7_75t_R FILLER_205_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_301 ();
 DECAPx6_ASAP7_75t_R FILLER_205_305 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_319 ();
 DECAPx2_ASAP7_75t_R FILLER_205_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_334 ();
 DECAPx4_ASAP7_75t_R FILLER_205_338 ();
 FILLER_ASAP7_75t_R FILLER_205_348 ();
 DECAPx4_ASAP7_75t_R FILLER_205_358 ();
 FILLER_ASAP7_75t_R FILLER_205_368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_376 ();
 FILLER_ASAP7_75t_R FILLER_205_382 ();
 FILLER_ASAP7_75t_R FILLER_205_387 ();
 DECAPx2_ASAP7_75t_R FILLER_205_395 ();
 FILLER_ASAP7_75t_R FILLER_205_401 ();
 DECAPx4_ASAP7_75t_R FILLER_205_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_439 ();
 DECAPx6_ASAP7_75t_R FILLER_205_446 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_460 ();
 DECAPx6_ASAP7_75t_R FILLER_205_466 ();
 DECAPx2_ASAP7_75t_R FILLER_205_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_486 ();
 DECAPx1_ASAP7_75t_R FILLER_205_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_497 ();
 DECAPx10_ASAP7_75t_R FILLER_205_501 ();
 DECAPx2_ASAP7_75t_R FILLER_205_523 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_529 ();
 FILLER_ASAP7_75t_R FILLER_205_535 ();
 DECAPx4_ASAP7_75t_R FILLER_205_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_550 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_559 ();
 FILLER_ASAP7_75t_R FILLER_205_568 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_578 ();
 DECAPx1_ASAP7_75t_R FILLER_205_607 ();
 DECAPx2_ASAP7_75t_R FILLER_205_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_620 ();
 DECAPx4_ASAP7_75t_R FILLER_205_629 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_639 ();
 DECAPx6_ASAP7_75t_R FILLER_205_650 ();
 DECAPx1_ASAP7_75t_R FILLER_205_664 ();
 DECAPx6_ASAP7_75t_R FILLER_205_674 ();
 FILLER_ASAP7_75t_R FILLER_205_688 ();
 DECAPx2_ASAP7_75t_R FILLER_205_697 ();
 FILLER_ASAP7_75t_R FILLER_205_709 ();
 DECAPx2_ASAP7_75t_R FILLER_205_715 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_721 ();
 DECAPx2_ASAP7_75t_R FILLER_205_728 ();
 FILLER_ASAP7_75t_R FILLER_205_734 ();
 DECAPx2_ASAP7_75t_R FILLER_205_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_748 ();
 DECAPx6_ASAP7_75t_R FILLER_205_752 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_766 ();
 FILLER_ASAP7_75t_R FILLER_205_775 ();
 DECAPx4_ASAP7_75t_R FILLER_205_783 ();
 FILLER_ASAP7_75t_R FILLER_205_793 ();
 DECAPx2_ASAP7_75t_R FILLER_205_801 ();
 FILLER_ASAP7_75t_R FILLER_205_807 ();
 DECAPx10_ASAP7_75t_R FILLER_205_816 ();
 DECAPx10_ASAP7_75t_R FILLER_205_838 ();
 DECAPx4_ASAP7_75t_R FILLER_205_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_870 ();
 DECAPx6_ASAP7_75t_R FILLER_205_877 ();
 FILLER_ASAP7_75t_R FILLER_205_891 ();
 FILLER_ASAP7_75t_R FILLER_205_896 ();
 DECAPx4_ASAP7_75t_R FILLER_205_901 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_911 ();
 DECAPx1_ASAP7_75t_R FILLER_205_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_924 ();
 DECAPx2_ASAP7_75t_R FILLER_205_927 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_933 ();
 DECAPx4_ASAP7_75t_R FILLER_205_942 ();
 FILLER_ASAP7_75t_R FILLER_205_952 ();
 FILLER_ASAP7_75t_R FILLER_205_960 ();
 DECAPx1_ASAP7_75t_R FILLER_205_965 ();
 DECAPx4_ASAP7_75t_R FILLER_205_977 ();
 FILLER_ASAP7_75t_R FILLER_205_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1022 ();
 DECAPx6_ASAP7_75t_R FILLER_205_1044 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_1058 ();
 DECAPx4_ASAP7_75t_R FILLER_205_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1078 ();
 FILLER_ASAP7_75t_R FILLER_205_1105 ();
 DECAPx2_ASAP7_75t_R FILLER_205_1133 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_205_1344 ();
 DECAPx4_ASAP7_75t_R FILLER_205_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_206_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_16 ();
 DECAPx1_ASAP7_75t_R FILLER_206_20 ();
 DECAPx2_ASAP7_75t_R FILLER_206_50 ();
 DECAPx2_ASAP7_75t_R FILLER_206_64 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_70 ();
 DECAPx2_ASAP7_75t_R FILLER_206_99 ();
 FILLER_ASAP7_75t_R FILLER_206_105 ();
 DECAPx2_ASAP7_75t_R FILLER_206_113 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_119 ();
 FILLER_ASAP7_75t_R FILLER_206_125 ();
 FILLER_ASAP7_75t_R FILLER_206_133 ();
 DECAPx2_ASAP7_75t_R FILLER_206_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_149 ();
 DECAPx2_ASAP7_75t_R FILLER_206_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_163 ();
 DECAPx6_ASAP7_75t_R FILLER_206_190 ();
 FILLER_ASAP7_75t_R FILLER_206_204 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_209 ();
 DECAPx2_ASAP7_75t_R FILLER_206_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_224 ();
 DECAPx2_ASAP7_75t_R FILLER_206_251 ();
 FILLER_ASAP7_75t_R FILLER_206_257 ();
 FILLER_ASAP7_75t_R FILLER_206_267 ();
 DECAPx2_ASAP7_75t_R FILLER_206_275 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_281 ();
 FILLER_ASAP7_75t_R FILLER_206_290 ();
 DECAPx10_ASAP7_75t_R FILLER_206_295 ();
 DECAPx2_ASAP7_75t_R FILLER_206_317 ();
 DECAPx10_ASAP7_75t_R FILLER_206_329 ();
 FILLER_ASAP7_75t_R FILLER_206_351 ();
 FILLER_ASAP7_75t_R FILLER_206_361 ();
 DECAPx2_ASAP7_75t_R FILLER_206_373 ();
 FILLER_ASAP7_75t_R FILLER_206_387 ();
 DECAPx4_ASAP7_75t_R FILLER_206_395 ();
 DECAPx2_ASAP7_75t_R FILLER_206_411 ();
 DECAPx4_ASAP7_75t_R FILLER_206_420 ();
 DECAPx2_ASAP7_75t_R FILLER_206_456 ();
 DECAPx2_ASAP7_75t_R FILLER_206_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_470 ();
 DECAPx6_ASAP7_75t_R FILLER_206_483 ();
 DECAPx2_ASAP7_75t_R FILLER_206_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_503 ();
 FILLER_ASAP7_75t_R FILLER_206_510 ();
 DECAPx1_ASAP7_75t_R FILLER_206_518 ();
 FILLER_ASAP7_75t_R FILLER_206_529 ();
 DECAPx1_ASAP7_75t_R FILLER_206_537 ();
 FILLER_ASAP7_75t_R FILLER_206_544 ();
 FILLER_ASAP7_75t_R FILLER_206_552 ();
 DECAPx4_ASAP7_75t_R FILLER_206_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_572 ();
 FILLER_ASAP7_75t_R FILLER_206_579 ();
 FILLER_ASAP7_75t_R FILLER_206_587 ();
 FILLER_ASAP7_75t_R FILLER_206_595 ();
 FILLER_ASAP7_75t_R FILLER_206_623 ();
 DECAPx1_ASAP7_75t_R FILLER_206_633 ();
 FILLER_ASAP7_75t_R FILLER_206_640 ();
 DECAPx4_ASAP7_75t_R FILLER_206_648 ();
 FILLER_ASAP7_75t_R FILLER_206_658 ();
 DECAPx1_ASAP7_75t_R FILLER_206_666 ();
 DECAPx4_ASAP7_75t_R FILLER_206_677 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_687 ();
 DECAPx1_ASAP7_75t_R FILLER_206_696 ();
 FILLER_ASAP7_75t_R FILLER_206_726 ();
 DECAPx4_ASAP7_75t_R FILLER_206_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_741 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_752 ();
 FILLER_ASAP7_75t_R FILLER_206_764 ();
 DECAPx6_ASAP7_75t_R FILLER_206_769 ();
 DECAPx1_ASAP7_75t_R FILLER_206_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_787 ();
 FILLER_ASAP7_75t_R FILLER_206_794 ();
 DECAPx2_ASAP7_75t_R FILLER_206_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_808 ();
 FILLER_ASAP7_75t_R FILLER_206_815 ();
 DECAPx2_ASAP7_75t_R FILLER_206_824 ();
 FILLER_ASAP7_75t_R FILLER_206_840 ();
 DECAPx6_ASAP7_75t_R FILLER_206_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_865 ();
 FILLER_ASAP7_75t_R FILLER_206_872 ();
 FILLER_ASAP7_75t_R FILLER_206_880 ();
 FILLER_ASAP7_75t_R FILLER_206_888 ();
 DECAPx1_ASAP7_75t_R FILLER_206_900 ();
 FILLER_ASAP7_75t_R FILLER_206_912 ();
 FILLER_ASAP7_75t_R FILLER_206_940 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_950 ();
 DECAPx2_ASAP7_75t_R FILLER_206_961 ();
 FILLER_ASAP7_75t_R FILLER_206_967 ();
 FILLER_ASAP7_75t_R FILLER_206_975 ();
 DECAPx1_ASAP7_75t_R FILLER_206_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_987 ();
 FILLER_ASAP7_75t_R FILLER_206_994 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_999 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1005 ();
 FILLER_ASAP7_75t_R FILLER_206_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1053 ();
 FILLER_ASAP7_75t_R FILLER_206_1064 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1114 ();
 DECAPx4_ASAP7_75t_R FILLER_206_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1128 ();
 FILLER_ASAP7_75t_R FILLER_206_1135 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1144 ();
 DECAPx2_ASAP7_75t_R FILLER_206_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_206_1336 ();
 DECAPx6_ASAP7_75t_R FILLER_206_1358 ();
 DECAPx1_ASAP7_75t_R FILLER_206_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_207_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_8 ();
 FILLER_ASAP7_75t_R FILLER_207_17 ();
 DECAPx4_ASAP7_75t_R FILLER_207_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_32 ();
 FILLER_ASAP7_75t_R FILLER_207_39 ();
 DECAPx4_ASAP7_75t_R FILLER_207_44 ();
 DECAPx6_ASAP7_75t_R FILLER_207_62 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_76 ();
 DECAPx1_ASAP7_75t_R FILLER_207_85 ();
 DECAPx1_ASAP7_75t_R FILLER_207_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_96 ();
 FILLER_ASAP7_75t_R FILLER_207_123 ();
 DECAPx6_ASAP7_75t_R FILLER_207_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_142 ();
 FILLER_ASAP7_75t_R FILLER_207_149 ();
 DECAPx2_ASAP7_75t_R FILLER_207_157 ();
 FILLER_ASAP7_75t_R FILLER_207_163 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_171 ();
 FILLER_ASAP7_75t_R FILLER_207_177 ();
 DECAPx1_ASAP7_75t_R FILLER_207_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_209 ();
 DECAPx6_ASAP7_75t_R FILLER_207_216 ();
 DECAPx1_ASAP7_75t_R FILLER_207_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_234 ();
 FILLER_ASAP7_75t_R FILLER_207_241 ();
 DECAPx6_ASAP7_75t_R FILLER_207_246 ();
 DECAPx2_ASAP7_75t_R FILLER_207_268 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_274 ();
 FILLER_ASAP7_75t_R FILLER_207_303 ();
 DECAPx2_ASAP7_75t_R FILLER_207_308 ();
 FILLER_ASAP7_75t_R FILLER_207_340 ();
 DECAPx1_ASAP7_75t_R FILLER_207_345 ();
 FILLER_ASAP7_75t_R FILLER_207_355 ();
 DECAPx10_ASAP7_75t_R FILLER_207_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_401 ();
 DECAPx2_ASAP7_75t_R FILLER_207_408 ();
 DECAPx2_ASAP7_75t_R FILLER_207_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_426 ();
 FILLER_ASAP7_75t_R FILLER_207_433 ();
 DECAPx1_ASAP7_75t_R FILLER_207_441 ();
 DECAPx2_ASAP7_75t_R FILLER_207_448 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_454 ();
 FILLER_ASAP7_75t_R FILLER_207_460 ();
 DECAPx2_ASAP7_75t_R FILLER_207_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_475 ();
 DECAPx6_ASAP7_75t_R FILLER_207_482 ();
 DECAPx2_ASAP7_75t_R FILLER_207_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_502 ();
 DECAPx4_ASAP7_75t_R FILLER_207_509 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_519 ();
 DECAPx1_ASAP7_75t_R FILLER_207_548 ();
 DECAPx6_ASAP7_75t_R FILLER_207_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_572 ();
 DECAPx1_ASAP7_75t_R FILLER_207_579 ();
 DECAPx2_ASAP7_75t_R FILLER_207_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_595 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_599 ();
 DECAPx4_ASAP7_75t_R FILLER_207_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_618 ();
 FILLER_ASAP7_75t_R FILLER_207_625 ();
 DECAPx4_ASAP7_75t_R FILLER_207_633 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_643 ();
 DECAPx2_ASAP7_75t_R FILLER_207_653 ();
 FILLER_ASAP7_75t_R FILLER_207_659 ();
 FILLER_ASAP7_75t_R FILLER_207_668 ();
 DECAPx6_ASAP7_75t_R FILLER_207_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_690 ();
 DECAPx4_ASAP7_75t_R FILLER_207_698 ();
 DECAPx6_ASAP7_75t_R FILLER_207_734 ();
 DECAPx1_ASAP7_75t_R FILLER_207_748 ();
 DECAPx6_ASAP7_75t_R FILLER_207_755 ();
 FILLER_ASAP7_75t_R FILLER_207_769 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_780 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_789 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_798 ();
 FILLER_ASAP7_75t_R FILLER_207_807 ();
 DECAPx2_ASAP7_75t_R FILLER_207_817 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_823 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_852 ();
 FILLER_ASAP7_75t_R FILLER_207_862 ();
 FILLER_ASAP7_75t_R FILLER_207_870 ();
 DECAPx10_ASAP7_75t_R FILLER_207_878 ();
 DECAPx2_ASAP7_75t_R FILLER_207_906 ();
 FILLER_ASAP7_75t_R FILLER_207_912 ();
 DECAPx1_ASAP7_75t_R FILLER_207_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_924 ();
 FILLER_ASAP7_75t_R FILLER_207_927 ();
 DECAPx10_ASAP7_75t_R FILLER_207_932 ();
 DECAPx10_ASAP7_75t_R FILLER_207_954 ();
 DECAPx10_ASAP7_75t_R FILLER_207_976 ();
 DECAPx6_ASAP7_75t_R FILLER_207_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1016 ();
 FILLER_ASAP7_75t_R FILLER_207_1022 ();
 FILLER_ASAP7_75t_R FILLER_207_1027 ();
 DECAPx4_ASAP7_75t_R FILLER_207_1036 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1058 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1114 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_207_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_207_1369 ();
 FILLER_ASAP7_75t_R FILLER_207_1375 ();
 FILLER_ASAP7_75t_R FILLER_208_2 ();
 FILLER_ASAP7_75t_R FILLER_208_30 ();
 DECAPx10_ASAP7_75t_R FILLER_208_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_57 ();
 DECAPx10_ASAP7_75t_R FILLER_208_64 ();
 FILLER_ASAP7_75t_R FILLER_208_86 ();
 DECAPx4_ASAP7_75t_R FILLER_208_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_101 ();
 DECAPx1_ASAP7_75t_R FILLER_208_108 ();
 DECAPx10_ASAP7_75t_R FILLER_208_115 ();
 DECAPx2_ASAP7_75t_R FILLER_208_137 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_143 ();
 DECAPx10_ASAP7_75t_R FILLER_208_154 ();
 DECAPx1_ASAP7_75t_R FILLER_208_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_180 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_187 ();
 DECAPx1_ASAP7_75t_R FILLER_208_196 ();
 DECAPx6_ASAP7_75t_R FILLER_208_226 ();
 FILLER_ASAP7_75t_R FILLER_208_240 ();
 FILLER_ASAP7_75t_R FILLER_208_248 ();
 DECAPx10_ASAP7_75t_R FILLER_208_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_278 ();
 DECAPx10_ASAP7_75t_R FILLER_208_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_307 ();
 FILLER_ASAP7_75t_R FILLER_208_314 ();
 DECAPx2_ASAP7_75t_R FILLER_208_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_328 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_332 ();
 DECAPx2_ASAP7_75t_R FILLER_208_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_347 ();
 DECAPx10_ASAP7_75t_R FILLER_208_354 ();
 DECAPx1_ASAP7_75t_R FILLER_208_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_380 ();
 DECAPx4_ASAP7_75t_R FILLER_208_387 ();
 FILLER_ASAP7_75t_R FILLER_208_397 ();
 DECAPx1_ASAP7_75t_R FILLER_208_425 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_451 ();
 FILLER_ASAP7_75t_R FILLER_208_460 ();
 FILLER_ASAP7_75t_R FILLER_208_464 ();
 FILLER_ASAP7_75t_R FILLER_208_474 ();
 FILLER_ASAP7_75t_R FILLER_208_491 ();
 DECAPx2_ASAP7_75t_R FILLER_208_499 ();
 DECAPx4_ASAP7_75t_R FILLER_208_513 ();
 FILLER_ASAP7_75t_R FILLER_208_523 ();
 DECAPx1_ASAP7_75t_R FILLER_208_531 ();
 DECAPx1_ASAP7_75t_R FILLER_208_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_545 ();
 DECAPx10_ASAP7_75t_R FILLER_208_552 ();
 DECAPx6_ASAP7_75t_R FILLER_208_574 ();
 DECAPx2_ASAP7_75t_R FILLER_208_588 ();
 DECAPx6_ASAP7_75t_R FILLER_208_600 ();
 FILLER_ASAP7_75t_R FILLER_208_614 ();
 DECAPx6_ASAP7_75t_R FILLER_208_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_633 ();
 FILLER_ASAP7_75t_R FILLER_208_640 ();
 DECAPx2_ASAP7_75t_R FILLER_208_652 ();
 FILLER_ASAP7_75t_R FILLER_208_658 ();
 FILLER_ASAP7_75t_R FILLER_208_667 ();
 DECAPx2_ASAP7_75t_R FILLER_208_707 ();
 FILLER_ASAP7_75t_R FILLER_208_713 ();
 DECAPx2_ASAP7_75t_R FILLER_208_718 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_724 ();
 DECAPx6_ASAP7_75t_R FILLER_208_733 ();
 FILLER_ASAP7_75t_R FILLER_208_747 ();
 FILLER_ASAP7_75t_R FILLER_208_758 ();
 DECAPx2_ASAP7_75t_R FILLER_208_763 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_769 ();
 DECAPx10_ASAP7_75t_R FILLER_208_775 ();
 DECAPx6_ASAP7_75t_R FILLER_208_797 ();
 DECAPx1_ASAP7_75t_R FILLER_208_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_821 ();
 DECAPx2_ASAP7_75t_R FILLER_208_830 ();
 FILLER_ASAP7_75t_R FILLER_208_846 ();
 DECAPx4_ASAP7_75t_R FILLER_208_851 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_861 ();
 DECAPx4_ASAP7_75t_R FILLER_208_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_877 ();
 DECAPx10_ASAP7_75t_R FILLER_208_886 ();
 DECAPx2_ASAP7_75t_R FILLER_208_908 ();
 DECAPx1_ASAP7_75t_R FILLER_208_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_924 ();
 DECAPx4_ASAP7_75t_R FILLER_208_931 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_948 ();
 FILLER_ASAP7_75t_R FILLER_208_958 ();
 DECAPx1_ASAP7_75t_R FILLER_208_966 ();
 FILLER_ASAP7_75t_R FILLER_208_976 ();
 DECAPx4_ASAP7_75t_R FILLER_208_986 ();
 FILLER_ASAP7_75t_R FILLER_208_996 ();
 FILLER_ASAP7_75t_R FILLER_208_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_208_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_208_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_208_1084 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_208_1338 ();
 DECAPx6_ASAP7_75t_R FILLER_208_1360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_1374 ();
 DECAPx1_ASAP7_75t_R FILLER_209_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_6 ();
 DECAPx2_ASAP7_75t_R FILLER_209_13 ();
 FILLER_ASAP7_75t_R FILLER_209_19 ();
 DECAPx6_ASAP7_75t_R FILLER_209_27 ();
 DECAPx1_ASAP7_75t_R FILLER_209_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_45 ();
 FILLER_ASAP7_75t_R FILLER_209_54 ();
 FILLER_ASAP7_75t_R FILLER_209_64 ();
 DECAPx2_ASAP7_75t_R FILLER_209_72 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_78 ();
 DECAPx6_ASAP7_75t_R FILLER_209_87 ();
 FILLER_ASAP7_75t_R FILLER_209_127 ();
 DECAPx4_ASAP7_75t_R FILLER_209_135 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_145 ();
 DECAPx2_ASAP7_75t_R FILLER_209_156 ();
 FILLER_ASAP7_75t_R FILLER_209_162 ();
 DECAPx10_ASAP7_75t_R FILLER_209_170 ();
 FILLER_ASAP7_75t_R FILLER_209_192 ();
 DECAPx2_ASAP7_75t_R FILLER_209_197 ();
 DECAPx2_ASAP7_75t_R FILLER_209_209 ();
 DECAPx6_ASAP7_75t_R FILLER_209_218 ();
 DECAPx2_ASAP7_75t_R FILLER_209_238 ();
 FILLER_ASAP7_75t_R FILLER_209_250 ();
 FILLER_ASAP7_75t_R FILLER_209_258 ();
 DECAPx4_ASAP7_75t_R FILLER_209_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_276 ();
 DECAPx6_ASAP7_75t_R FILLER_209_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_299 ();
 DECAPx1_ASAP7_75t_R FILLER_209_308 ();
 FILLER_ASAP7_75t_R FILLER_209_320 ();
 DECAPx1_ASAP7_75t_R FILLER_209_329 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_359 ();
 FILLER_ASAP7_75t_R FILLER_209_370 ();
 FILLER_ASAP7_75t_R FILLER_209_398 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_410 ();
 DECAPx6_ASAP7_75t_R FILLER_209_416 ();
 FILLER_ASAP7_75t_R FILLER_209_430 ();
 FILLER_ASAP7_75t_R FILLER_209_458 ();
 DECAPx6_ASAP7_75t_R FILLER_209_466 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_480 ();
 FILLER_ASAP7_75t_R FILLER_209_509 ();
 DECAPx6_ASAP7_75t_R FILLER_209_517 ();
 FILLER_ASAP7_75t_R FILLER_209_531 ();
 DECAPx2_ASAP7_75t_R FILLER_209_559 ();
 FILLER_ASAP7_75t_R FILLER_209_565 ();
 FILLER_ASAP7_75t_R FILLER_209_573 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_578 ();
 DECAPx2_ASAP7_75t_R FILLER_209_587 ();
 FILLER_ASAP7_75t_R FILLER_209_593 ();
 FILLER_ASAP7_75t_R FILLER_209_601 ();
 FILLER_ASAP7_75t_R FILLER_209_625 ();
 DECAPx4_ASAP7_75t_R FILLER_209_633 ();
 FILLER_ASAP7_75t_R FILLER_209_643 ();
 DECAPx4_ASAP7_75t_R FILLER_209_652 ();
 DECAPx1_ASAP7_75t_R FILLER_209_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_673 ();
 FILLER_ASAP7_75t_R FILLER_209_680 ();
 FILLER_ASAP7_75t_R FILLER_209_688 ();
 DECAPx4_ASAP7_75t_R FILLER_209_696 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_706 ();
 DECAPx4_ASAP7_75t_R FILLER_209_715 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_725 ();
 DECAPx1_ASAP7_75t_R FILLER_209_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_740 ();
 FILLER_ASAP7_75t_R FILLER_209_747 ();
 DECAPx6_ASAP7_75t_R FILLER_209_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_766 ();
 DECAPx2_ASAP7_75t_R FILLER_209_776 ();
 FILLER_ASAP7_75t_R FILLER_209_796 ();
 DECAPx10_ASAP7_75t_R FILLER_209_808 ();
 DECAPx6_ASAP7_75t_R FILLER_209_830 ();
 DECAPx2_ASAP7_75t_R FILLER_209_844 ();
 FILLER_ASAP7_75t_R FILLER_209_876 ();
 DECAPx2_ASAP7_75t_R FILLER_209_904 ();
 DECAPx4_ASAP7_75t_R FILLER_209_913 ();
 FILLER_ASAP7_75t_R FILLER_209_923 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_927 ();
 FILLER_ASAP7_75t_R FILLER_209_936 ();
 FILLER_ASAP7_75t_R FILLER_209_946 ();
 FILLER_ASAP7_75t_R FILLER_209_960 ();
 DECAPx2_ASAP7_75t_R FILLER_209_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_976 ();
 FILLER_ASAP7_75t_R FILLER_209_1003 ();
 FILLER_ASAP7_75t_R FILLER_209_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_209_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1056 ();
 DECAPx6_ASAP7_75t_R FILLER_209_1078 ();
 FILLER_ASAP7_75t_R FILLER_209_1092 ();
 FILLER_ASAP7_75t_R FILLER_209_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1142 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_209_1340 ();
 DECAPx6_ASAP7_75t_R FILLER_209_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_210_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_16 ();
 FILLER_ASAP7_75t_R FILLER_210_43 ();
 DECAPx6_ASAP7_75t_R FILLER_210_51 ();
 DECAPx1_ASAP7_75t_R FILLER_210_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_69 ();
 FILLER_ASAP7_75t_R FILLER_210_96 ();
 FILLER_ASAP7_75t_R FILLER_210_108 ();
 DECAPx1_ASAP7_75t_R FILLER_210_116 ();
 FILLER_ASAP7_75t_R FILLER_210_146 ();
 FILLER_ASAP7_75t_R FILLER_210_154 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_159 ();
 DECAPx10_ASAP7_75t_R FILLER_210_188 ();
 DECAPx2_ASAP7_75t_R FILLER_210_210 ();
 FILLER_ASAP7_75t_R FILLER_210_216 ();
 DECAPx2_ASAP7_75t_R FILLER_210_244 ();
 DECAPx6_ASAP7_75t_R FILLER_210_256 ();
 FILLER_ASAP7_75t_R FILLER_210_270 ();
 FILLER_ASAP7_75t_R FILLER_210_298 ();
 FILLER_ASAP7_75t_R FILLER_210_308 ();
 DECAPx10_ASAP7_75t_R FILLER_210_313 ();
 DECAPx2_ASAP7_75t_R FILLER_210_335 ();
 FILLER_ASAP7_75t_R FILLER_210_341 ();
 FILLER_ASAP7_75t_R FILLER_210_349 ();
 DECAPx1_ASAP7_75t_R FILLER_210_354 ();
 FILLER_ASAP7_75t_R FILLER_210_380 ();
 FILLER_ASAP7_75t_R FILLER_210_388 ();
 DECAPx2_ASAP7_75t_R FILLER_210_393 ();
 DECAPx2_ASAP7_75t_R FILLER_210_405 ();
 FILLER_ASAP7_75t_R FILLER_210_411 ();
 DECAPx2_ASAP7_75t_R FILLER_210_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_425 ();
 FILLER_ASAP7_75t_R FILLER_210_444 ();
 FILLER_ASAP7_75t_R FILLER_210_452 ();
 DECAPx1_ASAP7_75t_R FILLER_210_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_461 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_464 ();
 DECAPx6_ASAP7_75t_R FILLER_210_473 ();
 DECAPx1_ASAP7_75t_R FILLER_210_487 ();
 FILLER_ASAP7_75t_R FILLER_210_497 ();
 DECAPx2_ASAP7_75t_R FILLER_210_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_508 ();
 FILLER_ASAP7_75t_R FILLER_210_517 ();
 DECAPx10_ASAP7_75t_R FILLER_210_525 ();
 DECAPx4_ASAP7_75t_R FILLER_210_550 ();
 DECAPx1_ASAP7_75t_R FILLER_210_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_590 ();
 FILLER_ASAP7_75t_R FILLER_210_617 ();
 FILLER_ASAP7_75t_R FILLER_210_645 ();
 DECAPx10_ASAP7_75t_R FILLER_210_654 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_676 ();
 DECAPx1_ASAP7_75t_R FILLER_210_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_697 ();
 FILLER_ASAP7_75t_R FILLER_210_704 ();
 DECAPx6_ASAP7_75t_R FILLER_210_720 ();
 FILLER_ASAP7_75t_R FILLER_210_734 ();
 FILLER_ASAP7_75t_R FILLER_210_742 ();
 DECAPx4_ASAP7_75t_R FILLER_210_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_763 ();
 FILLER_ASAP7_75t_R FILLER_210_774 ();
 DECAPx6_ASAP7_75t_R FILLER_210_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_793 ();
 DECAPx1_ASAP7_75t_R FILLER_210_797 ();
 DECAPx1_ASAP7_75t_R FILLER_210_811 ();
 DECAPx1_ASAP7_75t_R FILLER_210_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_825 ();
 DECAPx2_ASAP7_75t_R FILLER_210_835 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_841 ();
 DECAPx10_ASAP7_75t_R FILLER_210_851 ();
 DECAPx6_ASAP7_75t_R FILLER_210_873 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_887 ();
 FILLER_ASAP7_75t_R FILLER_210_893 ();
 DECAPx2_ASAP7_75t_R FILLER_210_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_927 ();
 DECAPx1_ASAP7_75t_R FILLER_210_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_938 ();
 FILLER_ASAP7_75t_R FILLER_210_965 ();
 FILLER_ASAP7_75t_R FILLER_210_993 ();
 DECAPx4_ASAP7_75t_R FILLER_210_998 ();
 FILLER_ASAP7_75t_R FILLER_210_1011 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_1020 ();
 DECAPx6_ASAP7_75t_R FILLER_210_1030 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_210_1061 ();
 FILLER_ASAP7_75t_R FILLER_210_1067 ();
 FILLER_ASAP7_75t_R FILLER_210_1081 ();
 FILLER_ASAP7_75t_R FILLER_210_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_210_1351 ();
 DECAPx1_ASAP7_75t_R FILLER_210_1373 ();
 DECAPx1_ASAP7_75t_R FILLER_211_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_6 ();
 DECAPx1_ASAP7_75t_R FILLER_211_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_17 ();
 DECAPx2_ASAP7_75t_R FILLER_211_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_30 ();
 DECAPx2_ASAP7_75t_R FILLER_211_34 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_40 ();
 DECAPx10_ASAP7_75t_R FILLER_211_49 ();
 DECAPx1_ASAP7_75t_R FILLER_211_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_75 ();
 FILLER_ASAP7_75t_R FILLER_211_82 ();
 FILLER_ASAP7_75t_R FILLER_211_87 ();
 DECAPx2_ASAP7_75t_R FILLER_211_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_98 ();
 FILLER_ASAP7_75t_R FILLER_211_102 ();
 DECAPx2_ASAP7_75t_R FILLER_211_110 ();
 DECAPx2_ASAP7_75t_R FILLER_211_119 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_125 ();
 FILLER_ASAP7_75t_R FILLER_211_134 ();
 DECAPx2_ASAP7_75t_R FILLER_211_139 ();
 FILLER_ASAP7_75t_R FILLER_211_145 ();
 DECAPx6_ASAP7_75t_R FILLER_211_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_167 ();
 FILLER_ASAP7_75t_R FILLER_211_174 ();
 DECAPx2_ASAP7_75t_R FILLER_211_179 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_185 ();
 FILLER_ASAP7_75t_R FILLER_211_191 ();
 DECAPx1_ASAP7_75t_R FILLER_211_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_203 ();
 DECAPx2_ASAP7_75t_R FILLER_211_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_216 ();
 FILLER_ASAP7_75t_R FILLER_211_223 ();
 FILLER_ASAP7_75t_R FILLER_211_231 ();
 DECAPx2_ASAP7_75t_R FILLER_211_236 ();
 FILLER_ASAP7_75t_R FILLER_211_242 ();
 DECAPx4_ASAP7_75t_R FILLER_211_247 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_257 ();
 DECAPx2_ASAP7_75t_R FILLER_211_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_272 ();
 DECAPx2_ASAP7_75t_R FILLER_211_281 ();
 DECAPx1_ASAP7_75t_R FILLER_211_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_294 ();
 DECAPx1_ASAP7_75t_R FILLER_211_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_305 ();
 DECAPx10_ASAP7_75t_R FILLER_211_314 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_336 ();
 DECAPx4_ASAP7_75t_R FILLER_211_345 ();
 FILLER_ASAP7_75t_R FILLER_211_361 ();
 FILLER_ASAP7_75t_R FILLER_211_369 ();
 DECAPx10_ASAP7_75t_R FILLER_211_377 ();
 DECAPx4_ASAP7_75t_R FILLER_211_399 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_409 ();
 FILLER_ASAP7_75t_R FILLER_211_420 ();
 DECAPx2_ASAP7_75t_R FILLER_211_428 ();
 FILLER_ASAP7_75t_R FILLER_211_434 ();
 DECAPx1_ASAP7_75t_R FILLER_211_442 ();
 DECAPx2_ASAP7_75t_R FILLER_211_452 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_458 ();
 DECAPx10_ASAP7_75t_R FILLER_211_487 ();
 DECAPx1_ASAP7_75t_R FILLER_211_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_513 ();
 DECAPx10_ASAP7_75t_R FILLER_211_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_562 ();
 DECAPx1_ASAP7_75t_R FILLER_211_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_573 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_577 ();
 DECAPx6_ASAP7_75t_R FILLER_211_590 ();
 FILLER_ASAP7_75t_R FILLER_211_604 ();
 DECAPx6_ASAP7_75t_R FILLER_211_609 ();
 DECAPx1_ASAP7_75t_R FILLER_211_629 ();
 DECAPx6_ASAP7_75t_R FILLER_211_636 ();
 DECAPx1_ASAP7_75t_R FILLER_211_650 ();
 DECAPx6_ASAP7_75t_R FILLER_211_660 ();
 FILLER_ASAP7_75t_R FILLER_211_674 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_679 ();
 DECAPx4_ASAP7_75t_R FILLER_211_688 ();
 DECAPx2_ASAP7_75t_R FILLER_211_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_707 ();
 DECAPx2_ASAP7_75t_R FILLER_211_714 ();
 FILLER_ASAP7_75t_R FILLER_211_720 ();
 DECAPx10_ASAP7_75t_R FILLER_211_725 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_747 ();
 DECAPx4_ASAP7_75t_R FILLER_211_753 ();
 FILLER_ASAP7_75t_R FILLER_211_763 ();
 FILLER_ASAP7_75t_R FILLER_211_774 ();
 DECAPx2_ASAP7_75t_R FILLER_211_779 ();
 DECAPx6_ASAP7_75t_R FILLER_211_794 ();
 FILLER_ASAP7_75t_R FILLER_211_808 ();
 FILLER_ASAP7_75t_R FILLER_211_816 ();
 DECAPx2_ASAP7_75t_R FILLER_211_832 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_850 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_860 ();
 FILLER_ASAP7_75t_R FILLER_211_873 ();
 FILLER_ASAP7_75t_R FILLER_211_885 ();
 FILLER_ASAP7_75t_R FILLER_211_897 ();
 DECAPx2_ASAP7_75t_R FILLER_211_909 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_922 ();
 FILLER_ASAP7_75t_R FILLER_211_927 ();
 DECAPx6_ASAP7_75t_R FILLER_211_935 ();
 DECAPx1_ASAP7_75t_R FILLER_211_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_953 ();
 DECAPx10_ASAP7_75t_R FILLER_211_957 ();
 DECAPx2_ASAP7_75t_R FILLER_211_986 ();
 DECAPx10_ASAP7_75t_R FILLER_211_995 ();
 DECAPx6_ASAP7_75t_R FILLER_211_1017 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_1031 ();
 FILLER_ASAP7_75t_R FILLER_211_1040 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_1056 ();
 DECAPx4_ASAP7_75t_R FILLER_211_1073 ();
 FILLER_ASAP7_75t_R FILLER_211_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_211_1342 ();
 DECAPx4_ASAP7_75t_R FILLER_211_1364 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_1374 ();
 FILLER_ASAP7_75t_R FILLER_212_2 ();
 DECAPx2_ASAP7_75t_R FILLER_212_30 ();
 FILLER_ASAP7_75t_R FILLER_212_36 ();
 DECAPx4_ASAP7_75t_R FILLER_212_46 ();
 DECAPx1_ASAP7_75t_R FILLER_212_62 ();
 DECAPx10_ASAP7_75t_R FILLER_212_72 ();
 DECAPx6_ASAP7_75t_R FILLER_212_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_108 ();
 DECAPx10_ASAP7_75t_R FILLER_212_115 ();
 DECAPx2_ASAP7_75t_R FILLER_212_137 ();
 FILLER_ASAP7_75t_R FILLER_212_143 ();
 DECAPx6_ASAP7_75t_R FILLER_212_151 ();
 FILLER_ASAP7_75t_R FILLER_212_165 ();
 FILLER_ASAP7_75t_R FILLER_212_173 ();
 DECAPx2_ASAP7_75t_R FILLER_212_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_187 ();
 FILLER_ASAP7_75t_R FILLER_212_194 ();
 DECAPx2_ASAP7_75t_R FILLER_212_204 ();
 FILLER_ASAP7_75t_R FILLER_212_210 ();
 DECAPx6_ASAP7_75t_R FILLER_212_238 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_212_252 ();
 DECAPx10_ASAP7_75t_R FILLER_212_281 ();
 DECAPx2_ASAP7_75t_R FILLER_212_303 ();
 DECAPx2_ASAP7_75t_R FILLER_212_315 ();
 FILLER_ASAP7_75t_R FILLER_212_321 ();
 FILLER_ASAP7_75t_R FILLER_212_329 ();
 FILLER_ASAP7_75t_R FILLER_212_357 ();
 FILLER_ASAP7_75t_R FILLER_212_367 ();
 DECAPx4_ASAP7_75t_R FILLER_212_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_385 ();
 FILLER_ASAP7_75t_R FILLER_212_392 ();
 DECAPx2_ASAP7_75t_R FILLER_212_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_406 ();
 DECAPx1_ASAP7_75t_R FILLER_212_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_414 ();
 FILLER_ASAP7_75t_R FILLER_212_423 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_212_431 ();
 FILLER_ASAP7_75t_R FILLER_212_460 ();
 DECAPx4_ASAP7_75t_R FILLER_212_464 ();
 FILLER_ASAP7_75t_R FILLER_212_474 ();
 FILLER_ASAP7_75t_R FILLER_212_482 ();
 DECAPx6_ASAP7_75t_R FILLER_212_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_501 ();
 FILLER_ASAP7_75t_R FILLER_212_508 ();
 DECAPx2_ASAP7_75t_R FILLER_212_513 ();
 DECAPx2_ASAP7_75t_R FILLER_212_525 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_212_531 ();
 DECAPx2_ASAP7_75t_R FILLER_212_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_566 ();
 DECAPx10_ASAP7_75t_R FILLER_212_573 ();
 DECAPx1_ASAP7_75t_R FILLER_212_595 ();
 DECAPx6_ASAP7_75t_R FILLER_212_605 ();
 DECAPx2_ASAP7_75t_R FILLER_212_619 ();
 FILLER_ASAP7_75t_R FILLER_212_631 ();
 DECAPx2_ASAP7_75t_R FILLER_212_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_642 ();
 FILLER_ASAP7_75t_R FILLER_212_649 ();
 FILLER_ASAP7_75t_R FILLER_212_665 ();
 DECAPx6_ASAP7_75t_R FILLER_212_670 ();
 DECAPx4_ASAP7_75t_R FILLER_212_690 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_212_700 ();
 DECAPx2_ASAP7_75t_R FILLER_212_717 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_212_726 ();
 FILLER_ASAP7_75t_R FILLER_212_735 ();
 DECAPx6_ASAP7_75t_R FILLER_212_743 ();
 DECAPx1_ASAP7_75t_R FILLER_212_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_761 ();
 DECAPx4_ASAP7_75t_R FILLER_212_765 ();
 FILLER_ASAP7_75t_R FILLER_212_775 ();
 DECAPx1_ASAP7_75t_R FILLER_212_787 ();
 DECAPx1_ASAP7_75t_R FILLER_212_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_798 ();
 DECAPx6_ASAP7_75t_R FILLER_212_805 ();
 DECAPx2_ASAP7_75t_R FILLER_212_819 ();
 DECAPx1_ASAP7_75t_R FILLER_212_828 ();
 DECAPx4_ASAP7_75t_R FILLER_212_839 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_212_849 ();
 DECAPx10_ASAP7_75t_R FILLER_212_858 ();
 DECAPx10_ASAP7_75t_R FILLER_212_880 ();
 DECAPx2_ASAP7_75t_R FILLER_212_902 ();
 FILLER_ASAP7_75t_R FILLER_212_908 ();
 DECAPx10_ASAP7_75t_R FILLER_212_913 ();
 DECAPx10_ASAP7_75t_R FILLER_212_935 ();
 DECAPx10_ASAP7_75t_R FILLER_212_957 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_212_979 ();
 DECAPx10_ASAP7_75t_R FILLER_212_985 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1022 ();
 FILLER_ASAP7_75t_R FILLER_212_1030 ();
 DECAPx4_ASAP7_75t_R FILLER_212_1046 ();
 FILLER_ASAP7_75t_R FILLER_212_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_212_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_1076 ();
 FILLER_ASAP7_75t_R FILLER_212_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_212_1338 ();
 DECAPx6_ASAP7_75t_R FILLER_212_1360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_212_1374 ();
 DECAPx4_ASAP7_75t_R FILLER_213_2 ();
 FILLER_ASAP7_75t_R FILLER_213_18 ();
 DECAPx2_ASAP7_75t_R FILLER_213_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_29 ();
 DECAPx1_ASAP7_75t_R FILLER_213_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_37 ();
 DECAPx1_ASAP7_75t_R FILLER_213_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_50 ();
 FILLER_ASAP7_75t_R FILLER_213_59 ();
 FILLER_ASAP7_75t_R FILLER_213_69 ();
 DECAPx2_ASAP7_75t_R FILLER_213_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_83 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_213_91 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_213_100 ();
 FILLER_ASAP7_75t_R FILLER_213_129 ();
 DECAPx2_ASAP7_75t_R FILLER_213_157 ();
 FILLER_ASAP7_75t_R FILLER_213_163 ();
 DECAPx1_ASAP7_75t_R FILLER_213_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_195 ();
 DECAPx4_ASAP7_75t_R FILLER_213_204 ();
 DECAPx2_ASAP7_75t_R FILLER_213_220 ();
 DECAPx1_ASAP7_75t_R FILLER_213_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_233 ();
 DECAPx6_ASAP7_75t_R FILLER_213_237 ();
 FILLER_ASAP7_75t_R FILLER_213_251 ();
 FILLER_ASAP7_75t_R FILLER_213_256 ();
 DECAPx2_ASAP7_75t_R FILLER_213_264 ();
 DECAPx4_ASAP7_75t_R FILLER_213_273 ();
 FILLER_ASAP7_75t_R FILLER_213_283 ();
 DECAPx2_ASAP7_75t_R FILLER_213_291 ();
 DECAPx1_ASAP7_75t_R FILLER_213_303 ();
 FILLER_ASAP7_75t_R FILLER_213_313 ();
 DECAPx2_ASAP7_75t_R FILLER_213_341 ();
 FILLER_ASAP7_75t_R FILLER_213_369 ();
 DECAPx1_ASAP7_75t_R FILLER_213_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_383 ();
 DECAPx1_ASAP7_75t_R FILLER_213_410 ();
 FILLER_ASAP7_75t_R FILLER_213_420 ();
 FILLER_ASAP7_75t_R FILLER_213_428 ();
 DECAPx2_ASAP7_75t_R FILLER_213_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_442 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_213_449 ();
 DECAPx2_ASAP7_75t_R FILLER_213_455 ();
 DECAPx6_ASAP7_75t_R FILLER_213_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_213_478 ();
 DECAPx1_ASAP7_75t_R FILLER_213_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_488 ();
 DECAPx2_ASAP7_75t_R FILLER_213_515 ();
 FILLER_ASAP7_75t_R FILLER_213_521 ();
 FILLER_ASAP7_75t_R FILLER_213_529 ();
 DECAPx2_ASAP7_75t_R FILLER_213_534 ();
 FILLER_ASAP7_75t_R FILLER_213_546 ();
 FILLER_ASAP7_75t_R FILLER_213_554 ();
 DECAPx4_ASAP7_75t_R FILLER_213_559 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_213_575 ();
 DECAPx2_ASAP7_75t_R FILLER_213_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_587 ();
 DECAPx1_ASAP7_75t_R FILLER_213_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_618 ();
 DECAPx2_ASAP7_75t_R FILLER_213_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_651 ();
 FILLER_ASAP7_75t_R FILLER_213_658 ();
 FILLER_ASAP7_75t_R FILLER_213_663 ();
 FILLER_ASAP7_75t_R FILLER_213_679 ();
 DECAPx2_ASAP7_75t_R FILLER_213_695 ();
 DECAPx6_ASAP7_75t_R FILLER_213_710 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_213_724 ();
 DECAPx6_ASAP7_75t_R FILLER_213_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_755 ();
 DECAPx10_ASAP7_75t_R FILLER_213_765 ();
 DECAPx2_ASAP7_75t_R FILLER_213_787 ();
 FILLER_ASAP7_75t_R FILLER_213_802 ();
 DECAPx6_ASAP7_75t_R FILLER_213_813 ();
 DECAPx4_ASAP7_75t_R FILLER_213_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_840 ();
 DECAPx2_ASAP7_75t_R FILLER_213_848 ();
 FILLER_ASAP7_75t_R FILLER_213_861 ();
 DECAPx6_ASAP7_75t_R FILLER_213_873 ();
 DECAPx2_ASAP7_75t_R FILLER_213_887 ();
 DECAPx4_ASAP7_75t_R FILLER_213_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_913 ();
 DECAPx1_ASAP7_75t_R FILLER_213_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_924 ();
 FILLER_ASAP7_75t_R FILLER_213_927 ();
 FILLER_ASAP7_75t_R FILLER_213_935 ();
 DECAPx2_ASAP7_75t_R FILLER_213_944 ();
 FILLER_ASAP7_75t_R FILLER_213_950 ();
 DECAPx1_ASAP7_75t_R FILLER_213_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_963 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_213_970 ();
 FILLER_ASAP7_75t_R FILLER_213_980 ();
 FILLER_ASAP7_75t_R FILLER_213_989 ();
 FILLER_ASAP7_75t_R FILLER_213_998 ();
 FILLER_ASAP7_75t_R FILLER_213_1007 ();
 DECAPx6_ASAP7_75t_R FILLER_213_1016 ();
 FILLER_ASAP7_75t_R FILLER_213_1030 ();
 FILLER_ASAP7_75t_R FILLER_213_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1046 ();
 DECAPx4_ASAP7_75t_R FILLER_213_1068 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_213_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_213_1084 ();
 FILLER_ASAP7_75t_R FILLER_213_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_213_1337 ();
 DECAPx6_ASAP7_75t_R FILLER_213_1359 ();
 DECAPx1_ASAP7_75t_R FILLER_213_1373 ();
 DECAPx10_ASAP7_75t_R FILLER_214_2 ();
 DECAPx4_ASAP7_75t_R FILLER_214_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_34 ();
 FILLER_ASAP7_75t_R FILLER_214_41 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_49 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_55 ();
 DECAPx4_ASAP7_75t_R FILLER_214_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_74 ();
 FILLER_ASAP7_75t_R FILLER_214_81 ();
 DECAPx1_ASAP7_75t_R FILLER_214_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_95 ();
 FILLER_ASAP7_75t_R FILLER_214_106 ();
 DECAPx2_ASAP7_75t_R FILLER_214_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_120 ();
 DECAPx6_ASAP7_75t_R FILLER_214_124 ();
 FILLER_ASAP7_75t_R FILLER_214_144 ();
 DECAPx10_ASAP7_75t_R FILLER_214_149 ();
 DECAPx2_ASAP7_75t_R FILLER_214_171 ();
 FILLER_ASAP7_75t_R FILLER_214_177 ();
 DECAPx10_ASAP7_75t_R FILLER_214_182 ();
 DECAPx10_ASAP7_75t_R FILLER_214_204 ();
 DECAPx1_ASAP7_75t_R FILLER_214_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_230 ();
 FILLER_ASAP7_75t_R FILLER_214_237 ();
 DECAPx2_ASAP7_75t_R FILLER_214_247 ();
 DECAPx6_ASAP7_75t_R FILLER_214_259 ();
 DECAPx1_ASAP7_75t_R FILLER_214_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_277 ();
 DECAPx2_ASAP7_75t_R FILLER_214_304 ();
 FILLER_ASAP7_75t_R FILLER_214_316 ();
 DECAPx2_ASAP7_75t_R FILLER_214_324 ();
 DECAPx4_ASAP7_75t_R FILLER_214_333 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_343 ();
 DECAPx2_ASAP7_75t_R FILLER_214_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_355 ();
 FILLER_ASAP7_75t_R FILLER_214_378 ();
 DECAPx4_ASAP7_75t_R FILLER_214_386 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_396 ();
 DECAPx10_ASAP7_75t_R FILLER_214_402 ();
 DECAPx10_ASAP7_75t_R FILLER_214_424 ();
 DECAPx6_ASAP7_75t_R FILLER_214_446 ();
 FILLER_ASAP7_75t_R FILLER_214_460 ();
 FILLER_ASAP7_75t_R FILLER_214_464 ();
 DECAPx10_ASAP7_75t_R FILLER_214_473 ();
 FILLER_ASAP7_75t_R FILLER_214_501 ();
 DECAPx10_ASAP7_75t_R FILLER_214_506 ();
 DECAPx10_ASAP7_75t_R FILLER_214_528 ();
 DECAPx1_ASAP7_75t_R FILLER_214_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_562 ();
 DECAPx1_ASAP7_75t_R FILLER_214_589 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_599 ();
 FILLER_ASAP7_75t_R FILLER_214_605 ();
 DECAPx2_ASAP7_75t_R FILLER_214_613 ();
 FILLER_ASAP7_75t_R FILLER_214_619 ();
 DECAPx10_ASAP7_75t_R FILLER_214_627 ();
 DECAPx10_ASAP7_75t_R FILLER_214_649 ();
 DECAPx4_ASAP7_75t_R FILLER_214_671 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_681 ();
 DECAPx10_ASAP7_75t_R FILLER_214_690 ();
 DECAPx6_ASAP7_75t_R FILLER_214_712 ();
 DECAPx1_ASAP7_75t_R FILLER_214_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_730 ();
 DECAPx2_ASAP7_75t_R FILLER_214_737 ();
 DECAPx2_ASAP7_75t_R FILLER_214_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_752 ();
 FILLER_ASAP7_75t_R FILLER_214_759 ();
 FILLER_ASAP7_75t_R FILLER_214_767 ();
 DECAPx2_ASAP7_75t_R FILLER_214_772 ();
 FILLER_ASAP7_75t_R FILLER_214_778 ();
 FILLER_ASAP7_75t_R FILLER_214_789 ();
 DECAPx2_ASAP7_75t_R FILLER_214_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_800 ();
 DECAPx2_ASAP7_75t_R FILLER_214_804 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_810 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_816 ();
 DECAPx2_ASAP7_75t_R FILLER_214_828 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_834 ();
 DECAPx2_ASAP7_75t_R FILLER_214_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_852 ();
 DECAPx4_ASAP7_75t_R FILLER_214_863 ();
 FILLER_ASAP7_75t_R FILLER_214_873 ();
 FILLER_ASAP7_75t_R FILLER_214_885 ();
 FILLER_ASAP7_75t_R FILLER_214_897 ();
 DECAPx2_ASAP7_75t_R FILLER_214_909 ();
 FILLER_ASAP7_75t_R FILLER_214_915 ();
 DECAPx2_ASAP7_75t_R FILLER_214_924 ();
 DECAPx2_ASAP7_75t_R FILLER_214_936 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_942 ();
 DECAPx2_ASAP7_75t_R FILLER_214_951 ();
 FILLER_ASAP7_75t_R FILLER_214_957 ();
 FILLER_ASAP7_75t_R FILLER_214_966 ();
 DECAPx10_ASAP7_75t_R FILLER_214_975 ();
 DECAPx4_ASAP7_75t_R FILLER_214_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1007 ();
 FILLER_ASAP7_75t_R FILLER_214_1015 ();
 DECAPx6_ASAP7_75t_R FILLER_214_1024 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1044 ();
 DECAPx4_ASAP7_75t_R FILLER_214_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1058 ();
 FILLER_ASAP7_75t_R FILLER_214_1063 ();
 DECAPx4_ASAP7_75t_R FILLER_214_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_214_1346 ();
 DECAPx2_ASAP7_75t_R FILLER_214_1368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_1374 ();
 DECAPx4_ASAP7_75t_R FILLER_215_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_12 ();
 DECAPx10_ASAP7_75t_R FILLER_215_21 ();
 DECAPx2_ASAP7_75t_R FILLER_215_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_49 ();
 DECAPx2_ASAP7_75t_R FILLER_215_57 ();
 DECAPx4_ASAP7_75t_R FILLER_215_69 ();
 FILLER_ASAP7_75t_R FILLER_215_79 ();
 FILLER_ASAP7_75t_R FILLER_215_87 ();
 DECAPx6_ASAP7_75t_R FILLER_215_104 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_118 ();
 FILLER_ASAP7_75t_R FILLER_215_127 ();
 DECAPx6_ASAP7_75t_R FILLER_215_135 ();
 FILLER_ASAP7_75t_R FILLER_215_149 ();
 FILLER_ASAP7_75t_R FILLER_215_157 ();
 DECAPx4_ASAP7_75t_R FILLER_215_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_176 ();
 DECAPx2_ASAP7_75t_R FILLER_215_183 ();
 FILLER_ASAP7_75t_R FILLER_215_189 ();
 FILLER_ASAP7_75t_R FILLER_215_197 ();
 FILLER_ASAP7_75t_R FILLER_215_207 ();
 DECAPx1_ASAP7_75t_R FILLER_215_215 ();
 DECAPx4_ASAP7_75t_R FILLER_215_225 ();
 FILLER_ASAP7_75t_R FILLER_215_235 ();
 DECAPx1_ASAP7_75t_R FILLER_215_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_249 ();
 DECAPx2_ASAP7_75t_R FILLER_215_256 ();
 DECAPx4_ASAP7_75t_R FILLER_215_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_279 ();
 DECAPx2_ASAP7_75t_R FILLER_215_286 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_295 ();
 DECAPx10_ASAP7_75t_R FILLER_215_304 ();
 DECAPx4_ASAP7_75t_R FILLER_215_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_336 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_343 ();
 DECAPx1_ASAP7_75t_R FILLER_215_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_356 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_363 ();
 FILLER_ASAP7_75t_R FILLER_215_374 ();
 FILLER_ASAP7_75t_R FILLER_215_384 ();
 DECAPx2_ASAP7_75t_R FILLER_215_392 ();
 DECAPx2_ASAP7_75t_R FILLER_215_404 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_410 ();
 FILLER_ASAP7_75t_R FILLER_215_421 ();
 FILLER_ASAP7_75t_R FILLER_215_431 ();
 DECAPx1_ASAP7_75t_R FILLER_215_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_443 ();
 DECAPx2_ASAP7_75t_R FILLER_215_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_456 ();
 FILLER_ASAP7_75t_R FILLER_215_463 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_473 ();
 FILLER_ASAP7_75t_R FILLER_215_486 ();
 DECAPx10_ASAP7_75t_R FILLER_215_494 ();
 DECAPx4_ASAP7_75t_R FILLER_215_516 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_526 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_535 ();
 FILLER_ASAP7_75t_R FILLER_215_544 ();
 FILLER_ASAP7_75t_R FILLER_215_552 ();
 FILLER_ASAP7_75t_R FILLER_215_572 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_577 ();
 FILLER_ASAP7_75t_R FILLER_215_586 ();
 DECAPx2_ASAP7_75t_R FILLER_215_594 ();
 FILLER_ASAP7_75t_R FILLER_215_606 ();
 DECAPx6_ASAP7_75t_R FILLER_215_616 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_630 ();
 FILLER_ASAP7_75t_R FILLER_215_639 ();
 DECAPx2_ASAP7_75t_R FILLER_215_647 ();
 DECAPx10_ASAP7_75t_R FILLER_215_659 ();
 DECAPx10_ASAP7_75t_R FILLER_215_681 ();
 DECAPx2_ASAP7_75t_R FILLER_215_703 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_709 ();
 FILLER_ASAP7_75t_R FILLER_215_718 ();
 DECAPx10_ASAP7_75t_R FILLER_215_726 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_748 ();
 DECAPx6_ASAP7_75t_R FILLER_215_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_779 ();
 DECAPx10_ASAP7_75t_R FILLER_215_783 ();
 DECAPx2_ASAP7_75t_R FILLER_215_805 ();
 DECAPx6_ASAP7_75t_R FILLER_215_814 ();
 DECAPx1_ASAP7_75t_R FILLER_215_828 ();
 DECAPx2_ASAP7_75t_R FILLER_215_835 ();
 DECAPx10_ASAP7_75t_R FILLER_215_844 ();
 DECAPx2_ASAP7_75t_R FILLER_215_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_872 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_880 ();
 DECAPx6_ASAP7_75t_R FILLER_215_891 ();
 DECAPx1_ASAP7_75t_R FILLER_215_905 ();
 DECAPx4_ASAP7_75t_R FILLER_215_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_922 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_927 ();
 DECAPx2_ASAP7_75t_R FILLER_215_937 ();
 DECAPx10_ASAP7_75t_R FILLER_215_949 ();
 DECAPx6_ASAP7_75t_R FILLER_215_971 ();
 DECAPx1_ASAP7_75t_R FILLER_215_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_989 ();
 DECAPx6_ASAP7_75t_R FILLER_215_996 ();
 FILLER_ASAP7_75t_R FILLER_215_1016 ();
 DECAPx6_ASAP7_75t_R FILLER_215_1032 ();
 FILLER_ASAP7_75t_R FILLER_215_1060 ();
 DECAPx4_ASAP7_75t_R FILLER_215_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1075 ();
 DECAPx6_ASAP7_75t_R FILLER_215_1079 ();
 DECAPx1_ASAP7_75t_R FILLER_215_1093 ();
 FILLER_ASAP7_75t_R FILLER_215_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_215_1334 ();
 DECAPx6_ASAP7_75t_R FILLER_215_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_215_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_1376 ();
 DECAPx1_ASAP7_75t_R FILLER_216_2 ();
 DECAPx2_ASAP7_75t_R FILLER_216_32 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_38 ();
 DECAPx1_ASAP7_75t_R FILLER_216_47 ();
 DECAPx10_ASAP7_75t_R FILLER_216_77 ();
 FILLER_ASAP7_75t_R FILLER_216_105 ();
 FILLER_ASAP7_75t_R FILLER_216_114 ();
 DECAPx6_ASAP7_75t_R FILLER_216_142 ();
 FILLER_ASAP7_75t_R FILLER_216_156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_167 ();
 FILLER_ASAP7_75t_R FILLER_216_196 ();
 DECAPx1_ASAP7_75t_R FILLER_216_220 ();
 DECAPx1_ASAP7_75t_R FILLER_216_230 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_240 ();
 FILLER_ASAP7_75t_R FILLER_216_258 ();
 FILLER_ASAP7_75t_R FILLER_216_266 ();
 DECAPx10_ASAP7_75t_R FILLER_216_276 ();
 FILLER_ASAP7_75t_R FILLER_216_298 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_308 ();
 FILLER_ASAP7_75t_R FILLER_216_319 ();
 DECAPx2_ASAP7_75t_R FILLER_216_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_333 ();
 FILLER_ASAP7_75t_R FILLER_216_360 ();
 FILLER_ASAP7_75t_R FILLER_216_365 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_370 ();
 DECAPx2_ASAP7_75t_R FILLER_216_379 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_385 ();
 DECAPx2_ASAP7_75t_R FILLER_216_414 ();
 FILLER_ASAP7_75t_R FILLER_216_420 ();
 DECAPx1_ASAP7_75t_R FILLER_216_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_433 ();
 FILLER_ASAP7_75t_R FILLER_216_460 ();
 FILLER_ASAP7_75t_R FILLER_216_464 ();
 DECAPx2_ASAP7_75t_R FILLER_216_472 ();
 DECAPx2_ASAP7_75t_R FILLER_216_493 ();
 FILLER_ASAP7_75t_R FILLER_216_505 ();
 DECAPx2_ASAP7_75t_R FILLER_216_513 ();
 FILLER_ASAP7_75t_R FILLER_216_519 ();
 FILLER_ASAP7_75t_R FILLER_216_527 ();
 DECAPx1_ASAP7_75t_R FILLER_216_537 ();
 FILLER_ASAP7_75t_R FILLER_216_547 ();
 FILLER_ASAP7_75t_R FILLER_216_571 ();
 FILLER_ASAP7_75t_R FILLER_216_599 ();
 DECAPx1_ASAP7_75t_R FILLER_216_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_608 ();
 FILLER_ASAP7_75t_R FILLER_216_617 ();
 DECAPx2_ASAP7_75t_R FILLER_216_625 ();
 DECAPx2_ASAP7_75t_R FILLER_216_637 ();
 FILLER_ASAP7_75t_R FILLER_216_649 ();
 DECAPx4_ASAP7_75t_R FILLER_216_665 ();
 FILLER_ASAP7_75t_R FILLER_216_681 ();
 DECAPx2_ASAP7_75t_R FILLER_216_689 ();
 FILLER_ASAP7_75t_R FILLER_216_695 ();
 DECAPx2_ASAP7_75t_R FILLER_216_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_706 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_721 ();
 DECAPx6_ASAP7_75t_R FILLER_216_738 ();
 FILLER_ASAP7_75t_R FILLER_216_752 ();
 DECAPx6_ASAP7_75t_R FILLER_216_760 ();
 DECAPx4_ASAP7_75t_R FILLER_216_783 ();
 FILLER_ASAP7_75t_R FILLER_216_793 ();
 DECAPx6_ASAP7_75t_R FILLER_216_798 ();
 FILLER_ASAP7_75t_R FILLER_216_826 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_831 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_848 ();
 FILLER_ASAP7_75t_R FILLER_216_860 ();
 DECAPx10_ASAP7_75t_R FILLER_216_865 ();
 DECAPx6_ASAP7_75t_R FILLER_216_887 ();
 DECAPx1_ASAP7_75t_R FILLER_216_901 ();
 FILLER_ASAP7_75t_R FILLER_216_919 ();
 DECAPx4_ASAP7_75t_R FILLER_216_933 ();
 FILLER_ASAP7_75t_R FILLER_216_943 ();
 FILLER_ASAP7_75t_R FILLER_216_951 ();
 DECAPx4_ASAP7_75t_R FILLER_216_959 ();
 FILLER_ASAP7_75t_R FILLER_216_969 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_974 ();
 DECAPx2_ASAP7_75t_R FILLER_216_985 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_991 ();
 DECAPx4_ASAP7_75t_R FILLER_216_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1018 ();
 DECAPx6_ASAP7_75t_R FILLER_216_1025 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_1039 ();
 FILLER_ASAP7_75t_R FILLER_216_1045 ();
 DECAPx2_ASAP7_75t_R FILLER_216_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1060 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_1082 ();
 FILLER_ASAP7_75t_R FILLER_216_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_216_1353 ();
 FILLER_ASAP7_75t_R FILLER_216_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_217_2 ();
 FILLER_ASAP7_75t_R FILLER_217_8 ();
 DECAPx1_ASAP7_75t_R FILLER_217_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_20 ();
 DECAPx1_ASAP7_75t_R FILLER_217_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_28 ();
 FILLER_ASAP7_75t_R FILLER_217_55 ();
 FILLER_ASAP7_75t_R FILLER_217_64 ();
 FILLER_ASAP7_75t_R FILLER_217_73 ();
 FILLER_ASAP7_75t_R FILLER_217_81 ();
 DECAPx10_ASAP7_75t_R FILLER_217_86 ();
 DECAPx10_ASAP7_75t_R FILLER_217_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_130 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_134 ();
 FILLER_ASAP7_75t_R FILLER_217_140 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_150 ();
 DECAPx4_ASAP7_75t_R FILLER_217_159 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_169 ();
 DECAPx2_ASAP7_75t_R FILLER_217_178 ();
 DECAPx1_ASAP7_75t_R FILLER_217_187 ();
 FILLER_ASAP7_75t_R FILLER_217_197 ();
 DECAPx2_ASAP7_75t_R FILLER_217_207 ();
 FILLER_ASAP7_75t_R FILLER_217_213 ();
 DECAPx6_ASAP7_75t_R FILLER_217_241 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_255 ();
 DECAPx4_ASAP7_75t_R FILLER_217_266 ();
 FILLER_ASAP7_75t_R FILLER_217_282 ();
 DECAPx2_ASAP7_75t_R FILLER_217_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_296 ();
 DECAPx6_ASAP7_75t_R FILLER_217_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_314 ();
 FILLER_ASAP7_75t_R FILLER_217_321 ();
 DECAPx10_ASAP7_75t_R FILLER_217_329 ();
 FILLER_ASAP7_75t_R FILLER_217_351 ();
 DECAPx2_ASAP7_75t_R FILLER_217_359 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_365 ();
 DECAPx6_ASAP7_75t_R FILLER_217_371 ();
 DECAPx1_ASAP7_75t_R FILLER_217_385 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_398 ();
 FILLER_ASAP7_75t_R FILLER_217_404 ();
 FILLER_ASAP7_75t_R FILLER_217_412 ();
 FILLER_ASAP7_75t_R FILLER_217_420 ();
 FILLER_ASAP7_75t_R FILLER_217_429 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_438 ();
 DECAPx1_ASAP7_75t_R FILLER_217_447 ();
 DECAPx10_ASAP7_75t_R FILLER_217_454 ();
 DECAPx6_ASAP7_75t_R FILLER_217_476 ();
 DECAPx1_ASAP7_75t_R FILLER_217_490 ();
 FILLER_ASAP7_75t_R FILLER_217_520 ();
 FILLER_ASAP7_75t_R FILLER_217_530 ();
 FILLER_ASAP7_75t_R FILLER_217_535 ();
 DECAPx2_ASAP7_75t_R FILLER_217_543 ();
 FILLER_ASAP7_75t_R FILLER_217_549 ();
 DECAPx10_ASAP7_75t_R FILLER_217_559 ();
 DECAPx2_ASAP7_75t_R FILLER_217_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_587 ();
 DECAPx10_ASAP7_75t_R FILLER_217_591 ();
 FILLER_ASAP7_75t_R FILLER_217_613 ();
 DECAPx4_ASAP7_75t_R FILLER_217_621 ();
 DECAPx6_ASAP7_75t_R FILLER_217_637 ();
 FILLER_ASAP7_75t_R FILLER_217_651 ();
 DECAPx2_ASAP7_75t_R FILLER_217_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_665 ();
 FILLER_ASAP7_75t_R FILLER_217_669 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_685 ();
 DECAPx2_ASAP7_75t_R FILLER_217_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_708 ();
 DECAPx4_ASAP7_75t_R FILLER_217_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_725 ();
 FILLER_ASAP7_75t_R FILLER_217_729 ();
 FILLER_ASAP7_75t_R FILLER_217_740 ();
 DECAPx2_ASAP7_75t_R FILLER_217_745 ();
 DECAPx4_ASAP7_75t_R FILLER_217_757 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_767 ();
 FILLER_ASAP7_75t_R FILLER_217_784 ();
 FILLER_ASAP7_75t_R FILLER_217_792 ();
 DECAPx2_ASAP7_75t_R FILLER_217_797 ();
 FILLER_ASAP7_75t_R FILLER_217_812 ();
 DECAPx1_ASAP7_75t_R FILLER_217_817 ();
 DECAPx4_ASAP7_75t_R FILLER_217_824 ();
 FILLER_ASAP7_75t_R FILLER_217_837 ();
 DECAPx6_ASAP7_75t_R FILLER_217_842 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_856 ();
 DECAPx2_ASAP7_75t_R FILLER_217_873 ();
 DECAPx4_ASAP7_75t_R FILLER_217_882 ();
 FILLER_ASAP7_75t_R FILLER_217_892 ();
 DECAPx1_ASAP7_75t_R FILLER_217_897 ();
 FILLER_ASAP7_75t_R FILLER_217_905 ();
 DECAPx2_ASAP7_75t_R FILLER_217_916 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_922 ();
 DECAPx2_ASAP7_75t_R FILLER_217_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_933 ();
 FILLER_ASAP7_75t_R FILLER_217_940 ();
 DECAPx2_ASAP7_75t_R FILLER_217_949 ();
 FILLER_ASAP7_75t_R FILLER_217_955 ();
 DECAPx6_ASAP7_75t_R FILLER_217_965 ();
 FILLER_ASAP7_75t_R FILLER_217_985 ();
 DECAPx1_ASAP7_75t_R FILLER_217_993 ();
 FILLER_ASAP7_75t_R FILLER_217_1003 ();
 FILLER_ASAP7_75t_R FILLER_217_1008 ();
 DECAPx6_ASAP7_75t_R FILLER_217_1013 ();
 FILLER_ASAP7_75t_R FILLER_217_1030 ();
 FILLER_ASAP7_75t_R FILLER_217_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_217_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1061 ();
 FILLER_ASAP7_75t_R FILLER_217_1070 ();
 FILLER_ASAP7_75t_R FILLER_217_1086 ();
 FILLER_ASAP7_75t_R FILLER_217_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_217_1334 ();
 DECAPx6_ASAP7_75t_R FILLER_217_1356 ();
 DECAPx2_ASAP7_75t_R FILLER_217_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_1376 ();
 DECAPx4_ASAP7_75t_R FILLER_218_2 ();
 FILLER_ASAP7_75t_R FILLER_218_12 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_20 ();
 DECAPx2_ASAP7_75t_R FILLER_218_26 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_32 ();
 FILLER_ASAP7_75t_R FILLER_218_41 ();
 DECAPx1_ASAP7_75t_R FILLER_218_46 ();
 FILLER_ASAP7_75t_R FILLER_218_57 ();
 DECAPx1_ASAP7_75t_R FILLER_218_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_70 ();
 DECAPx6_ASAP7_75t_R FILLER_218_77 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_91 ();
 DECAPx6_ASAP7_75t_R FILLER_218_100 ();
 DECAPx2_ASAP7_75t_R FILLER_218_114 ();
 DECAPx2_ASAP7_75t_R FILLER_218_126 ();
 FILLER_ASAP7_75t_R FILLER_218_132 ();
 FILLER_ASAP7_75t_R FILLER_218_140 ();
 DECAPx2_ASAP7_75t_R FILLER_218_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_156 ();
 DECAPx6_ASAP7_75t_R FILLER_218_163 ();
 FILLER_ASAP7_75t_R FILLER_218_177 ();
 DECAPx4_ASAP7_75t_R FILLER_218_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_195 ();
 DECAPx4_ASAP7_75t_R FILLER_218_199 ();
 FILLER_ASAP7_75t_R FILLER_218_209 ();
 DECAPx4_ASAP7_75t_R FILLER_218_217 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_227 ();
 DECAPx10_ASAP7_75t_R FILLER_218_233 ();
 DECAPx6_ASAP7_75t_R FILLER_218_255 ();
 DECAPx2_ASAP7_75t_R FILLER_218_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_275 ();
 FILLER_ASAP7_75t_R FILLER_218_302 ();
 DECAPx4_ASAP7_75t_R FILLER_218_310 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_320 ();
 DECAPx6_ASAP7_75t_R FILLER_218_329 ();
 FILLER_ASAP7_75t_R FILLER_218_343 ();
 DECAPx1_ASAP7_75t_R FILLER_218_371 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_381 ();
 DECAPx4_ASAP7_75t_R FILLER_218_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_397 ();
 FILLER_ASAP7_75t_R FILLER_218_404 ();
 FILLER_ASAP7_75t_R FILLER_218_432 ();
 DECAPx4_ASAP7_75t_R FILLER_218_441 ();
 FILLER_ASAP7_75t_R FILLER_218_451 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_459 ();
 DECAPx4_ASAP7_75t_R FILLER_218_464 ();
 FILLER_ASAP7_75t_R FILLER_218_474 ();
 DECAPx6_ASAP7_75t_R FILLER_218_482 ();
 DECAPx1_ASAP7_75t_R FILLER_218_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_500 ();
 FILLER_ASAP7_75t_R FILLER_218_507 ();
 DECAPx2_ASAP7_75t_R FILLER_218_512 ();
 FILLER_ASAP7_75t_R FILLER_218_524 ();
 DECAPx1_ASAP7_75t_R FILLER_218_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_536 ();
 DECAPx6_ASAP7_75t_R FILLER_218_543 ();
 DECAPx1_ASAP7_75t_R FILLER_218_557 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_567 ();
 DECAPx4_ASAP7_75t_R FILLER_218_573 ();
 FILLER_ASAP7_75t_R FILLER_218_589 ();
 DECAPx6_ASAP7_75t_R FILLER_218_597 ();
 DECAPx2_ASAP7_75t_R FILLER_218_611 ();
 DECAPx1_ASAP7_75t_R FILLER_218_623 ();
 FILLER_ASAP7_75t_R FILLER_218_633 ();
 DECAPx6_ASAP7_75t_R FILLER_218_638 ();
 DECAPx1_ASAP7_75t_R FILLER_218_652 ();
 DECAPx1_ASAP7_75t_R FILLER_218_670 ();
 DECAPx2_ASAP7_75t_R FILLER_218_680 ();
 DECAPx1_ASAP7_75t_R FILLER_218_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_693 ();
 FILLER_ASAP7_75t_R FILLER_218_703 ();
 DECAPx10_ASAP7_75t_R FILLER_218_708 ();
 DECAPx2_ASAP7_75t_R FILLER_218_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_736 ();
 DECAPx1_ASAP7_75t_R FILLER_218_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_744 ();
 DECAPx1_ASAP7_75t_R FILLER_218_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_752 ();
 DECAPx4_ASAP7_75t_R FILLER_218_762 ();
 FILLER_ASAP7_75t_R FILLER_218_778 ();
 DECAPx4_ASAP7_75t_R FILLER_218_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_796 ();
 FILLER_ASAP7_75t_R FILLER_218_806 ();
 DECAPx10_ASAP7_75t_R FILLER_218_811 ();
 DECAPx6_ASAP7_75t_R FILLER_218_833 ();
 FILLER_ASAP7_75t_R FILLER_218_847 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_858 ();
 FILLER_ASAP7_75t_R FILLER_218_864 ();
 FILLER_ASAP7_75t_R FILLER_218_869 ();
 DECAPx1_ASAP7_75t_R FILLER_218_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_878 ();
 DECAPx4_ASAP7_75t_R FILLER_218_893 ();
 FILLER_ASAP7_75t_R FILLER_218_903 ();
 FILLER_ASAP7_75t_R FILLER_218_912 ();
 DECAPx2_ASAP7_75t_R FILLER_218_922 ();
 DECAPx4_ASAP7_75t_R FILLER_218_934 ();
 DECAPx1_ASAP7_75t_R FILLER_218_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_956 ();
 FILLER_ASAP7_75t_R FILLER_218_963 ();
 DECAPx2_ASAP7_75t_R FILLER_218_973 ();
 FILLER_ASAP7_75t_R FILLER_218_979 ();
 DECAPx6_ASAP7_75t_R FILLER_218_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1007 ();
 DECAPx6_ASAP7_75t_R FILLER_218_1014 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1037 ();
 DECAPx6_ASAP7_75t_R FILLER_218_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_218_1336 ();
 DECAPx6_ASAP7_75t_R FILLER_218_1358 ();
 DECAPx1_ASAP7_75t_R FILLER_218_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_219_2 ();
 DECAPx10_ASAP7_75t_R FILLER_219_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_56 ();
 FILLER_ASAP7_75t_R FILLER_219_83 ();
 FILLER_ASAP7_75t_R FILLER_219_111 ();
 FILLER_ASAP7_75t_R FILLER_219_139 ();
 DECAPx1_ASAP7_75t_R FILLER_219_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_151 ();
 FILLER_ASAP7_75t_R FILLER_219_158 ();
 DECAPx2_ASAP7_75t_R FILLER_219_166 ();
 DECAPx10_ASAP7_75t_R FILLER_219_198 ();
 DECAPx1_ASAP7_75t_R FILLER_219_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_224 ();
 FILLER_ASAP7_75t_R FILLER_219_231 ();
 DECAPx4_ASAP7_75t_R FILLER_219_236 ();
 FILLER_ASAP7_75t_R FILLER_219_246 ();
 FILLER_ASAP7_75t_R FILLER_219_254 ();
 DECAPx2_ASAP7_75t_R FILLER_219_262 ();
 DECAPx6_ASAP7_75t_R FILLER_219_274 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_219_288 ();
 DECAPx4_ASAP7_75t_R FILLER_219_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_304 ();
 DECAPx1_ASAP7_75t_R FILLER_219_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_317 ();
 DECAPx2_ASAP7_75t_R FILLER_219_326 ();
 FILLER_ASAP7_75t_R FILLER_219_332 ();
 DECAPx2_ASAP7_75t_R FILLER_219_340 ();
 FILLER_ASAP7_75t_R FILLER_219_346 ();
 DECAPx2_ASAP7_75t_R FILLER_219_354 ();
 DECAPx2_ASAP7_75t_R FILLER_219_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_369 ();
 DECAPx1_ASAP7_75t_R FILLER_219_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_400 ();
 DECAPx1_ASAP7_75t_R FILLER_219_404 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_219_414 ();
 FILLER_ASAP7_75t_R FILLER_219_420 ();
 DECAPx2_ASAP7_75t_R FILLER_219_429 ();
 FILLER_ASAP7_75t_R FILLER_219_435 ();
 FILLER_ASAP7_75t_R FILLER_219_463 ();
 FILLER_ASAP7_75t_R FILLER_219_491 ();
 DECAPx10_ASAP7_75t_R FILLER_219_499 ();
 DECAPx10_ASAP7_75t_R FILLER_219_521 ();
 DECAPx2_ASAP7_75t_R FILLER_219_543 ();
 FILLER_ASAP7_75t_R FILLER_219_549 ();
 FILLER_ASAP7_75t_R FILLER_219_577 ();
 DECAPx2_ASAP7_75t_R FILLER_219_605 ();
 DECAPx2_ASAP7_75t_R FILLER_219_637 ();
 FILLER_ASAP7_75t_R FILLER_219_643 ();
 FILLER_ASAP7_75t_R FILLER_219_651 ();
 DECAPx10_ASAP7_75t_R FILLER_219_656 ();
 DECAPx6_ASAP7_75t_R FILLER_219_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_692 ();
 FILLER_ASAP7_75t_R FILLER_219_702 ();
 FILLER_ASAP7_75t_R FILLER_219_707 ();
 FILLER_ASAP7_75t_R FILLER_219_723 ();
 DECAPx10_ASAP7_75t_R FILLER_219_728 ();
 FILLER_ASAP7_75t_R FILLER_219_750 ();
 FILLER_ASAP7_75t_R FILLER_219_761 ();
 DECAPx10_ASAP7_75t_R FILLER_219_766 ();
 FILLER_ASAP7_75t_R FILLER_219_797 ();
 FILLER_ASAP7_75t_R FILLER_219_802 ();
 DECAPx4_ASAP7_75t_R FILLER_219_807 ();
 FILLER_ASAP7_75t_R FILLER_219_817 ();
 DECAPx6_ASAP7_75t_R FILLER_219_825 ();
 FILLER_ASAP7_75t_R FILLER_219_839 ();
 DECAPx6_ASAP7_75t_R FILLER_219_844 ();
 DECAPx1_ASAP7_75t_R FILLER_219_858 ();
 DECAPx2_ASAP7_75t_R FILLER_219_871 ();
 FILLER_ASAP7_75t_R FILLER_219_877 ();
 FILLER_ASAP7_75t_R FILLER_219_882 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_219_887 ();
 FILLER_ASAP7_75t_R FILLER_219_893 ();
 DECAPx1_ASAP7_75t_R FILLER_219_904 ();
 DECAPx2_ASAP7_75t_R FILLER_219_916 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_219_922 ();
 DECAPx1_ASAP7_75t_R FILLER_219_927 ();
 DECAPx6_ASAP7_75t_R FILLER_219_937 ();
 FILLER_ASAP7_75t_R FILLER_219_951 ();
 DECAPx4_ASAP7_75t_R FILLER_219_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_969 ();
 DECAPx1_ASAP7_75t_R FILLER_219_976 ();
 DECAPx4_ASAP7_75t_R FILLER_219_994 ();
 FILLER_ASAP7_75t_R FILLER_219_1004 ();
 FILLER_ASAP7_75t_R FILLER_219_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_219_1025 ();
 FILLER_ASAP7_75t_R FILLER_219_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_219_1047 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_219_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1070 ();
 DECAPx4_ASAP7_75t_R FILLER_219_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_219_1335 ();
 DECAPx6_ASAP7_75t_R FILLER_219_1357 ();
 DECAPx2_ASAP7_75t_R FILLER_219_1371 ();
 DECAPx2_ASAP7_75t_R FILLER_220_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_220_8 ();
 DECAPx6_ASAP7_75t_R FILLER_220_17 ();
 DECAPx1_ASAP7_75t_R FILLER_220_31 ();
 DECAPx6_ASAP7_75t_R FILLER_220_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_52 ();
 DECAPx2_ASAP7_75t_R FILLER_220_59 ();
 DECAPx1_ASAP7_75t_R FILLER_220_71 ();
 DECAPx2_ASAP7_75t_R FILLER_220_78 ();
 FILLER_ASAP7_75t_R FILLER_220_87 ();
 DECAPx2_ASAP7_75t_R FILLER_220_95 ();
 DECAPx4_ASAP7_75t_R FILLER_220_104 ();
 FILLER_ASAP7_75t_R FILLER_220_114 ();
 DECAPx2_ASAP7_75t_R FILLER_220_122 ();
 DECAPx6_ASAP7_75t_R FILLER_220_131 ();
 DECAPx1_ASAP7_75t_R FILLER_220_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_149 ();
 DECAPx6_ASAP7_75t_R FILLER_220_158 ();
 FILLER_ASAP7_75t_R FILLER_220_172 ();
 DECAPx2_ASAP7_75t_R FILLER_220_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_186 ();
 DECAPx10_ASAP7_75t_R FILLER_220_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_212 ();
 FILLER_ASAP7_75t_R FILLER_220_239 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_220_244 ();
 FILLER_ASAP7_75t_R FILLER_220_255 ();
 FILLER_ASAP7_75t_R FILLER_220_263 ();
 DECAPx4_ASAP7_75t_R FILLER_220_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_301 ();
 FILLER_ASAP7_75t_R FILLER_220_308 ();
 DECAPx2_ASAP7_75t_R FILLER_220_316 ();
 FILLER_ASAP7_75t_R FILLER_220_322 ();
 FILLER_ASAP7_75t_R FILLER_220_330 ();
 DECAPx6_ASAP7_75t_R FILLER_220_358 ();
 DECAPx4_ASAP7_75t_R FILLER_220_378 ();
 FILLER_ASAP7_75t_R FILLER_220_388 ();
 DECAPx10_ASAP7_75t_R FILLER_220_396 ();
 DECAPx2_ASAP7_75t_R FILLER_220_418 ();
 FILLER_ASAP7_75t_R FILLER_220_424 ();
 FILLER_ASAP7_75t_R FILLER_220_452 ();
 FILLER_ASAP7_75t_R FILLER_220_460 ();
 DECAPx2_ASAP7_75t_R FILLER_220_464 ();
 FILLER_ASAP7_75t_R FILLER_220_476 ();
 FILLER_ASAP7_75t_R FILLER_220_481 ();
 FILLER_ASAP7_75t_R FILLER_220_489 ();
 FILLER_ASAP7_75t_R FILLER_220_499 ();
 DECAPx4_ASAP7_75t_R FILLER_220_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_517 ();
 DECAPx6_ASAP7_75t_R FILLER_220_524 ();
 DECAPx1_ASAP7_75t_R FILLER_220_538 ();
 DECAPx4_ASAP7_75t_R FILLER_220_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_558 ();
 FILLER_ASAP7_75t_R FILLER_220_565 ();
 DECAPx10_ASAP7_75t_R FILLER_220_570 ();
 FILLER_ASAP7_75t_R FILLER_220_592 ();
 DECAPx1_ASAP7_75t_R FILLER_220_597 ();
 DECAPx6_ASAP7_75t_R FILLER_220_607 ();
 DECAPx1_ASAP7_75t_R FILLER_220_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_625 ();
 DECAPx1_ASAP7_75t_R FILLER_220_629 ();
 FILLER_ASAP7_75t_R FILLER_220_639 ();
 DECAPx4_ASAP7_75t_R FILLER_220_655 ();
 FILLER_ASAP7_75t_R FILLER_220_665 ();
 DECAPx4_ASAP7_75t_R FILLER_220_676 ();
 DECAPx2_ASAP7_75t_R FILLER_220_689 ();
 FILLER_ASAP7_75t_R FILLER_220_695 ();
 DECAPx4_ASAP7_75t_R FILLER_220_711 ();
 DECAPx2_ASAP7_75t_R FILLER_220_724 ();
 DECAPx2_ASAP7_75t_R FILLER_220_744 ();
 DECAPx10_ASAP7_75t_R FILLER_220_753 ();
 FILLER_ASAP7_75t_R FILLER_220_775 ();
 DECAPx10_ASAP7_75t_R FILLER_220_783 ();
 DECAPx2_ASAP7_75t_R FILLER_220_805 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_220_811 ();
 FILLER_ASAP7_75t_R FILLER_220_820 ();
 DECAPx2_ASAP7_75t_R FILLER_220_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_837 ();
 FILLER_ASAP7_75t_R FILLER_220_847 ();
 DECAPx6_ASAP7_75t_R FILLER_220_852 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_220_866 ();
 DECAPx6_ASAP7_75t_R FILLER_220_872 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_220_886 ();
 DECAPx10_ASAP7_75t_R FILLER_220_892 ();
 DECAPx4_ASAP7_75t_R FILLER_220_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_924 ();
 DECAPx10_ASAP7_75t_R FILLER_220_932 ();
 DECAPx10_ASAP7_75t_R FILLER_220_954 ();
 DECAPx6_ASAP7_75t_R FILLER_220_976 ();
 DECAPx1_ASAP7_75t_R FILLER_220_990 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1001 ();
 FILLER_ASAP7_75t_R FILLER_220_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1015 ();
 FILLER_ASAP7_75t_R FILLER_220_1022 ();
 FILLER_ASAP7_75t_R FILLER_220_1030 ();
 FILLER_ASAP7_75t_R FILLER_220_1046 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1055 ();
 DECAPx1_ASAP7_75t_R FILLER_220_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_1074 ();
 DECAPx4_ASAP7_75t_R FILLER_220_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_220_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_220_1353 ();
 FILLER_ASAP7_75t_R FILLER_220_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_221_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_16 ();
 FILLER_ASAP7_75t_R FILLER_221_23 ();
 DECAPx2_ASAP7_75t_R FILLER_221_31 ();
 FILLER_ASAP7_75t_R FILLER_221_37 ();
 DECAPx1_ASAP7_75t_R FILLER_221_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_49 ();
 DECAPx6_ASAP7_75t_R FILLER_221_76 ();
 DECAPx1_ASAP7_75t_R FILLER_221_90 ();
 FILLER_ASAP7_75t_R FILLER_221_102 ();
 DECAPx10_ASAP7_75t_R FILLER_221_110 ();
 DECAPx6_ASAP7_75t_R FILLER_221_132 ();
 DECAPx1_ASAP7_75t_R FILLER_221_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_150 ();
 DECAPx6_ASAP7_75t_R FILLER_221_159 ();
 FILLER_ASAP7_75t_R FILLER_221_173 ();
 DECAPx4_ASAP7_75t_R FILLER_221_181 ();
 FILLER_ASAP7_75t_R FILLER_221_197 ();
 FILLER_ASAP7_75t_R FILLER_221_207 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_215 ();
 FILLER_ASAP7_75t_R FILLER_221_224 ();
 DECAPx6_ASAP7_75t_R FILLER_221_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_246 ();
 DECAPx4_ASAP7_75t_R FILLER_221_255 ();
 FILLER_ASAP7_75t_R FILLER_221_265 ();
 DECAPx2_ASAP7_75t_R FILLER_221_273 ();
 DECAPx2_ASAP7_75t_R FILLER_221_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_288 ();
 DECAPx2_ASAP7_75t_R FILLER_221_295 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_301 ();
 DECAPx2_ASAP7_75t_R FILLER_221_307 ();
 FILLER_ASAP7_75t_R FILLER_221_313 ();
 DECAPx4_ASAP7_75t_R FILLER_221_323 ();
 DECAPx2_ASAP7_75t_R FILLER_221_339 ();
 FILLER_ASAP7_75t_R FILLER_221_345 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_350 ();
 DECAPx4_ASAP7_75t_R FILLER_221_359 ();
 FILLER_ASAP7_75t_R FILLER_221_369 ();
 DECAPx1_ASAP7_75t_R FILLER_221_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_381 ();
 FILLER_ASAP7_75t_R FILLER_221_408 ();
 DECAPx4_ASAP7_75t_R FILLER_221_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_428 ();
 FILLER_ASAP7_75t_R FILLER_221_435 ();
 FILLER_ASAP7_75t_R FILLER_221_443 ();
 DECAPx4_ASAP7_75t_R FILLER_221_448 ();
 DECAPx4_ASAP7_75t_R FILLER_221_461 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_471 ();
 DECAPx6_ASAP7_75t_R FILLER_221_477 ();
 DECAPx1_ASAP7_75t_R FILLER_221_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_495 ();
 DECAPx1_ASAP7_75t_R FILLER_221_504 ();
 FILLER_ASAP7_75t_R FILLER_221_534 ();
 FILLER_ASAP7_75t_R FILLER_221_539 ();
 DECAPx2_ASAP7_75t_R FILLER_221_547 ();
 FILLER_ASAP7_75t_R FILLER_221_553 ();
 DECAPx6_ASAP7_75t_R FILLER_221_563 ();
 DECAPx1_ASAP7_75t_R FILLER_221_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_581 ();
 DECAPx2_ASAP7_75t_R FILLER_221_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_594 ();
 FILLER_ASAP7_75t_R FILLER_221_601 ();
 DECAPx10_ASAP7_75t_R FILLER_221_611 ();
 DECAPx4_ASAP7_75t_R FILLER_221_633 ();
 FILLER_ASAP7_75t_R FILLER_221_643 ();
 FILLER_ASAP7_75t_R FILLER_221_651 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_667 ();
 FILLER_ASAP7_75t_R FILLER_221_676 ();
 DECAPx6_ASAP7_75t_R FILLER_221_687 ();
 DECAPx2_ASAP7_75t_R FILLER_221_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_707 ();
 DECAPx6_ASAP7_75t_R FILLER_221_711 ();
 DECAPx1_ASAP7_75t_R FILLER_221_725 ();
 FILLER_ASAP7_75t_R FILLER_221_732 ();
 DECAPx2_ASAP7_75t_R FILLER_221_748 ();
 FILLER_ASAP7_75t_R FILLER_221_754 ();
 FILLER_ASAP7_75t_R FILLER_221_762 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_767 ();
 FILLER_ASAP7_75t_R FILLER_221_776 ();
 DECAPx2_ASAP7_75t_R FILLER_221_792 ();
 FILLER_ASAP7_75t_R FILLER_221_798 ();
 FILLER_ASAP7_75t_R FILLER_221_809 ();
 DECAPx2_ASAP7_75t_R FILLER_221_814 ();
 FILLER_ASAP7_75t_R FILLER_221_834 ();
 DECAPx10_ASAP7_75t_R FILLER_221_839 ();
 DECAPx2_ASAP7_75t_R FILLER_221_861 ();
 FILLER_ASAP7_75t_R FILLER_221_867 ();
 DECAPx2_ASAP7_75t_R FILLER_221_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_889 ();
 FILLER_ASAP7_75t_R FILLER_221_894 ();
 FILLER_ASAP7_75t_R FILLER_221_910 ();
 DECAPx2_ASAP7_75t_R FILLER_221_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_924 ();
 DECAPx4_ASAP7_75t_R FILLER_221_927 ();
 DECAPx4_ASAP7_75t_R FILLER_221_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_959 ();
 DECAPx10_ASAP7_75t_R FILLER_221_972 ();
 FILLER_ASAP7_75t_R FILLER_221_994 ();
 DECAPx10_ASAP7_75t_R FILLER_221_999 ();
 DECAPx4_ASAP7_75t_R FILLER_221_1021 ();
 DECAPx6_ASAP7_75t_R FILLER_221_1041 ();
 DECAPx4_ASAP7_75t_R FILLER_221_1058 ();
 FILLER_ASAP7_75t_R FILLER_221_1068 ();
 FILLER_ASAP7_75t_R FILLER_221_1073 ();
 DECAPx1_ASAP7_75t_R FILLER_221_1089 ();
 FILLER_ASAP7_75t_R FILLER_221_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_221_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_1376 ();
 DECAPx4_ASAP7_75t_R FILLER_222_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_12 ();
 DECAPx1_ASAP7_75t_R FILLER_222_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_43 ();
 DECAPx2_ASAP7_75t_R FILLER_222_52 ();
 FILLER_ASAP7_75t_R FILLER_222_64 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_69 ();
 DECAPx6_ASAP7_75t_R FILLER_222_75 ();
 FILLER_ASAP7_75t_R FILLER_222_89 ();
 FILLER_ASAP7_75t_R FILLER_222_99 ();
 DECAPx4_ASAP7_75t_R FILLER_222_107 ();
 FILLER_ASAP7_75t_R FILLER_222_117 ();
 DECAPx4_ASAP7_75t_R FILLER_222_125 ();
 FILLER_ASAP7_75t_R FILLER_222_135 ();
 DECAPx4_ASAP7_75t_R FILLER_222_140 ();
 FILLER_ASAP7_75t_R FILLER_222_150 ();
 FILLER_ASAP7_75t_R FILLER_222_158 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_166 ();
 FILLER_ASAP7_75t_R FILLER_222_195 ();
 DECAPx2_ASAP7_75t_R FILLER_222_219 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_225 ();
 DECAPx2_ASAP7_75t_R FILLER_222_234 ();
 DECAPx6_ASAP7_75t_R FILLER_222_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_257 ();
 DECAPx6_ASAP7_75t_R FILLER_222_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_278 ();
 DECAPx10_ASAP7_75t_R FILLER_222_305 ();
 DECAPx10_ASAP7_75t_R FILLER_222_327 ();
 FILLER_ASAP7_75t_R FILLER_222_349 ();
 DECAPx2_ASAP7_75t_R FILLER_222_377 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_383 ();
 DECAPx1_ASAP7_75t_R FILLER_222_392 ();
 DECAPx2_ASAP7_75t_R FILLER_222_399 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_408 ();
 FILLER_ASAP7_75t_R FILLER_222_419 ();
 DECAPx6_ASAP7_75t_R FILLER_222_427 ();
 DECAPx1_ASAP7_75t_R FILLER_222_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_445 ();
 FILLER_ASAP7_75t_R FILLER_222_452 ();
 FILLER_ASAP7_75t_R FILLER_222_460 ();
 DECAPx2_ASAP7_75t_R FILLER_222_464 ();
 FILLER_ASAP7_75t_R FILLER_222_470 ();
 DECAPx2_ASAP7_75t_R FILLER_222_478 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_484 ();
 DECAPx10_ASAP7_75t_R FILLER_222_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_512 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_519 ();
 DECAPx2_ASAP7_75t_R FILLER_222_525 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_531 ();
 DECAPx4_ASAP7_75t_R FILLER_222_542 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_552 ();
 DECAPx2_ASAP7_75t_R FILLER_222_563 ();
 FILLER_ASAP7_75t_R FILLER_222_595 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_600 ();
 DECAPx2_ASAP7_75t_R FILLER_222_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_617 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_626 ();
 DECAPx2_ASAP7_75t_R FILLER_222_638 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_644 ();
 DECAPx1_ASAP7_75t_R FILLER_222_650 ();
 DECAPx6_ASAP7_75t_R FILLER_222_657 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_671 ();
 FILLER_ASAP7_75t_R FILLER_222_680 ();
 DECAPx2_ASAP7_75t_R FILLER_222_685 ();
 FILLER_ASAP7_75t_R FILLER_222_691 ();
 DECAPx4_ASAP7_75t_R FILLER_222_696 ();
 FILLER_ASAP7_75t_R FILLER_222_706 ();
 FILLER_ASAP7_75t_R FILLER_222_722 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_727 ();
 DECAPx6_ASAP7_75t_R FILLER_222_744 ();
 DECAPx4_ASAP7_75t_R FILLER_222_767 ();
 DECAPx4_ASAP7_75t_R FILLER_222_783 ();
 FILLER_ASAP7_75t_R FILLER_222_793 ();
 FILLER_ASAP7_75t_R FILLER_222_809 ();
 DECAPx2_ASAP7_75t_R FILLER_222_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_824 ();
 DECAPx2_ASAP7_75t_R FILLER_222_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_834 ();
 DECAPx2_ASAP7_75t_R FILLER_222_838 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_844 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_850 ();
 FILLER_ASAP7_75t_R FILLER_222_862 ();
 DECAPx4_ASAP7_75t_R FILLER_222_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_877 ();
 DECAPx2_ASAP7_75t_R FILLER_222_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_898 ();
 FILLER_ASAP7_75t_R FILLER_222_910 ();
 DECAPx1_ASAP7_75t_R FILLER_222_918 ();
 FILLER_ASAP7_75t_R FILLER_222_931 ();
 FILLER_ASAP7_75t_R FILLER_222_947 ();
 DECAPx2_ASAP7_75t_R FILLER_222_952 ();
 FILLER_ASAP7_75t_R FILLER_222_961 ();
 FILLER_ASAP7_75t_R FILLER_222_977 ();
 DECAPx2_ASAP7_75t_R FILLER_222_986 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_992 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1010 ();
 FILLER_ASAP7_75t_R FILLER_222_1017 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_222_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_1091 ();
 FILLER_ASAP7_75t_R FILLER_222_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_222_1335 ();
 DECAPx6_ASAP7_75t_R FILLER_222_1357 ();
 DECAPx2_ASAP7_75t_R FILLER_222_1371 ();
 DECAPx2_ASAP7_75t_R FILLER_223_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_8 ();
 DECAPx4_ASAP7_75t_R FILLER_223_15 ();
 FILLER_ASAP7_75t_R FILLER_223_25 ();
 DECAPx1_ASAP7_75t_R FILLER_223_30 ();
 FILLER_ASAP7_75t_R FILLER_223_40 ();
 DECAPx10_ASAP7_75t_R FILLER_223_50 ();
 DECAPx1_ASAP7_75t_R FILLER_223_72 ();
 DECAPx2_ASAP7_75t_R FILLER_223_84 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_90 ();
 DECAPx4_ASAP7_75t_R FILLER_223_99 ();
 FILLER_ASAP7_75t_R FILLER_223_109 ();
 DECAPx2_ASAP7_75t_R FILLER_223_137 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_143 ();
 DECAPx10_ASAP7_75t_R FILLER_223_149 ();
 DECAPx1_ASAP7_75t_R FILLER_223_177 ();
 FILLER_ASAP7_75t_R FILLER_223_184 ();
 FILLER_ASAP7_75t_R FILLER_223_189 ();
 FILLER_ASAP7_75t_R FILLER_223_197 ();
 DECAPx2_ASAP7_75t_R FILLER_223_207 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_213 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_242 ();
 FILLER_ASAP7_75t_R FILLER_223_253 ();
 DECAPx2_ASAP7_75t_R FILLER_223_262 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_268 ();
 DECAPx1_ASAP7_75t_R FILLER_223_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_281 ();
 DECAPx2_ASAP7_75t_R FILLER_223_288 ();
 DECAPx1_ASAP7_75t_R FILLER_223_297 ();
 DECAPx1_ASAP7_75t_R FILLER_223_307 ();
 FILLER_ASAP7_75t_R FILLER_223_317 ();
 DECAPx4_ASAP7_75t_R FILLER_223_322 ();
 FILLER_ASAP7_75t_R FILLER_223_332 ();
 FILLER_ASAP7_75t_R FILLER_223_340 ();
 DECAPx6_ASAP7_75t_R FILLER_223_345 ();
 DECAPx2_ASAP7_75t_R FILLER_223_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_365 ();
 FILLER_ASAP7_75t_R FILLER_223_372 ();
 DECAPx10_ASAP7_75t_R FILLER_223_377 ();
 DECAPx2_ASAP7_75t_R FILLER_223_399 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_405 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_414 ();
 DECAPx2_ASAP7_75t_R FILLER_223_423 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_429 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_438 ();
 FILLER_ASAP7_75t_R FILLER_223_447 ();
 DECAPx1_ASAP7_75t_R FILLER_223_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_461 ();
 DECAPx1_ASAP7_75t_R FILLER_223_488 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_500 ();
 DECAPx6_ASAP7_75t_R FILLER_223_509 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_523 ();
 FILLER_ASAP7_75t_R FILLER_223_532 ();
 FILLER_ASAP7_75t_R FILLER_223_542 ();
 DECAPx2_ASAP7_75t_R FILLER_223_550 ();
 FILLER_ASAP7_75t_R FILLER_223_562 ();
 DECAPx1_ASAP7_75t_R FILLER_223_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_574 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_581 ();
 DECAPx4_ASAP7_75t_R FILLER_223_587 ();
 DECAPx2_ASAP7_75t_R FILLER_223_604 ();
 FILLER_ASAP7_75t_R FILLER_223_616 ();
 FILLER_ASAP7_75t_R FILLER_223_626 ();
 DECAPx10_ASAP7_75t_R FILLER_223_637 ();
 DECAPx10_ASAP7_75t_R FILLER_223_659 ();
 DECAPx2_ASAP7_75t_R FILLER_223_681 ();
 FILLER_ASAP7_75t_R FILLER_223_687 ();
 DECAPx1_ASAP7_75t_R FILLER_223_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_707 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_711 ();
 DECAPx6_ASAP7_75t_R FILLER_223_717 ();
 DECAPx1_ASAP7_75t_R FILLER_223_731 ();
 DECAPx4_ASAP7_75t_R FILLER_223_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_756 ();
 DECAPx4_ASAP7_75t_R FILLER_223_763 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_773 ();
 DECAPx6_ASAP7_75t_R FILLER_223_782 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_796 ();
 DECAPx10_ASAP7_75t_R FILLER_223_802 ();
 DECAPx10_ASAP7_75t_R FILLER_223_824 ();
 DECAPx1_ASAP7_75t_R FILLER_223_846 ();
 DECAPx2_ASAP7_75t_R FILLER_223_853 ();
 FILLER_ASAP7_75t_R FILLER_223_859 ();
 DECAPx4_ASAP7_75t_R FILLER_223_864 ();
 FILLER_ASAP7_75t_R FILLER_223_877 ();
 DECAPx6_ASAP7_75t_R FILLER_223_882 ();
 DECAPx2_ASAP7_75t_R FILLER_223_896 ();
 FILLER_ASAP7_75t_R FILLER_223_911 ();
 DECAPx2_ASAP7_75t_R FILLER_223_919 ();
 FILLER_ASAP7_75t_R FILLER_223_927 ();
 DECAPx10_ASAP7_75t_R FILLER_223_937 ();
 DECAPx2_ASAP7_75t_R FILLER_223_959 ();
 DECAPx2_ASAP7_75t_R FILLER_223_974 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_980 ();
 DECAPx6_ASAP7_75t_R FILLER_223_992 ();
 DECAPx1_ASAP7_75t_R FILLER_223_1006 ();
 FILLER_ASAP7_75t_R FILLER_223_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_223_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1057 ();
 FILLER_ASAP7_75t_R FILLER_223_1062 ();
 FILLER_ASAP7_75t_R FILLER_223_1068 ();
 DECAPx4_ASAP7_75t_R FILLER_223_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1083 ();
 DECAPx6_ASAP7_75t_R FILLER_223_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_223_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_223_1350 ();
 DECAPx1_ASAP7_75t_R FILLER_223_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_1376 ();
 FILLER_ASAP7_75t_R FILLER_224_2 ();
 DECAPx6_ASAP7_75t_R FILLER_224_30 ();
 DECAPx2_ASAP7_75t_R FILLER_224_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_50 ();
 DECAPx4_ASAP7_75t_R FILLER_224_57 ();
 FILLER_ASAP7_75t_R FILLER_224_67 ();
 FILLER_ASAP7_75t_R FILLER_224_75 ();
 DECAPx2_ASAP7_75t_R FILLER_224_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_91 ();
 DECAPx2_ASAP7_75t_R FILLER_224_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_104 ();
 DECAPx1_ASAP7_75t_R FILLER_224_111 ();
 DECAPx1_ASAP7_75t_R FILLER_224_121 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_224_128 ();
 FILLER_ASAP7_75t_R FILLER_224_157 ();
 DECAPx4_ASAP7_75t_R FILLER_224_165 ();
 FILLER_ASAP7_75t_R FILLER_224_175 ();
 DECAPx1_ASAP7_75t_R FILLER_224_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_187 ();
 FILLER_ASAP7_75t_R FILLER_224_195 ();
 FILLER_ASAP7_75t_R FILLER_224_204 ();
 DECAPx2_ASAP7_75t_R FILLER_224_214 ();
 FILLER_ASAP7_75t_R FILLER_224_220 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_224_228 ();
 DECAPx4_ASAP7_75t_R FILLER_224_234 ();
 FILLER_ASAP7_75t_R FILLER_224_244 ();
 DECAPx4_ASAP7_75t_R FILLER_224_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_264 ();
 DECAPx2_ASAP7_75t_R FILLER_224_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_297 ();
 DECAPx1_ASAP7_75t_R FILLER_224_324 ();
 DECAPx2_ASAP7_75t_R FILLER_224_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_360 ();
 DECAPx1_ASAP7_75t_R FILLER_224_367 ();
 DECAPx6_ASAP7_75t_R FILLER_224_377 ();
 FILLER_ASAP7_75t_R FILLER_224_391 ();
 FILLER_ASAP7_75t_R FILLER_224_399 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_224_404 ();
 DECAPx2_ASAP7_75t_R FILLER_224_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_419 ();
 DECAPx1_ASAP7_75t_R FILLER_224_446 ();
 DECAPx1_ASAP7_75t_R FILLER_224_458 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_224_464 ();
 DECAPx1_ASAP7_75t_R FILLER_224_473 ();
 DECAPx2_ASAP7_75t_R FILLER_224_480 ();
 FILLER_ASAP7_75t_R FILLER_224_486 ();
 FILLER_ASAP7_75t_R FILLER_224_494 ();
 DECAPx6_ASAP7_75t_R FILLER_224_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_518 ();
 DECAPx2_ASAP7_75t_R FILLER_224_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_531 ();
 DECAPx2_ASAP7_75t_R FILLER_224_538 ();
 DECAPx10_ASAP7_75t_R FILLER_224_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_572 ();
 DECAPx2_ASAP7_75t_R FILLER_224_579 ();
 FILLER_ASAP7_75t_R FILLER_224_585 ();
 FILLER_ASAP7_75t_R FILLER_224_590 ();
 FILLER_ASAP7_75t_R FILLER_224_599 ();
 FILLER_ASAP7_75t_R FILLER_224_609 ();
 DECAPx2_ASAP7_75t_R FILLER_224_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_623 ();
 DECAPx6_ASAP7_75t_R FILLER_224_630 ();
 DECAPx1_ASAP7_75t_R FILLER_224_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_648 ();
 DECAPx2_ASAP7_75t_R FILLER_224_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_661 ();
 FILLER_ASAP7_75t_R FILLER_224_671 ();
 DECAPx4_ASAP7_75t_R FILLER_224_676 ();
 FILLER_ASAP7_75t_R FILLER_224_686 ();
 FILLER_ASAP7_75t_R FILLER_224_697 ();
 DECAPx2_ASAP7_75t_R FILLER_224_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_708 ();
 DECAPx4_ASAP7_75t_R FILLER_224_723 ();
 DECAPx1_ASAP7_75t_R FILLER_224_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_751 ();
 DECAPx1_ASAP7_75t_R FILLER_224_761 ();
 FILLER_ASAP7_75t_R FILLER_224_771 ();
 DECAPx4_ASAP7_75t_R FILLER_224_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_797 ();
 DECAPx1_ASAP7_75t_R FILLER_224_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_816 ();
 DECAPx1_ASAP7_75t_R FILLER_224_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_824 ();
 FILLER_ASAP7_75t_R FILLER_224_839 ();
 DECAPx2_ASAP7_75t_R FILLER_224_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_856 ();
 DECAPx4_ASAP7_75t_R FILLER_224_860 ();
 DECAPx10_ASAP7_75t_R FILLER_224_879 ();
 DECAPx10_ASAP7_75t_R FILLER_224_901 ();
 FILLER_ASAP7_75t_R FILLER_224_923 ();
 DECAPx6_ASAP7_75t_R FILLER_224_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_945 ();
 DECAPx6_ASAP7_75t_R FILLER_224_958 ();
 FILLER_ASAP7_75t_R FILLER_224_972 ();
 DECAPx4_ASAP7_75t_R FILLER_224_981 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_224_991 ();
 DECAPx4_ASAP7_75t_R FILLER_224_1008 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_224_1018 ();
 FILLER_ASAP7_75t_R FILLER_224_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_224_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1053 ();
 FILLER_ASAP7_75t_R FILLER_224_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_224_1344 ();
 DECAPx4_ASAP7_75t_R FILLER_224_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_1376 ();
 DECAPx1_ASAP7_75t_R FILLER_225_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_6 ();
 DECAPx1_ASAP7_75t_R FILLER_225_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_17 ();
 DECAPx4_ASAP7_75t_R FILLER_225_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_31 ();
 DECAPx2_ASAP7_75t_R FILLER_225_35 ();
 FILLER_ASAP7_75t_R FILLER_225_49 ();
 DECAPx1_ASAP7_75t_R FILLER_225_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_61 ();
 DECAPx2_ASAP7_75t_R FILLER_225_68 ();
 DECAPx6_ASAP7_75t_R FILLER_225_80 ();
 DECAPx6_ASAP7_75t_R FILLER_225_101 ();
 DECAPx1_ASAP7_75t_R FILLER_225_115 ();
 DECAPx2_ASAP7_75t_R FILLER_225_125 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_225_131 ();
 DECAPx10_ASAP7_75t_R FILLER_225_140 ();
 DECAPx2_ASAP7_75t_R FILLER_225_162 ();
 FILLER_ASAP7_75t_R FILLER_225_168 ();
 FILLER_ASAP7_75t_R FILLER_225_196 ();
 FILLER_ASAP7_75t_R FILLER_225_205 ();
 DECAPx10_ASAP7_75t_R FILLER_225_215 ();
 DECAPx2_ASAP7_75t_R FILLER_225_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_243 ();
 FILLER_ASAP7_75t_R FILLER_225_250 ();
 DECAPx2_ASAP7_75t_R FILLER_225_258 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_225_264 ();
 DECAPx2_ASAP7_75t_R FILLER_225_273 ();
 DECAPx1_ASAP7_75t_R FILLER_225_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_286 ();
 DECAPx6_ASAP7_75t_R FILLER_225_290 ();
 FILLER_ASAP7_75t_R FILLER_225_304 ();
 FILLER_ASAP7_75t_R FILLER_225_309 ();
 FILLER_ASAP7_75t_R FILLER_225_317 ();
 FILLER_ASAP7_75t_R FILLER_225_326 ();
 FILLER_ASAP7_75t_R FILLER_225_335 ();
 DECAPx2_ASAP7_75t_R FILLER_225_344 ();
 DECAPx2_ASAP7_75t_R FILLER_225_356 ();
 FILLER_ASAP7_75t_R FILLER_225_368 ();
 DECAPx2_ASAP7_75t_R FILLER_225_378 ();
 FILLER_ASAP7_75t_R FILLER_225_384 ();
 DECAPx6_ASAP7_75t_R FILLER_225_412 ();
 FILLER_ASAP7_75t_R FILLER_225_426 ();
 FILLER_ASAP7_75t_R FILLER_225_434 ();
 DECAPx1_ASAP7_75t_R FILLER_225_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_443 ();
 DECAPx10_ASAP7_75t_R FILLER_225_447 ();
 DECAPx2_ASAP7_75t_R FILLER_225_469 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_225_475 ();
 DECAPx4_ASAP7_75t_R FILLER_225_484 ();
 DECAPx4_ASAP7_75t_R FILLER_225_500 ();
 FILLER_ASAP7_75t_R FILLER_225_510 ();
 DECAPx6_ASAP7_75t_R FILLER_225_538 ();
 DECAPx1_ASAP7_75t_R FILLER_225_552 ();
 DECAPx2_ASAP7_75t_R FILLER_225_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_568 ();
 DECAPx2_ASAP7_75t_R FILLER_225_595 ();
 FILLER_ASAP7_75t_R FILLER_225_609 ();
 DECAPx10_ASAP7_75t_R FILLER_225_618 ();
 FILLER_ASAP7_75t_R FILLER_225_640 ();
 DECAPx2_ASAP7_75t_R FILLER_225_656 ();
 FILLER_ASAP7_75t_R FILLER_225_662 ();
 FILLER_ASAP7_75t_R FILLER_225_678 ();
 DECAPx2_ASAP7_75t_R FILLER_225_683 ();
 FILLER_ASAP7_75t_R FILLER_225_703 ();
 DECAPx10_ASAP7_75t_R FILLER_225_708 ();
 DECAPx4_ASAP7_75t_R FILLER_225_730 ();
 DECAPx10_ASAP7_75t_R FILLER_225_743 ();
 DECAPx1_ASAP7_75t_R FILLER_225_765 ();
 FILLER_ASAP7_75t_R FILLER_225_772 ();
 DECAPx4_ASAP7_75t_R FILLER_225_780 ();
 FILLER_ASAP7_75t_R FILLER_225_790 ();
 DECAPx2_ASAP7_75t_R FILLER_225_806 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_225_812 ();
 FILLER_ASAP7_75t_R FILLER_225_821 ();
 DECAPx2_ASAP7_75t_R FILLER_225_837 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_225_843 ();
 FILLER_ASAP7_75t_R FILLER_225_849 ();
 DECAPx4_ASAP7_75t_R FILLER_225_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_875 ();
 FILLER_ASAP7_75t_R FILLER_225_879 ();
 DECAPx4_ASAP7_75t_R FILLER_225_884 ();
 FILLER_ASAP7_75t_R FILLER_225_894 ();
 FILLER_ASAP7_75t_R FILLER_225_899 ();
 DECAPx6_ASAP7_75t_R FILLER_225_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_924 ();
 DECAPx10_ASAP7_75t_R FILLER_225_927 ();
 DECAPx6_ASAP7_75t_R FILLER_225_949 ();
 DECAPx2_ASAP7_75t_R FILLER_225_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_976 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_225_991 ();
 FILLER_ASAP7_75t_R FILLER_225_997 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1013 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_225_1019 ();
 FILLER_ASAP7_75t_R FILLER_225_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_225_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1048 ();
 FILLER_ASAP7_75t_R FILLER_225_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_225_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_225_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1083 ();
 DECAPx1_ASAP7_75t_R FILLER_225_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_1102 ();
 DECAPx1_ASAP7_75t_R FILLER_225_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_225_1355 ();
 DECAPx2_ASAP7_75t_R FILLER_226_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_8 ();
 FILLER_ASAP7_75t_R FILLER_226_17 ();
 DECAPx2_ASAP7_75t_R FILLER_226_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_31 ();
 FILLER_ASAP7_75t_R FILLER_226_38 ();
 DECAPx2_ASAP7_75t_R FILLER_226_48 ();
 FILLER_ASAP7_75t_R FILLER_226_54 ();
 DECAPx6_ASAP7_75t_R FILLER_226_82 ();
 DECAPx1_ASAP7_75t_R FILLER_226_107 ();
 DECAPx2_ASAP7_75t_R FILLER_226_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_143 ();
 DECAPx1_ASAP7_75t_R FILLER_226_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_156 ();
 DECAPx2_ASAP7_75t_R FILLER_226_163 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_169 ();
 DECAPx1_ASAP7_75t_R FILLER_226_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_182 ();
 FILLER_ASAP7_75t_R FILLER_226_186 ();
 FILLER_ASAP7_75t_R FILLER_226_195 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_204 ();
 FILLER_ASAP7_75t_R FILLER_226_213 ();
 DECAPx2_ASAP7_75t_R FILLER_226_221 ();
 DECAPx1_ASAP7_75t_R FILLER_226_233 ();
 DECAPx10_ASAP7_75t_R FILLER_226_240 ();
 DECAPx10_ASAP7_75t_R FILLER_226_262 ();
 DECAPx2_ASAP7_75t_R FILLER_226_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_290 ();
 DECAPx6_ASAP7_75t_R FILLER_226_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_313 ();
 DECAPx2_ASAP7_75t_R FILLER_226_322 ();
 FILLER_ASAP7_75t_R FILLER_226_335 ();
 FILLER_ASAP7_75t_R FILLER_226_344 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_349 ();
 DECAPx4_ASAP7_75t_R FILLER_226_360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_370 ();
 DECAPx2_ASAP7_75t_R FILLER_226_381 ();
 FILLER_ASAP7_75t_R FILLER_226_387 ();
 DECAPx6_ASAP7_75t_R FILLER_226_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_409 ();
 DECAPx10_ASAP7_75t_R FILLER_226_416 ();
 DECAPx10_ASAP7_75t_R FILLER_226_438 ();
 FILLER_ASAP7_75t_R FILLER_226_460 ();
 DECAPx2_ASAP7_75t_R FILLER_226_464 ();
 FILLER_ASAP7_75t_R FILLER_226_470 ();
 DECAPx6_ASAP7_75t_R FILLER_226_498 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_512 ();
 DECAPx1_ASAP7_75t_R FILLER_226_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_525 ();
 DECAPx6_ASAP7_75t_R FILLER_226_529 ();
 FILLER_ASAP7_75t_R FILLER_226_569 ();
 DECAPx2_ASAP7_75t_R FILLER_226_577 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_586 ();
 FILLER_ASAP7_75t_R FILLER_226_595 ();
 FILLER_ASAP7_75t_R FILLER_226_604 ();
 FILLER_ASAP7_75t_R FILLER_226_613 ();
 FILLER_ASAP7_75t_R FILLER_226_621 ();
 DECAPx6_ASAP7_75t_R FILLER_226_629 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_643 ();
 FILLER_ASAP7_75t_R FILLER_226_652 ();
 DECAPx6_ASAP7_75t_R FILLER_226_660 ();
 DECAPx1_ASAP7_75t_R FILLER_226_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_681 ();
 DECAPx10_ASAP7_75t_R FILLER_226_685 ();
 DECAPx10_ASAP7_75t_R FILLER_226_707 ();
 DECAPx1_ASAP7_75t_R FILLER_226_729 ();
 DECAPx10_ASAP7_75t_R FILLER_226_742 ();
 DECAPx10_ASAP7_75t_R FILLER_226_764 ();
 DECAPx1_ASAP7_75t_R FILLER_226_786 ();
 DECAPx4_ASAP7_75t_R FILLER_226_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_809 ();
 DECAPx2_ASAP7_75t_R FILLER_226_813 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_819 ();
 FILLER_ASAP7_75t_R FILLER_226_828 ();
 DECAPx6_ASAP7_75t_R FILLER_226_836 ();
 DECAPx1_ASAP7_75t_R FILLER_226_850 ();
 DECAPx4_ASAP7_75t_R FILLER_226_863 ();
 FILLER_ASAP7_75t_R FILLER_226_887 ();
 FILLER_ASAP7_75t_R FILLER_226_903 ();
 DECAPx10_ASAP7_75t_R FILLER_226_908 ();
 FILLER_ASAP7_75t_R FILLER_226_930 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_944 ();
 FILLER_ASAP7_75t_R FILLER_226_961 ();
 DECAPx6_ASAP7_75t_R FILLER_226_972 ();
 FILLER_ASAP7_75t_R FILLER_226_986 ();
 FILLER_ASAP7_75t_R FILLER_226_991 ();
 DECAPx1_ASAP7_75t_R FILLER_226_996 ();
 DECAPx6_ASAP7_75t_R FILLER_226_1014 ();
 FILLER_ASAP7_75t_R FILLER_226_1028 ();
 FILLER_ASAP7_75t_R FILLER_226_1036 ();
 DECAPx1_ASAP7_75t_R FILLER_226_1041 ();
 FILLER_ASAP7_75t_R FILLER_226_1048 ();
 DECAPx1_ASAP7_75t_R FILLER_226_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_1068 ();
 FILLER_ASAP7_75t_R FILLER_226_1073 ();
 FILLER_ASAP7_75t_R FILLER_226_1089 ();
 FILLER_ASAP7_75t_R FILLER_226_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_226_1341 ();
 DECAPx6_ASAP7_75t_R FILLER_226_1363 ();
 DECAPx2_ASAP7_75t_R FILLER_227_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_227_8 ();
 FILLER_ASAP7_75t_R FILLER_227_37 ();
 DECAPx10_ASAP7_75t_R FILLER_227_45 ();
 FILLER_ASAP7_75t_R FILLER_227_73 ();
 DECAPx6_ASAP7_75t_R FILLER_227_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_92 ();
 DECAPx6_ASAP7_75t_R FILLER_227_101 ();
 DECAPx1_ASAP7_75t_R FILLER_227_121 ();
 DECAPx2_ASAP7_75t_R FILLER_227_128 ();
 FILLER_ASAP7_75t_R FILLER_227_134 ();
 FILLER_ASAP7_75t_R FILLER_227_142 ();
 DECAPx2_ASAP7_75t_R FILLER_227_152 ();
 FILLER_ASAP7_75t_R FILLER_227_158 ();
 FILLER_ASAP7_75t_R FILLER_227_168 ();
 DECAPx2_ASAP7_75t_R FILLER_227_176 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_227_182 ();
 FILLER_ASAP7_75t_R FILLER_227_191 ();
 DECAPx2_ASAP7_75t_R FILLER_227_196 ();
 DECAPx6_ASAP7_75t_R FILLER_227_205 ();
 DECAPx1_ASAP7_75t_R FILLER_227_219 ();
 FILLER_ASAP7_75t_R FILLER_227_249 ();
 DECAPx4_ASAP7_75t_R FILLER_227_257 ();
 FILLER_ASAP7_75t_R FILLER_227_267 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_227_275 ();
 FILLER_ASAP7_75t_R FILLER_227_281 ();
 FILLER_ASAP7_75t_R FILLER_227_289 ();
 FILLER_ASAP7_75t_R FILLER_227_299 ();
 FILLER_ASAP7_75t_R FILLER_227_307 ();
 FILLER_ASAP7_75t_R FILLER_227_315 ();
 FILLER_ASAP7_75t_R FILLER_227_326 ();
 FILLER_ASAP7_75t_R FILLER_227_354 ();
 DECAPx4_ASAP7_75t_R FILLER_227_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_372 ();
 DECAPx6_ASAP7_75t_R FILLER_227_376 ();
 DECAPx2_ASAP7_75t_R FILLER_227_390 ();
 DECAPx1_ASAP7_75t_R FILLER_227_402 ();
 FILLER_ASAP7_75t_R FILLER_227_412 ();
 DECAPx4_ASAP7_75t_R FILLER_227_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_432 ();
 DECAPx2_ASAP7_75t_R FILLER_227_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_445 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_227_449 ();
 FILLER_ASAP7_75t_R FILLER_227_460 ();
 DECAPx2_ASAP7_75t_R FILLER_227_468 ();
 DECAPx2_ASAP7_75t_R FILLER_227_480 ();
 DECAPx2_ASAP7_75t_R FILLER_227_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_495 ();
 DECAPx2_ASAP7_75t_R FILLER_227_502 ();
 FILLER_ASAP7_75t_R FILLER_227_508 ();
 DECAPx2_ASAP7_75t_R FILLER_227_516 ();
 FILLER_ASAP7_75t_R FILLER_227_522 ();
 DECAPx6_ASAP7_75t_R FILLER_227_530 ();
 FILLER_ASAP7_75t_R FILLER_227_544 ();
 FILLER_ASAP7_75t_R FILLER_227_553 ();
 FILLER_ASAP7_75t_R FILLER_227_561 ();
 DECAPx4_ASAP7_75t_R FILLER_227_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_576 ();
 DECAPx6_ASAP7_75t_R FILLER_227_583 ();
 DECAPx2_ASAP7_75t_R FILLER_227_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_603 ();
 FILLER_ASAP7_75t_R FILLER_227_610 ();
 DECAPx4_ASAP7_75t_R FILLER_227_638 ();
 DECAPx2_ASAP7_75t_R FILLER_227_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_657 ();
 DECAPx10_ASAP7_75t_R FILLER_227_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_689 ();
 FILLER_ASAP7_75t_R FILLER_227_693 ();
 FILLER_ASAP7_75t_R FILLER_227_698 ();
 FILLER_ASAP7_75t_R FILLER_227_714 ();
 FILLER_ASAP7_75t_R FILLER_227_725 ();
 FILLER_ASAP7_75t_R FILLER_227_735 ();
 FILLER_ASAP7_75t_R FILLER_227_744 ();
 DECAPx2_ASAP7_75t_R FILLER_227_752 ();
 DECAPx2_ASAP7_75t_R FILLER_227_772 ();
 DECAPx6_ASAP7_75t_R FILLER_227_787 ();
 DECAPx2_ASAP7_75t_R FILLER_227_804 ();
 DECAPx6_ASAP7_75t_R FILLER_227_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_833 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_227_843 ();
 FILLER_ASAP7_75t_R FILLER_227_849 ();
 DECAPx6_ASAP7_75t_R FILLER_227_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_868 ();
 DECAPx6_ASAP7_75t_R FILLER_227_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_886 ();
 FILLER_ASAP7_75t_R FILLER_227_890 ();
 DECAPx6_ASAP7_75t_R FILLER_227_895 ();
 DECAPx1_ASAP7_75t_R FILLER_227_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_913 ();
 DECAPx1_ASAP7_75t_R FILLER_227_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_924 ();
 FILLER_ASAP7_75t_R FILLER_227_927 ();
 FILLER_ASAP7_75t_R FILLER_227_943 ();
 FILLER_ASAP7_75t_R FILLER_227_951 ();
 DECAPx1_ASAP7_75t_R FILLER_227_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_963 ();
 DECAPx2_ASAP7_75t_R FILLER_227_978 ();
 DECAPx6_ASAP7_75t_R FILLER_227_998 ();
 FILLER_ASAP7_75t_R FILLER_227_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1020 ();
 DECAPx4_ASAP7_75t_R FILLER_227_1042 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_227_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1058 ();
 FILLER_ASAP7_75t_R FILLER_227_1064 ();
 FILLER_ASAP7_75t_R FILLER_227_1080 ();
 DECAPx6_ASAP7_75t_R FILLER_227_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_227_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_227_1351 ();
 DECAPx1_ASAP7_75t_R FILLER_227_1373 ();
 DECAPx10_ASAP7_75t_R FILLER_228_2 ();
 FILLER_ASAP7_75t_R FILLER_228_24 ();
 DECAPx10_ASAP7_75t_R FILLER_228_29 ();
 DECAPx4_ASAP7_75t_R FILLER_228_51 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_61 ();
 DECAPx6_ASAP7_75t_R FILLER_228_70 ();
 FILLER_ASAP7_75t_R FILLER_228_92 ();
 FILLER_ASAP7_75t_R FILLER_228_100 ();
 DECAPx6_ASAP7_75t_R FILLER_228_108 ();
 DECAPx1_ASAP7_75t_R FILLER_228_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_126 ();
 DECAPx2_ASAP7_75t_R FILLER_228_133 ();
 FILLER_ASAP7_75t_R FILLER_228_145 ();
 DECAPx4_ASAP7_75t_R FILLER_228_150 ();
 DECAPx4_ASAP7_75t_R FILLER_228_168 ();
 FILLER_ASAP7_75t_R FILLER_228_204 ();
 FILLER_ASAP7_75t_R FILLER_228_212 ();
 DECAPx2_ASAP7_75t_R FILLER_228_217 ();
 FILLER_ASAP7_75t_R FILLER_228_223 ();
 DECAPx1_ASAP7_75t_R FILLER_228_231 ();
 FILLER_ASAP7_75t_R FILLER_228_261 ();
 FILLER_ASAP7_75t_R FILLER_228_289 ();
 DECAPx4_ASAP7_75t_R FILLER_228_297 ();
 DECAPx4_ASAP7_75t_R FILLER_228_313 ();
 FILLER_ASAP7_75t_R FILLER_228_323 ();
 FILLER_ASAP7_75t_R FILLER_228_331 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_339 ();
 DECAPx2_ASAP7_75t_R FILLER_228_345 ();
 DECAPx4_ASAP7_75t_R FILLER_228_357 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_367 ();
 FILLER_ASAP7_75t_R FILLER_228_376 ();
 DECAPx2_ASAP7_75t_R FILLER_228_381 ();
 FILLER_ASAP7_75t_R FILLER_228_387 ();
 DECAPx2_ASAP7_75t_R FILLER_228_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_421 ();
 DECAPx1_ASAP7_75t_R FILLER_228_448 ();
 FILLER_ASAP7_75t_R FILLER_228_460 ();
 DECAPx2_ASAP7_75t_R FILLER_228_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_470 ();
 DECAPx4_ASAP7_75t_R FILLER_228_477 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_487 ();
 FILLER_ASAP7_75t_R FILLER_228_498 ();
 DECAPx2_ASAP7_75t_R FILLER_228_526 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_532 ();
 FILLER_ASAP7_75t_R FILLER_228_541 ();
 FILLER_ASAP7_75t_R FILLER_228_554 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_563 ();
 FILLER_ASAP7_75t_R FILLER_228_572 ();
 DECAPx10_ASAP7_75t_R FILLER_228_600 ();
 DECAPx1_ASAP7_75t_R FILLER_228_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_626 ();
 FILLER_ASAP7_75t_R FILLER_228_630 ();
 DECAPx2_ASAP7_75t_R FILLER_228_635 ();
 FILLER_ASAP7_75t_R FILLER_228_641 ();
 FILLER_ASAP7_75t_R FILLER_228_657 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_662 ();
 DECAPx2_ASAP7_75t_R FILLER_228_668 ();
 FILLER_ASAP7_75t_R FILLER_228_674 ();
 DECAPx10_ASAP7_75t_R FILLER_228_685 ();
 DECAPx4_ASAP7_75t_R FILLER_228_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_717 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_732 ();
 FILLER_ASAP7_75t_R FILLER_228_741 ();
 DECAPx1_ASAP7_75t_R FILLER_228_749 ();
 FILLER_ASAP7_75t_R FILLER_228_767 ();
 FILLER_ASAP7_75t_R FILLER_228_775 ();
 DECAPx2_ASAP7_75t_R FILLER_228_780 ();
 DECAPx2_ASAP7_75t_R FILLER_228_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_795 ();
 DECAPx6_ASAP7_75t_R FILLER_228_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_819 ();
 DECAPx4_ASAP7_75t_R FILLER_228_823 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_833 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_850 ();
 FILLER_ASAP7_75t_R FILLER_228_867 ();
 FILLER_ASAP7_75t_R FILLER_228_878 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_883 ();
 DECAPx6_ASAP7_75t_R FILLER_228_889 ();
 DECAPx2_ASAP7_75t_R FILLER_228_903 ();
 DECAPx1_ASAP7_75t_R FILLER_228_921 ();
 DECAPx4_ASAP7_75t_R FILLER_228_932 ();
 DECAPx1_ASAP7_75t_R FILLER_228_948 ();
 DECAPx6_ASAP7_75t_R FILLER_228_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_975 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_979 ();
 DECAPx2_ASAP7_75t_R FILLER_228_996 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_1002 ();
 FILLER_ASAP7_75t_R FILLER_228_1011 ();
 DECAPx4_ASAP7_75t_R FILLER_228_1027 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1065 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_1087 ();
 DECAPx2_ASAP7_75t_R FILLER_228_1099 ();
 FILLER_ASAP7_75t_R FILLER_228_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_228_1355 ();
 DECAPx6_ASAP7_75t_R FILLER_229_2 ();
 DECAPx2_ASAP7_75t_R FILLER_229_16 ();
 DECAPx1_ASAP7_75t_R FILLER_229_28 ();
 DECAPx2_ASAP7_75t_R FILLER_229_38 ();
 DECAPx2_ASAP7_75t_R FILLER_229_47 ();
 DECAPx1_ASAP7_75t_R FILLER_229_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_83 ();
 DECAPx2_ASAP7_75t_R FILLER_229_92 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_98 ();
 DECAPx2_ASAP7_75t_R FILLER_229_107 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_113 ();
 DECAPx10_ASAP7_75t_R FILLER_229_142 ();
 FILLER_ASAP7_75t_R FILLER_229_170 ();
 FILLER_ASAP7_75t_R FILLER_229_178 ();
 DECAPx2_ASAP7_75t_R FILLER_229_186 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_192 ();
 DECAPx10_ASAP7_75t_R FILLER_229_221 ();
 DECAPx1_ASAP7_75t_R FILLER_229_243 ();
 FILLER_ASAP7_75t_R FILLER_229_253 ();
 DECAPx2_ASAP7_75t_R FILLER_229_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_264 ();
 DECAPx10_ASAP7_75t_R FILLER_229_271 ();
 DECAPx4_ASAP7_75t_R FILLER_229_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_303 ();
 DECAPx4_ASAP7_75t_R FILLER_229_312 ();
 FILLER_ASAP7_75t_R FILLER_229_322 ();
 DECAPx10_ASAP7_75t_R FILLER_229_330 ();
 DECAPx4_ASAP7_75t_R FILLER_229_352 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_388 ();
 DECAPx2_ASAP7_75t_R FILLER_229_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_403 ();
 DECAPx1_ASAP7_75t_R FILLER_229_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_411 ();
 DECAPx2_ASAP7_75t_R FILLER_229_420 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_426 ();
 FILLER_ASAP7_75t_R FILLER_229_435 ();
 DECAPx4_ASAP7_75t_R FILLER_229_440 ();
 FILLER_ASAP7_75t_R FILLER_229_456 ();
 FILLER_ASAP7_75t_R FILLER_229_464 ();
 DECAPx4_ASAP7_75t_R FILLER_229_492 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_502 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_511 ();
 FILLER_ASAP7_75t_R FILLER_229_517 ();
 FILLER_ASAP7_75t_R FILLER_229_525 ();
 FILLER_ASAP7_75t_R FILLER_229_535 ();
 FILLER_ASAP7_75t_R FILLER_229_543 ();
 FILLER_ASAP7_75t_R FILLER_229_552 ();
 FILLER_ASAP7_75t_R FILLER_229_562 ();
 DECAPx1_ASAP7_75t_R FILLER_229_571 ();
 DECAPx2_ASAP7_75t_R FILLER_229_581 ();
 FILLER_ASAP7_75t_R FILLER_229_587 ();
 DECAPx6_ASAP7_75t_R FILLER_229_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_606 ();
 DECAPx6_ASAP7_75t_R FILLER_229_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_627 ();
 DECAPx10_ASAP7_75t_R FILLER_229_636 ();
 DECAPx2_ASAP7_75t_R FILLER_229_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_664 ();
 DECAPx2_ASAP7_75t_R FILLER_229_679 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_685 ();
 FILLER_ASAP7_75t_R FILLER_229_702 ();
 DECAPx6_ASAP7_75t_R FILLER_229_707 ();
 DECAPx1_ASAP7_75t_R FILLER_229_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_725 ();
 DECAPx10_ASAP7_75t_R FILLER_229_735 ();
 FILLER_ASAP7_75t_R FILLER_229_757 ();
 FILLER_ASAP7_75t_R FILLER_229_765 ();
 DECAPx6_ASAP7_75t_R FILLER_229_773 ();
 FILLER_ASAP7_75t_R FILLER_229_787 ();
 DECAPx10_ASAP7_75t_R FILLER_229_792 ();
 DECAPx10_ASAP7_75t_R FILLER_229_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_836 ();
 DECAPx6_ASAP7_75t_R FILLER_229_846 ();
 DECAPx2_ASAP7_75t_R FILLER_229_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_866 ();
 DECAPx10_ASAP7_75t_R FILLER_229_870 ();
 DECAPx1_ASAP7_75t_R FILLER_229_892 ();
 DECAPx2_ASAP7_75t_R FILLER_229_905 ();
 FILLER_ASAP7_75t_R FILLER_229_911 ();
 DECAPx1_ASAP7_75t_R FILLER_229_921 ();
 FILLER_ASAP7_75t_R FILLER_229_927 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_938 ();
 FILLER_ASAP7_75t_R FILLER_229_951 ();
 DECAPx6_ASAP7_75t_R FILLER_229_959 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_973 ();
 DECAPx10_ASAP7_75t_R FILLER_229_979 ();
 DECAPx2_ASAP7_75t_R FILLER_229_1001 ();
 FILLER_ASAP7_75t_R FILLER_229_1007 ();
 DECAPx4_ASAP7_75t_R FILLER_229_1012 ();
 FILLER_ASAP7_75t_R FILLER_229_1022 ();
 FILLER_ASAP7_75t_R FILLER_229_1027 ();
 DECAPx6_ASAP7_75t_R FILLER_229_1043 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_1061 ();
 FILLER_ASAP7_75t_R FILLER_229_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1070 ();
 DECAPx1_ASAP7_75t_R FILLER_229_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1264 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1286 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1308 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_229_1352 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_1374 ();
 DECAPx6_ASAP7_75t_R FILLER_230_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_16 ();
 DECAPx1_ASAP7_75t_R FILLER_230_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_49 ();
 FILLER_ASAP7_75t_R FILLER_230_58 ();
 FILLER_ASAP7_75t_R FILLER_230_66 ();
 DECAPx2_ASAP7_75t_R FILLER_230_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_77 ();
 FILLER_ASAP7_75t_R FILLER_230_84 ();
 DECAPx2_ASAP7_75t_R FILLER_230_92 ();
 FILLER_ASAP7_75t_R FILLER_230_98 ();
 DECAPx4_ASAP7_75t_R FILLER_230_108 ();
 FILLER_ASAP7_75t_R FILLER_230_118 ();
 DECAPx1_ASAP7_75t_R FILLER_230_126 ();
 DECAPx2_ASAP7_75t_R FILLER_230_133 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_139 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_148 ();
 FILLER_ASAP7_75t_R FILLER_230_157 ();
 DECAPx4_ASAP7_75t_R FILLER_230_162 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_172 ();
 DECAPx1_ASAP7_75t_R FILLER_230_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_185 ();
 DECAPx6_ASAP7_75t_R FILLER_230_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_203 ();
 DECAPx1_ASAP7_75t_R FILLER_230_210 ();
 DECAPx6_ASAP7_75t_R FILLER_230_240 ();
 DECAPx2_ASAP7_75t_R FILLER_230_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_293 ();
 DECAPx2_ASAP7_75t_R FILLER_230_299 ();
 FILLER_ASAP7_75t_R FILLER_230_305 ();
 DECAPx2_ASAP7_75t_R FILLER_230_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_321 ();
 DECAPx6_ASAP7_75t_R FILLER_230_348 ();
 FILLER_ASAP7_75t_R FILLER_230_362 ();
 DECAPx2_ASAP7_75t_R FILLER_230_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_376 ();
 DECAPx10_ASAP7_75t_R FILLER_230_383 ();
 DECAPx1_ASAP7_75t_R FILLER_230_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_409 ();
 DECAPx10_ASAP7_75t_R FILLER_230_413 ();
 DECAPx10_ASAP7_75t_R FILLER_230_435 ();
 DECAPx1_ASAP7_75t_R FILLER_230_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_461 ();
 DECAPx4_ASAP7_75t_R FILLER_230_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_474 ();
 FILLER_ASAP7_75t_R FILLER_230_481 ();
 DECAPx10_ASAP7_75t_R FILLER_230_486 ();
 DECAPx6_ASAP7_75t_R FILLER_230_508 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_522 ();
 DECAPx2_ASAP7_75t_R FILLER_230_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_539 ();
 FILLER_ASAP7_75t_R FILLER_230_547 ();
 DECAPx1_ASAP7_75t_R FILLER_230_560 ();
 DECAPx2_ASAP7_75t_R FILLER_230_590 ();
 FILLER_ASAP7_75t_R FILLER_230_596 ();
 DECAPx2_ASAP7_75t_R FILLER_230_624 ();
 DECAPx2_ASAP7_75t_R FILLER_230_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_642 ();
 FILLER_ASAP7_75t_R FILLER_230_649 ();
 DECAPx2_ASAP7_75t_R FILLER_230_657 ();
 DECAPx4_ASAP7_75t_R FILLER_230_677 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_687 ();
 DECAPx10_ASAP7_75t_R FILLER_230_704 ();
 DECAPx10_ASAP7_75t_R FILLER_230_726 ();
 DECAPx4_ASAP7_75t_R FILLER_230_748 ();
 FILLER_ASAP7_75t_R FILLER_230_758 ();
 DECAPx4_ASAP7_75t_R FILLER_230_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_773 ();
 DECAPx6_ASAP7_75t_R FILLER_230_777 ();
 FILLER_ASAP7_75t_R FILLER_230_791 ();
 FILLER_ASAP7_75t_R FILLER_230_807 ();
 FILLER_ASAP7_75t_R FILLER_230_815 ();
 DECAPx2_ASAP7_75t_R FILLER_230_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_829 ();
 FILLER_ASAP7_75t_R FILLER_230_839 ();
 DECAPx6_ASAP7_75t_R FILLER_230_844 ();
 DECAPx1_ASAP7_75t_R FILLER_230_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_862 ();
 FILLER_ASAP7_75t_R FILLER_230_866 ();
 DECAPx6_ASAP7_75t_R FILLER_230_871 ();
 DECAPx1_ASAP7_75t_R FILLER_230_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_889 ();
 FILLER_ASAP7_75t_R FILLER_230_904 ();
 DECAPx1_ASAP7_75t_R FILLER_230_913 ();
 FILLER_ASAP7_75t_R FILLER_230_923 ();
 DECAPx10_ASAP7_75t_R FILLER_230_931 ();
 DECAPx1_ASAP7_75t_R FILLER_230_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_971 ();
 DECAPx2_ASAP7_75t_R FILLER_230_986 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_992 ();
 DECAPx2_ASAP7_75t_R FILLER_230_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1004 ();
 DECAPx6_ASAP7_75t_R FILLER_230_1019 ();
 FILLER_ASAP7_75t_R FILLER_230_1033 ();
 FILLER_ASAP7_75t_R FILLER_230_1038 ();
 FILLER_ASAP7_75t_R FILLER_230_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_230_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1083 ();
 FILLER_ASAP7_75t_R FILLER_230_1087 ();
 FILLER_ASAP7_75t_R FILLER_230_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1174 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_230_1350 ();
 DECAPx1_ASAP7_75t_R FILLER_230_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_231_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_16 ();
 DECAPx2_ASAP7_75t_R FILLER_231_25 ();
 FILLER_ASAP7_75t_R FILLER_231_31 ();
 DECAPx2_ASAP7_75t_R FILLER_231_36 ();
 FILLER_ASAP7_75t_R FILLER_231_48 ();
 DECAPx10_ASAP7_75t_R FILLER_231_58 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_80 ();
 DECAPx6_ASAP7_75t_R FILLER_231_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_100 ();
 DECAPx2_ASAP7_75t_R FILLER_231_109 ();
 FILLER_ASAP7_75t_R FILLER_231_115 ();
 DECAPx6_ASAP7_75t_R FILLER_231_123 ();
 DECAPx2_ASAP7_75t_R FILLER_231_163 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_169 ();
 DECAPx6_ASAP7_75t_R FILLER_231_198 ();
 DECAPx2_ASAP7_75t_R FILLER_231_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_218 ();
 FILLER_ASAP7_75t_R FILLER_231_225 ();
 FILLER_ASAP7_75t_R FILLER_231_233 ();
 FILLER_ASAP7_75t_R FILLER_231_238 ();
 FILLER_ASAP7_75t_R FILLER_231_243 ();
 FILLER_ASAP7_75t_R FILLER_231_251 ();
 DECAPx2_ASAP7_75t_R FILLER_231_261 ();
 FILLER_ASAP7_75t_R FILLER_231_267 ();
 FILLER_ASAP7_75t_R FILLER_231_275 ();
 FILLER_ASAP7_75t_R FILLER_231_283 ();
 FILLER_ASAP7_75t_R FILLER_231_311 ();
 DECAPx4_ASAP7_75t_R FILLER_231_319 ();
 FILLER_ASAP7_75t_R FILLER_231_335 ();
 DECAPx2_ASAP7_75t_R FILLER_231_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_346 ();
 DECAPx2_ASAP7_75t_R FILLER_231_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_356 ();
 DECAPx6_ASAP7_75t_R FILLER_231_363 ();
 FILLER_ASAP7_75t_R FILLER_231_385 ();
 DECAPx1_ASAP7_75t_R FILLER_231_394 ();
 DECAPx1_ASAP7_75t_R FILLER_231_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_408 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_435 ();
 DECAPx1_ASAP7_75t_R FILLER_231_444 ();
 DECAPx2_ASAP7_75t_R FILLER_231_474 ();
 FILLER_ASAP7_75t_R FILLER_231_480 ();
 DECAPx6_ASAP7_75t_R FILLER_231_490 ();
 DECAPx2_ASAP7_75t_R FILLER_231_504 ();
 DECAPx1_ASAP7_75t_R FILLER_231_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_520 ();
 DECAPx2_ASAP7_75t_R FILLER_231_524 ();
 FILLER_ASAP7_75t_R FILLER_231_530 ();
 DECAPx1_ASAP7_75t_R FILLER_231_538 ();
 DECAPx6_ASAP7_75t_R FILLER_231_550 ();
 DECAPx2_ASAP7_75t_R FILLER_231_564 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_576 ();
 DECAPx2_ASAP7_75t_R FILLER_231_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_588 ();
 DECAPx4_ASAP7_75t_R FILLER_231_592 ();
 DECAPx1_ASAP7_75t_R FILLER_231_608 ();
 FILLER_ASAP7_75t_R FILLER_231_615 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_625 ();
 DECAPx4_ASAP7_75t_R FILLER_231_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_644 ();
 FILLER_ASAP7_75t_R FILLER_231_659 ();
 DECAPx2_ASAP7_75t_R FILLER_231_667 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_673 ();
 DECAPx6_ASAP7_75t_R FILLER_231_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_696 ();
 FILLER_ASAP7_75t_R FILLER_231_700 ();
 DECAPx1_ASAP7_75t_R FILLER_231_716 ();
 DECAPx2_ASAP7_75t_R FILLER_231_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_737 ();
 FILLER_ASAP7_75t_R FILLER_231_746 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_756 ();
 FILLER_ASAP7_75t_R FILLER_231_765 ();
 DECAPx1_ASAP7_75t_R FILLER_231_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_777 ();
 FILLER_ASAP7_75t_R FILLER_231_784 ();
 FILLER_ASAP7_75t_R FILLER_231_792 ();
 DECAPx4_ASAP7_75t_R FILLER_231_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_807 ();
 DECAPx1_ASAP7_75t_R FILLER_231_822 ();
 FILLER_ASAP7_75t_R FILLER_231_832 ();
 DECAPx10_ASAP7_75t_R FILLER_231_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_859 ();
 DECAPx4_ASAP7_75t_R FILLER_231_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_876 ();
 DECAPx4_ASAP7_75t_R FILLER_231_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_893 ();
 DECAPx6_ASAP7_75t_R FILLER_231_897 ();
 DECAPx1_ASAP7_75t_R FILLER_231_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_924 ();
 DECAPx4_ASAP7_75t_R FILLER_231_927 ();
 DECAPx6_ASAP7_75t_R FILLER_231_946 ();
 FILLER_ASAP7_75t_R FILLER_231_960 ();
 FILLER_ASAP7_75t_R FILLER_231_965 ();
 DECAPx10_ASAP7_75t_R FILLER_231_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1003 ();
 FILLER_ASAP7_75t_R FILLER_231_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1023 ();
 FILLER_ASAP7_75t_R FILLER_231_1035 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1043 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_231_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_231_1343 ();
 DECAPx4_ASAP7_75t_R FILLER_231_1365 ();
 FILLER_ASAP7_75t_R FILLER_231_1375 ();
 DECAPx4_ASAP7_75t_R FILLER_232_2 ();
 DECAPx2_ASAP7_75t_R FILLER_232_38 ();
 FILLER_ASAP7_75t_R FILLER_232_44 ();
 DECAPx6_ASAP7_75t_R FILLER_232_52 ();
 DECAPx1_ASAP7_75t_R FILLER_232_66 ();
 FILLER_ASAP7_75t_R FILLER_232_76 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_84 ();
 DECAPx4_ASAP7_75t_R FILLER_232_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_103 ();
 DECAPx1_ASAP7_75t_R FILLER_232_110 ();
 DECAPx4_ASAP7_75t_R FILLER_232_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_150 ();
 DECAPx6_ASAP7_75t_R FILLER_232_154 ();
 DECAPx2_ASAP7_75t_R FILLER_232_168 ();
 DECAPx4_ASAP7_75t_R FILLER_232_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_190 ();
 DECAPx6_ASAP7_75t_R FILLER_232_197 ();
 DECAPx1_ASAP7_75t_R FILLER_232_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_215 ();
 FILLER_ASAP7_75t_R FILLER_232_222 ();
 DECAPx6_ASAP7_75t_R FILLER_232_227 ();
 DECAPx1_ASAP7_75t_R FILLER_232_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_245 ();
 DECAPx2_ASAP7_75t_R FILLER_232_254 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_266 ();
 DECAPx2_ASAP7_75t_R FILLER_232_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_281 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_285 ();
 DECAPx2_ASAP7_75t_R FILLER_232_294 ();
 FILLER_ASAP7_75t_R FILLER_232_303 ();
 DECAPx6_ASAP7_75t_R FILLER_232_311 ();
 DECAPx2_ASAP7_75t_R FILLER_232_325 ();
 DECAPx2_ASAP7_75t_R FILLER_232_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_343 ();
 FILLER_ASAP7_75t_R FILLER_232_350 ();
 FILLER_ASAP7_75t_R FILLER_232_360 ();
 FILLER_ASAP7_75t_R FILLER_232_370 ();
 DECAPx4_ASAP7_75t_R FILLER_232_378 ();
 FILLER_ASAP7_75t_R FILLER_232_388 ();
 FILLER_ASAP7_75t_R FILLER_232_416 ();
 DECAPx1_ASAP7_75t_R FILLER_232_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_428 ();
 DECAPx2_ASAP7_75t_R FILLER_232_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_461 ();
 FILLER_ASAP7_75t_R FILLER_232_464 ();
 DECAPx1_ASAP7_75t_R FILLER_232_472 ();
 FILLER_ASAP7_75t_R FILLER_232_482 ();
 DECAPx2_ASAP7_75t_R FILLER_232_492 ();
 DECAPx2_ASAP7_75t_R FILLER_232_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_530 ();
 DECAPx10_ASAP7_75t_R FILLER_232_539 ();
 DECAPx10_ASAP7_75t_R FILLER_232_561 ();
 DECAPx4_ASAP7_75t_R FILLER_232_583 ();
 DECAPx6_ASAP7_75t_R FILLER_232_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_615 ();
 DECAPx1_ASAP7_75t_R FILLER_232_622 ();
 DECAPx4_ASAP7_75t_R FILLER_232_632 ();
 FILLER_ASAP7_75t_R FILLER_232_642 ();
 DECAPx4_ASAP7_75t_R FILLER_232_658 ();
 FILLER_ASAP7_75t_R FILLER_232_668 ();
 FILLER_ASAP7_75t_R FILLER_232_684 ();
 FILLER_ASAP7_75t_R FILLER_232_692 ();
 DECAPx2_ASAP7_75t_R FILLER_232_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_703 ();
 DECAPx2_ASAP7_75t_R FILLER_232_707 ();
 FILLER_ASAP7_75t_R FILLER_232_713 ();
 DECAPx6_ASAP7_75t_R FILLER_232_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_738 ();
 DECAPx4_ASAP7_75t_R FILLER_232_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_756 ();
 DECAPx2_ASAP7_75t_R FILLER_232_771 ();
 FILLER_ASAP7_75t_R FILLER_232_777 ();
 DECAPx6_ASAP7_75t_R FILLER_232_793 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_807 ();
 DECAPx2_ASAP7_75t_R FILLER_232_816 ();
 DECAPx10_ASAP7_75t_R FILLER_232_825 ();
 FILLER_ASAP7_75t_R FILLER_232_847 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_855 ();
 DECAPx2_ASAP7_75t_R FILLER_232_864 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_870 ();
 FILLER_ASAP7_75t_R FILLER_232_887 ();
 DECAPx6_ASAP7_75t_R FILLER_232_892 ();
 DECAPx6_ASAP7_75t_R FILLER_232_920 ();
 DECAPx1_ASAP7_75t_R FILLER_232_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_938 ();
 DECAPx4_ASAP7_75t_R FILLER_232_953 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_963 ();
 DECAPx6_ASAP7_75t_R FILLER_232_969 ();
 FILLER_ASAP7_75t_R FILLER_232_986 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_232_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_232_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_1052 ();
 FILLER_ASAP7_75t_R FILLER_232_1056 ();
 FILLER_ASAP7_75t_R FILLER_232_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_232_1066 ();
 DECAPx4_ASAP7_75t_R FILLER_232_1075 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_232_1355 ();
 DECAPx4_ASAP7_75t_R FILLER_233_2 ();
 FILLER_ASAP7_75t_R FILLER_233_12 ();
 DECAPx2_ASAP7_75t_R FILLER_233_20 ();
 DECAPx10_ASAP7_75t_R FILLER_233_29 ();
 DECAPx6_ASAP7_75t_R FILLER_233_51 ();
 FILLER_ASAP7_75t_R FILLER_233_65 ();
 DECAPx4_ASAP7_75t_R FILLER_233_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_103 ();
 DECAPx2_ASAP7_75t_R FILLER_233_110 ();
 DECAPx2_ASAP7_75t_R FILLER_233_122 ();
 DECAPx2_ASAP7_75t_R FILLER_233_131 ();
 DECAPx6_ASAP7_75t_R FILLER_233_143 ();
 DECAPx2_ASAP7_75t_R FILLER_233_157 ();
 DECAPx2_ASAP7_75t_R FILLER_233_169 ();
 FILLER_ASAP7_75t_R FILLER_233_175 ();
 FILLER_ASAP7_75t_R FILLER_233_203 ();
 FILLER_ASAP7_75t_R FILLER_233_231 ();
 DECAPx10_ASAP7_75t_R FILLER_233_239 ();
 DECAPx10_ASAP7_75t_R FILLER_233_261 ();
 DECAPx10_ASAP7_75t_R FILLER_233_283 ();
 DECAPx6_ASAP7_75t_R FILLER_233_305 ();
 DECAPx2_ASAP7_75t_R FILLER_233_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_325 ();
 FILLER_ASAP7_75t_R FILLER_233_352 ();
 DECAPx6_ASAP7_75t_R FILLER_233_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_374 ();
 DECAPx4_ASAP7_75t_R FILLER_233_383 ();
 DECAPx1_ASAP7_75t_R FILLER_233_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_403 ();
 DECAPx4_ASAP7_75t_R FILLER_233_407 ();
 FILLER_ASAP7_75t_R FILLER_233_417 ();
 FILLER_ASAP7_75t_R FILLER_233_425 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_233_430 ();
 DECAPx1_ASAP7_75t_R FILLER_233_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_443 ();
 DECAPx2_ASAP7_75t_R FILLER_233_447 ();
 DECAPx1_ASAP7_75t_R FILLER_233_459 ();
 DECAPx2_ASAP7_75t_R FILLER_233_466 ();
 FILLER_ASAP7_75t_R FILLER_233_472 ();
 DECAPx1_ASAP7_75t_R FILLER_233_477 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_233_487 ();
 DECAPx2_ASAP7_75t_R FILLER_233_496 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_233_502 ();
 FILLER_ASAP7_75t_R FILLER_233_511 ();
 DECAPx4_ASAP7_75t_R FILLER_233_516 ();
 FILLER_ASAP7_75t_R FILLER_233_532 ();
 DECAPx2_ASAP7_75t_R FILLER_233_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_548 ();
 FILLER_ASAP7_75t_R FILLER_233_575 ();
 DECAPx1_ASAP7_75t_R FILLER_233_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_587 ();
 FILLER_ASAP7_75t_R FILLER_233_594 ();
 FILLER_ASAP7_75t_R FILLER_233_604 ();
 DECAPx1_ASAP7_75t_R FILLER_233_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_616 ();
 DECAPx2_ASAP7_75t_R FILLER_233_623 ();
 DECAPx10_ASAP7_75t_R FILLER_233_635 ();
 DECAPx1_ASAP7_75t_R FILLER_233_657 ();
 DECAPx4_ASAP7_75t_R FILLER_233_664 ();
 FILLER_ASAP7_75t_R FILLER_233_674 ();
 DECAPx10_ASAP7_75t_R FILLER_233_682 ();
 DECAPx6_ASAP7_75t_R FILLER_233_704 ();
 DECAPx4_ASAP7_75t_R FILLER_233_724 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_233_734 ();
 FILLER_ASAP7_75t_R FILLER_233_743 ();
 DECAPx2_ASAP7_75t_R FILLER_233_751 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_233_757 ();
 DECAPx4_ASAP7_75t_R FILLER_233_766 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_233_776 ();
 DECAPx6_ASAP7_75t_R FILLER_233_785 ();
 DECAPx2_ASAP7_75t_R FILLER_233_799 ();
 DECAPx10_ASAP7_75t_R FILLER_233_811 ();
 FILLER_ASAP7_75t_R FILLER_233_833 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_233_841 ();
 DECAPx1_ASAP7_75t_R FILLER_233_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_854 ();
 DECAPx4_ASAP7_75t_R FILLER_233_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_879 ();
 DECAPx10_ASAP7_75t_R FILLER_233_883 ();
 DECAPx4_ASAP7_75t_R FILLER_233_905 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_233_915 ();
 DECAPx1_ASAP7_75t_R FILLER_233_921 ();
 FILLER_ASAP7_75t_R FILLER_233_927 ();
 DECAPx4_ASAP7_75t_R FILLER_233_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_953 ();
 DECAPx6_ASAP7_75t_R FILLER_233_968 ();
 DECAPx1_ASAP7_75t_R FILLER_233_982 ();
 FILLER_ASAP7_75t_R FILLER_233_1000 ();
 DECAPx2_ASAP7_75t_R FILLER_233_1012 ();
 DECAPx4_ASAP7_75t_R FILLER_233_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1059 ();
 DECAPx4_ASAP7_75t_R FILLER_233_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_233_1337 ();
 DECAPx6_ASAP7_75t_R FILLER_233_1359 ();
 DECAPx1_ASAP7_75t_R FILLER_233_1373 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_2 ();
 DECAPx2_ASAP7_75t_R FILLER_234_31 ();
 DECAPx2_ASAP7_75t_R FILLER_234_43 ();
 FILLER_ASAP7_75t_R FILLER_234_55 ();
 DECAPx6_ASAP7_75t_R FILLER_234_65 ();
 FILLER_ASAP7_75t_R FILLER_234_79 ();
 DECAPx4_ASAP7_75t_R FILLER_234_84 ();
 FILLER_ASAP7_75t_R FILLER_234_94 ();
 DECAPx6_ASAP7_75t_R FILLER_234_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_132 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_159 ();
 FILLER_ASAP7_75t_R FILLER_234_170 ();
 DECAPx2_ASAP7_75t_R FILLER_234_178 ();
 FILLER_ASAP7_75t_R FILLER_234_184 ();
 FILLER_ASAP7_75t_R FILLER_234_192 ();
 DECAPx2_ASAP7_75t_R FILLER_234_197 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_206 ();
 DECAPx2_ASAP7_75t_R FILLER_234_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_221 ();
 DECAPx2_ASAP7_75t_R FILLER_234_248 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_254 ();
 DECAPx2_ASAP7_75t_R FILLER_234_265 ();
 FILLER_ASAP7_75t_R FILLER_234_271 ();
 DECAPx4_ASAP7_75t_R FILLER_234_279 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_289 ();
 DECAPx2_ASAP7_75t_R FILLER_234_298 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_310 ();
 DECAPx4_ASAP7_75t_R FILLER_234_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_326 ();
 DECAPx2_ASAP7_75t_R FILLER_234_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_339 ();
 DECAPx10_ASAP7_75t_R FILLER_234_343 ();
 DECAPx2_ASAP7_75t_R FILLER_234_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_371 ();
 FILLER_ASAP7_75t_R FILLER_234_380 ();
 DECAPx10_ASAP7_75t_R FILLER_234_388 ();
 DECAPx10_ASAP7_75t_R FILLER_234_410 ();
 DECAPx10_ASAP7_75t_R FILLER_234_432 ();
 DECAPx2_ASAP7_75t_R FILLER_234_454 ();
 FILLER_ASAP7_75t_R FILLER_234_460 ();
 DECAPx10_ASAP7_75t_R FILLER_234_464 ();
 DECAPx10_ASAP7_75t_R FILLER_234_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_508 ();
 DECAPx4_ASAP7_75t_R FILLER_234_515 ();
 FILLER_ASAP7_75t_R FILLER_234_525 ();
 DECAPx2_ASAP7_75t_R FILLER_234_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_536 ();
 DECAPx4_ASAP7_75t_R FILLER_234_543 ();
 DECAPx1_ASAP7_75t_R FILLER_234_559 ();
 FILLER_ASAP7_75t_R FILLER_234_566 ();
 FILLER_ASAP7_75t_R FILLER_234_594 ();
 DECAPx4_ASAP7_75t_R FILLER_234_602 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_612 ();
 DECAPx2_ASAP7_75t_R FILLER_234_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_627 ();
 DECAPx2_ASAP7_75t_R FILLER_234_637 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_643 ();
 FILLER_ASAP7_75t_R FILLER_234_649 ();
 DECAPx10_ASAP7_75t_R FILLER_234_660 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_682 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_688 ();
 DECAPx6_ASAP7_75t_R FILLER_234_700 ();
 FILLER_ASAP7_75t_R FILLER_234_717 ();
 DECAPx4_ASAP7_75t_R FILLER_234_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_738 ();
 DECAPx1_ASAP7_75t_R FILLER_234_742 ();
 DECAPx10_ASAP7_75t_R FILLER_234_758 ();
 DECAPx10_ASAP7_75t_R FILLER_234_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_802 ();
 FILLER_ASAP7_75t_R FILLER_234_809 ();
 DECAPx2_ASAP7_75t_R FILLER_234_817 ();
 FILLER_ASAP7_75t_R FILLER_234_823 ();
 DECAPx2_ASAP7_75t_R FILLER_234_831 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_837 ();
 DECAPx4_ASAP7_75t_R FILLER_234_854 ();
 FILLER_ASAP7_75t_R FILLER_234_864 ();
 DECAPx2_ASAP7_75t_R FILLER_234_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_875 ();
 DECAPx1_ASAP7_75t_R FILLER_234_890 ();
 FILLER_ASAP7_75t_R FILLER_234_900 ();
 FILLER_ASAP7_75t_R FILLER_234_908 ();
 DECAPx1_ASAP7_75t_R FILLER_234_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_917 ();
 DECAPx1_ASAP7_75t_R FILLER_234_932 ();
 DECAPx4_ASAP7_75t_R FILLER_234_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_949 ();
 FILLER_ASAP7_75t_R FILLER_234_953 ();
 FILLER_ASAP7_75t_R FILLER_234_958 ();
 DECAPx2_ASAP7_75t_R FILLER_234_974 ();
 FILLER_ASAP7_75t_R FILLER_234_980 ();
 DECAPx2_ASAP7_75t_R FILLER_234_985 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_991 ();
 FILLER_ASAP7_75t_R FILLER_234_997 ();
 DECAPx4_ASAP7_75t_R FILLER_234_1002 ();
 FILLER_ASAP7_75t_R FILLER_234_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1017 ();
 DECAPx6_ASAP7_75t_R FILLER_234_1039 ();
 FILLER_ASAP7_75t_R FILLER_234_1053 ();
 FILLER_ASAP7_75t_R FILLER_234_1058 ();
 FILLER_ASAP7_75t_R FILLER_234_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_234_1068 ();
 FILLER_ASAP7_75t_R FILLER_234_1075 ();
 FILLER_ASAP7_75t_R FILLER_234_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_234_1338 ();
 DECAPx6_ASAP7_75t_R FILLER_234_1360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_1374 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_2 ();
 FILLER_ASAP7_75t_R FILLER_235_11 ();
 DECAPx1_ASAP7_75t_R FILLER_235_19 ();
 FILLER_ASAP7_75t_R FILLER_235_26 ();
 FILLER_ASAP7_75t_R FILLER_235_54 ();
 DECAPx2_ASAP7_75t_R FILLER_235_64 ();
 DECAPx6_ASAP7_75t_R FILLER_235_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_90 ();
 FILLER_ASAP7_75t_R FILLER_235_101 ();
 FILLER_ASAP7_75t_R FILLER_235_109 ();
 DECAPx2_ASAP7_75t_R FILLER_235_114 ();
 DECAPx6_ASAP7_75t_R FILLER_235_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_140 ();
 FILLER_ASAP7_75t_R FILLER_235_147 ();
 DECAPx6_ASAP7_75t_R FILLER_235_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_185 ();
 DECAPx10_ASAP7_75t_R FILLER_235_192 ();
 DECAPx6_ASAP7_75t_R FILLER_235_214 ();
 DECAPx2_ASAP7_75t_R FILLER_235_228 ();
 DECAPx1_ASAP7_75t_R FILLER_235_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_244 ();
 FILLER_ASAP7_75t_R FILLER_235_248 ();
 DECAPx1_ASAP7_75t_R FILLER_235_256 ();
 DECAPx2_ASAP7_75t_R FILLER_235_266 ();
 FILLER_ASAP7_75t_R FILLER_235_272 ();
 DECAPx1_ASAP7_75t_R FILLER_235_280 ();
 FILLER_ASAP7_75t_R FILLER_235_287 ();
 FILLER_ASAP7_75t_R FILLER_235_315 ();
 DECAPx10_ASAP7_75t_R FILLER_235_323 ();
 DECAPx4_ASAP7_75t_R FILLER_235_345 ();
 FILLER_ASAP7_75t_R FILLER_235_355 ();
 DECAPx4_ASAP7_75t_R FILLER_235_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_373 ();
 DECAPx10_ASAP7_75t_R FILLER_235_380 ();
 FILLER_ASAP7_75t_R FILLER_235_402 ();
 DECAPx4_ASAP7_75t_R FILLER_235_410 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_420 ();
 DECAPx4_ASAP7_75t_R FILLER_235_429 ();
 FILLER_ASAP7_75t_R FILLER_235_439 ();
 DECAPx1_ASAP7_75t_R FILLER_235_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_451 ();
 DECAPx10_ASAP7_75t_R FILLER_235_455 ();
 FILLER_ASAP7_75t_R FILLER_235_477 ();
 FILLER_ASAP7_75t_R FILLER_235_487 ();
 DECAPx2_ASAP7_75t_R FILLER_235_495 ();
 DECAPx10_ASAP7_75t_R FILLER_235_527 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_549 ();
 DECAPx6_ASAP7_75t_R FILLER_235_558 ();
 DECAPx1_ASAP7_75t_R FILLER_235_572 ();
 FILLER_ASAP7_75t_R FILLER_235_582 ();
 DECAPx10_ASAP7_75t_R FILLER_235_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_609 ();
 DECAPx10_ASAP7_75t_R FILLER_235_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_658 ();
 DECAPx1_ASAP7_75t_R FILLER_235_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_666 ();
 FILLER_ASAP7_75t_R FILLER_235_681 ();
 FILLER_ASAP7_75t_R FILLER_235_692 ();
 DECAPx2_ASAP7_75t_R FILLER_235_697 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_703 ();
 DECAPx2_ASAP7_75t_R FILLER_235_720 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_726 ();
 FILLER_ASAP7_75t_R FILLER_235_738 ();
 DECAPx4_ASAP7_75t_R FILLER_235_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_764 ();
 DECAPx2_ASAP7_75t_R FILLER_235_771 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_777 ();
 FILLER_ASAP7_75t_R FILLER_235_786 ();
 DECAPx2_ASAP7_75t_R FILLER_235_797 ();
 DECAPx4_ASAP7_75t_R FILLER_235_817 ();
 DECAPx6_ASAP7_75t_R FILLER_235_841 ();
 DECAPx1_ASAP7_75t_R FILLER_235_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_859 ();
 DECAPx10_ASAP7_75t_R FILLER_235_863 ();
 DECAPx2_ASAP7_75t_R FILLER_235_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_891 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_906 ();
 FILLER_ASAP7_75t_R FILLER_235_923 ();
 FILLER_ASAP7_75t_R FILLER_235_927 ();
 FILLER_ASAP7_75t_R FILLER_235_932 ();
 FILLER_ASAP7_75t_R FILLER_235_948 ();
 FILLER_ASAP7_75t_R FILLER_235_964 ();
 FILLER_ASAP7_75t_R FILLER_235_969 ();
 DECAPx6_ASAP7_75t_R FILLER_235_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_999 ();
 DECAPx2_ASAP7_75t_R FILLER_235_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1009 ();
 DECAPx4_ASAP7_75t_R FILLER_235_1013 ();
 DECAPx6_ASAP7_75t_R FILLER_235_1026 ();
 FILLER_ASAP7_75t_R FILLER_235_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_235_1048 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_1068 ();
 FILLER_ASAP7_75t_R FILLER_235_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_235_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_236_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_16 ();
 DECAPx4_ASAP7_75t_R FILLER_236_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_32 ();
 DECAPx1_ASAP7_75t_R FILLER_236_39 ();
 DECAPx1_ASAP7_75t_R FILLER_236_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_50 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_57 ();
 DECAPx2_ASAP7_75t_R FILLER_236_66 ();
 FILLER_ASAP7_75t_R FILLER_236_81 ();
 FILLER_ASAP7_75t_R FILLER_236_109 ();
 FILLER_ASAP7_75t_R FILLER_236_137 ();
 FILLER_ASAP7_75t_R FILLER_236_142 ();
 FILLER_ASAP7_75t_R FILLER_236_147 ();
 DECAPx1_ASAP7_75t_R FILLER_236_155 ();
 DECAPx6_ASAP7_75t_R FILLER_236_165 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_179 ();
 FILLER_ASAP7_75t_R FILLER_236_208 ();
 DECAPx6_ASAP7_75t_R FILLER_236_216 ();
 DECAPx2_ASAP7_75t_R FILLER_236_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_236 ();
 DECAPx4_ASAP7_75t_R FILLER_236_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_250 ();
 FILLER_ASAP7_75t_R FILLER_236_259 ();
 FILLER_ASAP7_75t_R FILLER_236_267 ();
 DECAPx2_ASAP7_75t_R FILLER_236_295 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_301 ();
 DECAPx4_ASAP7_75t_R FILLER_236_307 ();
 FILLER_ASAP7_75t_R FILLER_236_325 ();
 DECAPx1_ASAP7_75t_R FILLER_236_333 ();
 DECAPx1_ASAP7_75t_R FILLER_236_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_347 ();
 DECAPx1_ASAP7_75t_R FILLER_236_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_355 ();
 FILLER_ASAP7_75t_R FILLER_236_382 ();
 DECAPx2_ASAP7_75t_R FILLER_236_390 ();
 DECAPx1_ASAP7_75t_R FILLER_236_422 ();
 FILLER_ASAP7_75t_R FILLER_236_432 ();
 FILLER_ASAP7_75t_R FILLER_236_460 ();
 FILLER_ASAP7_75t_R FILLER_236_464 ();
 FILLER_ASAP7_75t_R FILLER_236_469 ();
 FILLER_ASAP7_75t_R FILLER_236_477 ();
 DECAPx2_ASAP7_75t_R FILLER_236_487 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_493 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_502 ();
 DECAPx1_ASAP7_75t_R FILLER_236_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_515 ();
 DECAPx2_ASAP7_75t_R FILLER_236_519 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_525 ();
 DECAPx2_ASAP7_75t_R FILLER_236_534 ();
 DECAPx1_ASAP7_75t_R FILLER_236_543 ();
 DECAPx10_ASAP7_75t_R FILLER_236_553 ();
 DECAPx10_ASAP7_75t_R FILLER_236_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_597 ();
 DECAPx2_ASAP7_75t_R FILLER_236_604 ();
 FILLER_ASAP7_75t_R FILLER_236_610 ();
 DECAPx1_ASAP7_75t_R FILLER_236_618 ();
 FILLER_ASAP7_75t_R FILLER_236_630 ();
 DECAPx2_ASAP7_75t_R FILLER_236_635 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_641 ();
 FILLER_ASAP7_75t_R FILLER_236_650 ();
 DECAPx4_ASAP7_75t_R FILLER_236_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_668 ();
 DECAPx4_ASAP7_75t_R FILLER_236_683 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_707 ();
 DECAPx2_ASAP7_75t_R FILLER_236_713 ();
 DECAPx4_ASAP7_75t_R FILLER_236_722 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_732 ();
 FILLER_ASAP7_75t_R FILLER_236_738 ();
 DECAPx4_ASAP7_75t_R FILLER_236_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_756 ();
 FILLER_ASAP7_75t_R FILLER_236_763 ();
 DECAPx2_ASAP7_75t_R FILLER_236_779 ();
 FILLER_ASAP7_75t_R FILLER_236_785 ();
 DECAPx2_ASAP7_75t_R FILLER_236_790 ();
 DECAPx2_ASAP7_75t_R FILLER_236_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_805 ();
 DECAPx10_ASAP7_75t_R FILLER_236_809 ();
 DECAPx6_ASAP7_75t_R FILLER_236_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_851 ();
 FILLER_ASAP7_75t_R FILLER_236_855 ();
 DECAPx4_ASAP7_75t_R FILLER_236_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_870 ();
 FILLER_ASAP7_75t_R FILLER_236_877 ();
 DECAPx1_ASAP7_75t_R FILLER_236_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_889 ();
 FILLER_ASAP7_75t_R FILLER_236_893 ();
 DECAPx10_ASAP7_75t_R FILLER_236_901 ();
 DECAPx10_ASAP7_75t_R FILLER_236_923 ();
 DECAPx6_ASAP7_75t_R FILLER_236_945 ();
 DECAPx2_ASAP7_75t_R FILLER_236_959 ();
 DECAPx10_ASAP7_75t_R FILLER_236_968 ();
 DECAPx10_ASAP7_75t_R FILLER_236_990 ();
 FILLER_ASAP7_75t_R FILLER_236_1026 ();
 FILLER_ASAP7_75t_R FILLER_236_1042 ();
 FILLER_ASAP7_75t_R FILLER_236_1058 ();
 DECAPx4_ASAP7_75t_R FILLER_236_1063 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_236_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_237_2 ();
 DECAPx2_ASAP7_75t_R FILLER_237_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_22 ();
 DECAPx10_ASAP7_75t_R FILLER_237_29 ();
 DECAPx1_ASAP7_75t_R FILLER_237_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_55 ();
 DECAPx10_ASAP7_75t_R FILLER_237_64 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_237_86 ();
 DECAPx1_ASAP7_75t_R FILLER_237_95 ();
 DECAPx4_ASAP7_75t_R FILLER_237_102 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_237_112 ();
 DECAPx1_ASAP7_75t_R FILLER_237_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_125 ();
 DECAPx6_ASAP7_75t_R FILLER_237_129 ();
 DECAPx2_ASAP7_75t_R FILLER_237_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_149 ();
 DECAPx4_ASAP7_75t_R FILLER_237_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_168 ();
 DECAPx4_ASAP7_75t_R FILLER_237_177 ();
 FILLER_ASAP7_75t_R FILLER_237_187 ();
 DECAPx2_ASAP7_75t_R FILLER_237_195 ();
 FILLER_ASAP7_75t_R FILLER_237_207 ();
 DECAPx2_ASAP7_75t_R FILLER_237_217 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_237_223 ();
 DECAPx6_ASAP7_75t_R FILLER_237_232 ();
 DECAPx1_ASAP7_75t_R FILLER_237_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_250 ();
 FILLER_ASAP7_75t_R FILLER_237_257 ();
 DECAPx6_ASAP7_75t_R FILLER_237_270 ();
 DECAPx1_ASAP7_75t_R FILLER_237_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_288 ();
 DECAPx2_ASAP7_75t_R FILLER_237_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_301 ();
 DECAPx6_ASAP7_75t_R FILLER_237_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_322 ();
 FILLER_ASAP7_75t_R FILLER_237_331 ();
 DECAPx4_ASAP7_75t_R FILLER_237_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_369 ();
 DECAPx6_ASAP7_75t_R FILLER_237_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_387 ();
 DECAPx1_ASAP7_75t_R FILLER_237_394 ();
 DECAPx2_ASAP7_75t_R FILLER_237_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_410 ();
 DECAPx2_ASAP7_75t_R FILLER_237_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_420 ();
 DECAPx1_ASAP7_75t_R FILLER_237_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_428 ();
 FILLER_ASAP7_75t_R FILLER_237_437 ();
 DECAPx2_ASAP7_75t_R FILLER_237_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_451 ();
 FILLER_ASAP7_75t_R FILLER_237_478 ();
 FILLER_ASAP7_75t_R FILLER_237_486 ();
 DECAPx6_ASAP7_75t_R FILLER_237_494 ();
 DECAPx2_ASAP7_75t_R FILLER_237_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_514 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_237_541 ();
 DECAPx2_ASAP7_75t_R FILLER_237_552 ();
 FILLER_ASAP7_75t_R FILLER_237_558 ();
 FILLER_ASAP7_75t_R FILLER_237_586 ();
 DECAPx1_ASAP7_75t_R FILLER_237_594 ();
 DECAPx10_ASAP7_75t_R FILLER_237_606 ();
 DECAPx4_ASAP7_75t_R FILLER_237_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_638 ();
 FILLER_ASAP7_75t_R FILLER_237_653 ();
 FILLER_ASAP7_75t_R FILLER_237_661 ();
 FILLER_ASAP7_75t_R FILLER_237_666 ();
 DECAPx6_ASAP7_75t_R FILLER_237_671 ();
 DECAPx2_ASAP7_75t_R FILLER_237_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_691 ();
 FILLER_ASAP7_75t_R FILLER_237_706 ();
 DECAPx10_ASAP7_75t_R FILLER_237_711 ();
 DECAPx10_ASAP7_75t_R FILLER_237_733 ();
 DECAPx4_ASAP7_75t_R FILLER_237_755 ();
 FILLER_ASAP7_75t_R FILLER_237_765 ();
 FILLER_ASAP7_75t_R FILLER_237_773 ();
 DECAPx6_ASAP7_75t_R FILLER_237_778 ();
 DECAPx2_ASAP7_75t_R FILLER_237_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_798 ();
 DECAPx2_ASAP7_75t_R FILLER_237_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_819 ();
 FILLER_ASAP7_75t_R FILLER_237_834 ();
 FILLER_ASAP7_75t_R FILLER_237_839 ();
 FILLER_ASAP7_75t_R FILLER_237_844 ();
 DECAPx1_ASAP7_75t_R FILLER_237_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_853 ();
 FILLER_ASAP7_75t_R FILLER_237_868 ();
 DECAPx10_ASAP7_75t_R FILLER_237_884 ();
 DECAPx4_ASAP7_75t_R FILLER_237_906 ();
 DECAPx2_ASAP7_75t_R FILLER_237_919 ();
 FILLER_ASAP7_75t_R FILLER_237_927 ();
 DECAPx4_ASAP7_75t_R FILLER_237_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_942 ();
 DECAPx2_ASAP7_75t_R FILLER_237_946 ();
 FILLER_ASAP7_75t_R FILLER_237_952 ();
 DECAPx6_ASAP7_75t_R FILLER_237_957 ();
 FILLER_ASAP7_75t_R FILLER_237_971 ();
 FILLER_ASAP7_75t_R FILLER_237_987 ();
 DECAPx2_ASAP7_75t_R FILLER_237_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_998 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_237_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_237_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_1023 ();
 DECAPx4_ASAP7_75t_R FILLER_237_1027 ();
 FILLER_ASAP7_75t_R FILLER_237_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_237_1353 ();
 FILLER_ASAP7_75t_R FILLER_237_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_238_2 ();
 DECAPx1_ASAP7_75t_R FILLER_238_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_20 ();
 FILLER_ASAP7_75t_R FILLER_238_47 ();
 FILLER_ASAP7_75t_R FILLER_238_55 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_65 ();
 DECAPx6_ASAP7_75t_R FILLER_238_74 ();
 FILLER_ASAP7_75t_R FILLER_238_94 ();
 DECAPx1_ASAP7_75t_R FILLER_238_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_110 ();
 DECAPx4_ASAP7_75t_R FILLER_238_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_127 ();
 DECAPx2_ASAP7_75t_R FILLER_238_134 ();
 FILLER_ASAP7_75t_R FILLER_238_140 ();
 DECAPx2_ASAP7_75t_R FILLER_238_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_154 ();
 DECAPx2_ASAP7_75t_R FILLER_238_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_167 ();
 FILLER_ASAP7_75t_R FILLER_238_176 ();
 DECAPx4_ASAP7_75t_R FILLER_238_184 ();
 FILLER_ASAP7_75t_R FILLER_238_194 ();
 DECAPx4_ASAP7_75t_R FILLER_238_199 ();
 FILLER_ASAP7_75t_R FILLER_238_217 ();
 FILLER_ASAP7_75t_R FILLER_238_225 ();
 FILLER_ASAP7_75t_R FILLER_238_235 ();
 DECAPx1_ASAP7_75t_R FILLER_238_243 ();
 DECAPx10_ASAP7_75t_R FILLER_238_255 ();
 DECAPx2_ASAP7_75t_R FILLER_238_277 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_283 ();
 DECAPx4_ASAP7_75t_R FILLER_238_312 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_322 ();
 DECAPx1_ASAP7_75t_R FILLER_238_331 ();
 DECAPx4_ASAP7_75t_R FILLER_238_341 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_351 ();
 DECAPx2_ASAP7_75t_R FILLER_238_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_366 ();
 DECAPx1_ASAP7_75t_R FILLER_238_370 ();
 DECAPx2_ASAP7_75t_R FILLER_238_377 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_383 ();
 DECAPx4_ASAP7_75t_R FILLER_238_412 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_422 ();
 DECAPx6_ASAP7_75t_R FILLER_238_433 ();
 DECAPx2_ASAP7_75t_R FILLER_238_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_453 ();
 FILLER_ASAP7_75t_R FILLER_238_460 ();
 FILLER_ASAP7_75t_R FILLER_238_464 ();
 FILLER_ASAP7_75t_R FILLER_238_472 ();
 DECAPx10_ASAP7_75t_R FILLER_238_477 ();
 DECAPx2_ASAP7_75t_R FILLER_238_499 ();
 DECAPx4_ASAP7_75t_R FILLER_238_511 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_527 ();
 DECAPx4_ASAP7_75t_R FILLER_238_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_543 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_550 ();
 FILLER_ASAP7_75t_R FILLER_238_561 ();
 DECAPx2_ASAP7_75t_R FILLER_238_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_575 ();
 DECAPx1_ASAP7_75t_R FILLER_238_602 ();
 FILLER_ASAP7_75t_R FILLER_238_614 ();
 FILLER_ASAP7_75t_R FILLER_238_622 ();
 DECAPx6_ASAP7_75t_R FILLER_238_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_644 ();
 FILLER_ASAP7_75t_R FILLER_238_648 ();
 DECAPx4_ASAP7_75t_R FILLER_238_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_674 ();
 DECAPx6_ASAP7_75t_R FILLER_238_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_695 ();
 DECAPx6_ASAP7_75t_R FILLER_238_699 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_713 ();
 DECAPx2_ASAP7_75t_R FILLER_238_719 ();
 FILLER_ASAP7_75t_R FILLER_238_725 ();
 DECAPx10_ASAP7_75t_R FILLER_238_733 ();
 DECAPx10_ASAP7_75t_R FILLER_238_755 ();
 FILLER_ASAP7_75t_R FILLER_238_786 ();
 DECAPx10_ASAP7_75t_R FILLER_238_791 ();
 DECAPx4_ASAP7_75t_R FILLER_238_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_823 ();
 FILLER_ASAP7_75t_R FILLER_238_830 ();
 DECAPx10_ASAP7_75t_R FILLER_238_835 ();
 DECAPx6_ASAP7_75t_R FILLER_238_857 ();
 FILLER_ASAP7_75t_R FILLER_238_871 ();
 DECAPx2_ASAP7_75t_R FILLER_238_879 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_885 ();
 FILLER_ASAP7_75t_R FILLER_238_902 ();
 DECAPx2_ASAP7_75t_R FILLER_238_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_916 ();
 DECAPx2_ASAP7_75t_R FILLER_238_923 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_929 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_938 ();
 DECAPx2_ASAP7_75t_R FILLER_238_947 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_959 ();
 FILLER_ASAP7_75t_R FILLER_238_968 ();
 DECAPx2_ASAP7_75t_R FILLER_238_976 ();
 FILLER_ASAP7_75t_R FILLER_238_985 ();
 DECAPx4_ASAP7_75t_R FILLER_238_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1003 ();
 DECAPx4_ASAP7_75t_R FILLER_238_1018 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_1028 ();
 DECAPx6_ASAP7_75t_R FILLER_238_1034 ();
 FILLER_ASAP7_75t_R FILLER_238_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_238_1053 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1142 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_238_1340 ();
 DECAPx6_ASAP7_75t_R FILLER_238_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_239_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_24 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_33 ();
 DECAPx2_ASAP7_75t_R FILLER_239_39 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_45 ();
 FILLER_ASAP7_75t_R FILLER_239_51 ();
 DECAPx4_ASAP7_75t_R FILLER_239_59 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_69 ();
 FILLER_ASAP7_75t_R FILLER_239_80 ();
 DECAPx2_ASAP7_75t_R FILLER_239_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_96 ();
 DECAPx2_ASAP7_75t_R FILLER_239_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_131 ();
 DECAPx2_ASAP7_75t_R FILLER_239_140 ();
 FILLER_ASAP7_75t_R FILLER_239_146 ();
 FILLER_ASAP7_75t_R FILLER_239_154 ();
 DECAPx2_ASAP7_75t_R FILLER_239_162 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_168 ();
 DECAPx10_ASAP7_75t_R FILLER_239_177 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_199 ();
 DECAPx4_ASAP7_75t_R FILLER_239_208 ();
 FILLER_ASAP7_75t_R FILLER_239_218 ();
 DECAPx1_ASAP7_75t_R FILLER_239_223 ();
 FILLER_ASAP7_75t_R FILLER_239_235 ();
 DECAPx1_ASAP7_75t_R FILLER_239_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_247 ();
 DECAPx2_ASAP7_75t_R FILLER_239_254 ();
 FILLER_ASAP7_75t_R FILLER_239_286 ();
 DECAPx2_ASAP7_75t_R FILLER_239_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_300 ();
 DECAPx1_ASAP7_75t_R FILLER_239_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_308 ();
 FILLER_ASAP7_75t_R FILLER_239_312 ();
 DECAPx2_ASAP7_75t_R FILLER_239_322 ();
 DECAPx6_ASAP7_75t_R FILLER_239_334 ();
 DECAPx1_ASAP7_75t_R FILLER_239_348 ();
 FILLER_ASAP7_75t_R FILLER_239_378 ();
 DECAPx2_ASAP7_75t_R FILLER_239_386 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_398 ();
 DECAPx2_ASAP7_75t_R FILLER_239_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_410 ();
 FILLER_ASAP7_75t_R FILLER_239_414 ();
 FILLER_ASAP7_75t_R FILLER_239_424 ();
 DECAPx1_ASAP7_75t_R FILLER_239_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_436 ();
 DECAPx6_ASAP7_75t_R FILLER_239_443 ();
 DECAPx2_ASAP7_75t_R FILLER_239_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_463 ();
 DECAPx6_ASAP7_75t_R FILLER_239_470 ();
 DECAPx1_ASAP7_75t_R FILLER_239_484 ();
 DECAPx1_ASAP7_75t_R FILLER_239_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_500 ();
 DECAPx10_ASAP7_75t_R FILLER_239_527 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_549 ();
 DECAPx1_ASAP7_75t_R FILLER_239_558 ();
 DECAPx2_ASAP7_75t_R FILLER_239_568 ();
 DECAPx1_ASAP7_75t_R FILLER_239_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_581 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_588 ();
 DECAPx2_ASAP7_75t_R FILLER_239_594 ();
 FILLER_ASAP7_75t_R FILLER_239_600 ();
 DECAPx6_ASAP7_75t_R FILLER_239_608 ();
 FILLER_ASAP7_75t_R FILLER_239_622 ();
 DECAPx10_ASAP7_75t_R FILLER_239_630 ();
 DECAPx4_ASAP7_75t_R FILLER_239_652 ();
 FILLER_ASAP7_75t_R FILLER_239_662 ();
 FILLER_ASAP7_75t_R FILLER_239_670 ();
 DECAPx2_ASAP7_75t_R FILLER_239_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_692 ();
 FILLER_ASAP7_75t_R FILLER_239_707 ();
 FILLER_ASAP7_75t_R FILLER_239_712 ();
 FILLER_ASAP7_75t_R FILLER_239_723 ();
 FILLER_ASAP7_75t_R FILLER_239_731 ();
 FILLER_ASAP7_75t_R FILLER_239_739 ();
 FILLER_ASAP7_75t_R FILLER_239_747 ();
 FILLER_ASAP7_75t_R FILLER_239_755 ();
 DECAPx6_ASAP7_75t_R FILLER_239_763 ();
 FILLER_ASAP7_75t_R FILLER_239_777 ();
 FILLER_ASAP7_75t_R FILLER_239_782 ();
 DECAPx2_ASAP7_75t_R FILLER_239_787 ();
 FILLER_ASAP7_75t_R FILLER_239_793 ();
 DECAPx1_ASAP7_75t_R FILLER_239_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_805 ();
 DECAPx10_ASAP7_75t_R FILLER_239_818 ();
 DECAPx10_ASAP7_75t_R FILLER_239_854 ();
 DECAPx2_ASAP7_75t_R FILLER_239_876 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_882 ();
 DECAPx2_ASAP7_75t_R FILLER_239_888 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_894 ();
 DECAPx2_ASAP7_75t_R FILLER_239_900 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_906 ();
 FILLER_ASAP7_75t_R FILLER_239_923 ();
 DECAPx2_ASAP7_75t_R FILLER_239_927 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_933 ();
 DECAPx2_ASAP7_75t_R FILLER_239_950 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_956 ();
 DECAPx4_ASAP7_75t_R FILLER_239_973 ();
 FILLER_ASAP7_75t_R FILLER_239_983 ();
 FILLER_ASAP7_75t_R FILLER_239_999 ();
 DECAPx4_ASAP7_75t_R FILLER_239_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_239_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_1046 ();
 FILLER_ASAP7_75t_R FILLER_239_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1176 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1220 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1264 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1286 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1308 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_239_1352 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_1374 ();
 DECAPx10_ASAP7_75t_R FILLER_240_2 ();
 FILLER_ASAP7_75t_R FILLER_240_24 ();
 DECAPx10_ASAP7_75t_R FILLER_240_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_74 ();
 FILLER_ASAP7_75t_R FILLER_240_81 ();
 DECAPx6_ASAP7_75t_R FILLER_240_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_103 ();
 DECAPx1_ASAP7_75t_R FILLER_240_110 ();
 DECAPx2_ASAP7_75t_R FILLER_240_117 ();
 FILLER_ASAP7_75t_R FILLER_240_129 ();
 DECAPx1_ASAP7_75t_R FILLER_240_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_143 ();
 DECAPx10_ASAP7_75t_R FILLER_240_150 ();
 DECAPx2_ASAP7_75t_R FILLER_240_172 ();
 DECAPx2_ASAP7_75t_R FILLER_240_184 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_240_190 ();
 DECAPx10_ASAP7_75t_R FILLER_240_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_241 ();
 FILLER_ASAP7_75t_R FILLER_240_248 ();
 FILLER_ASAP7_75t_R FILLER_240_288 ();
 FILLER_ASAP7_75t_R FILLER_240_293 ();
 DECAPx4_ASAP7_75t_R FILLER_240_301 ();
 FILLER_ASAP7_75t_R FILLER_240_311 ();
 DECAPx2_ASAP7_75t_R FILLER_240_319 ();
 FILLER_ASAP7_75t_R FILLER_240_325 ();
 FILLER_ASAP7_75t_R FILLER_240_335 ();
 DECAPx2_ASAP7_75t_R FILLER_240_343 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_240_349 ();
 DECAPx10_ASAP7_75t_R FILLER_240_358 ();
 DECAPx2_ASAP7_75t_R FILLER_240_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_386 ();
 FILLER_ASAP7_75t_R FILLER_240_396 ();
 DECAPx1_ASAP7_75t_R FILLER_240_404 ();
 FILLER_ASAP7_75t_R FILLER_240_414 ();
 DECAPx1_ASAP7_75t_R FILLER_240_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_428 ();
 FILLER_ASAP7_75t_R FILLER_240_435 ();
 FILLER_ASAP7_75t_R FILLER_240_443 ();
 DECAPx2_ASAP7_75t_R FILLER_240_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_240_459 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_240_464 ();
 FILLER_ASAP7_75t_R FILLER_240_476 ();
 FILLER_ASAP7_75t_R FILLER_240_481 ();
 FILLER_ASAP7_75t_R FILLER_240_489 ();
 DECAPx2_ASAP7_75t_R FILLER_240_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_503 ();
 DECAPx2_ASAP7_75t_R FILLER_240_510 ();
 DECAPx2_ASAP7_75t_R FILLER_240_519 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_240_525 ();
 DECAPx4_ASAP7_75t_R FILLER_240_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_544 ();
 DECAPx10_ASAP7_75t_R FILLER_240_551 ();
 DECAPx6_ASAP7_75t_R FILLER_240_573 ();
 DECAPx2_ASAP7_75t_R FILLER_240_587 ();
 FILLER_ASAP7_75t_R FILLER_240_599 ();
 DECAPx4_ASAP7_75t_R FILLER_240_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_614 ();
 DECAPx1_ASAP7_75t_R FILLER_240_621 ();
 FILLER_ASAP7_75t_R FILLER_240_631 ();
 DECAPx6_ASAP7_75t_R FILLER_240_636 ();
 FILLER_ASAP7_75t_R FILLER_240_650 ();
 DECAPx6_ASAP7_75t_R FILLER_240_655 ();
 DECAPx2_ASAP7_75t_R FILLER_240_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_675 ();
 DECAPx10_ASAP7_75t_R FILLER_240_682 ();
 DECAPx2_ASAP7_75t_R FILLER_240_704 ();
 FILLER_ASAP7_75t_R FILLER_240_710 ();
 DECAPx2_ASAP7_75t_R FILLER_240_721 ();
 FILLER_ASAP7_75t_R FILLER_240_741 ();
 DECAPx1_ASAP7_75t_R FILLER_240_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_753 ();
 DECAPx10_ASAP7_75t_R FILLER_240_769 ();
 FILLER_ASAP7_75t_R FILLER_240_791 ();
 FILLER_ASAP7_75t_R FILLER_240_807 ();
 DECAPx4_ASAP7_75t_R FILLER_240_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_825 ();
 DECAPx2_ASAP7_75t_R FILLER_240_832 ();
 FILLER_ASAP7_75t_R FILLER_240_838 ();
 DECAPx4_ASAP7_75t_R FILLER_240_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_853 ();
 FILLER_ASAP7_75t_R FILLER_240_860 ();
 FILLER_ASAP7_75t_R FILLER_240_868 ();
 DECAPx2_ASAP7_75t_R FILLER_240_873 ();
 DECAPx6_ASAP7_75t_R FILLER_240_882 ();
 DECAPx4_ASAP7_75t_R FILLER_240_910 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_240_923 ();
 DECAPx6_ASAP7_75t_R FILLER_240_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_943 ();
 FILLER_ASAP7_75t_R FILLER_240_947 ();
 DECAPx6_ASAP7_75t_R FILLER_240_952 ();
 FILLER_ASAP7_75t_R FILLER_240_966 ();
 DECAPx4_ASAP7_75t_R FILLER_240_971 ();
 FILLER_ASAP7_75t_R FILLER_240_981 ();
 DECAPx6_ASAP7_75t_R FILLER_240_986 ();
 DECAPx2_ASAP7_75t_R FILLER_240_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_240_1010 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_240_1020 ();
 FILLER_ASAP7_75t_R FILLER_240_1029 ();
 FILLER_ASAP7_75t_R FILLER_240_1037 ();
 FILLER_ASAP7_75t_R FILLER_240_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1072 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_240_1336 ();
 DECAPx6_ASAP7_75t_R FILLER_240_1358 ();
 DECAPx1_ASAP7_75t_R FILLER_240_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_241_2 ();
 FILLER_ASAP7_75t_R FILLER_241_24 ();
 FILLER_ASAP7_75t_R FILLER_241_32 ();
 FILLER_ASAP7_75t_R FILLER_241_40 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_45 ();
 DECAPx2_ASAP7_75t_R FILLER_241_74 ();
 FILLER_ASAP7_75t_R FILLER_241_86 ();
 DECAPx6_ASAP7_75t_R FILLER_241_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_105 ();
 DECAPx4_ASAP7_75t_R FILLER_241_112 ();
 FILLER_ASAP7_75t_R FILLER_241_122 ();
 DECAPx4_ASAP7_75t_R FILLER_241_127 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_137 ();
 DECAPx4_ASAP7_75t_R FILLER_241_148 ();
 DECAPx2_ASAP7_75t_R FILLER_241_164 ();
 FILLER_ASAP7_75t_R FILLER_241_196 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_204 ();
 DECAPx10_ASAP7_75t_R FILLER_241_210 ();
 DECAPx10_ASAP7_75t_R FILLER_241_232 ();
 DECAPx1_ASAP7_75t_R FILLER_241_254 ();
 FILLER_ASAP7_75t_R FILLER_241_264 ();
 DECAPx2_ASAP7_75t_R FILLER_241_272 ();
 FILLER_ASAP7_75t_R FILLER_241_284 ();
 DECAPx6_ASAP7_75t_R FILLER_241_294 ();
 DECAPx1_ASAP7_75t_R FILLER_241_308 ();
 DECAPx1_ASAP7_75t_R FILLER_241_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_322 ();
 DECAPx2_ASAP7_75t_R FILLER_241_326 ();
 FILLER_ASAP7_75t_R FILLER_241_332 ();
 DECAPx2_ASAP7_75t_R FILLER_241_340 ();
 DECAPx6_ASAP7_75t_R FILLER_241_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_386 ();
 FILLER_ASAP7_75t_R FILLER_241_413 ();
 DECAPx10_ASAP7_75t_R FILLER_241_421 ();
 FILLER_ASAP7_75t_R FILLER_241_443 ();
 FILLER_ASAP7_75t_R FILLER_241_454 ();
 DECAPx2_ASAP7_75t_R FILLER_241_482 ();
 FILLER_ASAP7_75t_R FILLER_241_496 ();
 DECAPx6_ASAP7_75t_R FILLER_241_504 ();
 FILLER_ASAP7_75t_R FILLER_241_544 ();
 DECAPx1_ASAP7_75t_R FILLER_241_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_558 ();
 FILLER_ASAP7_75t_R FILLER_241_567 ();
 DECAPx2_ASAP7_75t_R FILLER_241_575 ();
 FILLER_ASAP7_75t_R FILLER_241_581 ();
 FILLER_ASAP7_75t_R FILLER_241_609 ();
 DECAPx4_ASAP7_75t_R FILLER_241_637 ();
 FILLER_ASAP7_75t_R FILLER_241_653 ();
 DECAPx2_ASAP7_75t_R FILLER_241_661 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_667 ();
 DECAPx6_ASAP7_75t_R FILLER_241_676 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_690 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_696 ();
 DECAPx4_ASAP7_75t_R FILLER_241_702 ();
 FILLER_ASAP7_75t_R FILLER_241_712 ();
 DECAPx10_ASAP7_75t_R FILLER_241_717 ();
 DECAPx1_ASAP7_75t_R FILLER_241_739 ();
 FILLER_ASAP7_75t_R FILLER_241_749 ();
 FILLER_ASAP7_75t_R FILLER_241_758 ();
 FILLER_ASAP7_75t_R FILLER_241_774 ();
 DECAPx2_ASAP7_75t_R FILLER_241_788 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_794 ();
 FILLER_ASAP7_75t_R FILLER_241_806 ();
 DECAPx2_ASAP7_75t_R FILLER_241_814 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_820 ();
 DECAPx2_ASAP7_75t_R FILLER_241_837 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_843 ();
 FILLER_ASAP7_75t_R FILLER_241_849 ();
 DECAPx2_ASAP7_75t_R FILLER_241_865 ();
 DECAPx4_ASAP7_75t_R FILLER_241_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_895 ();
 DECAPx2_ASAP7_75t_R FILLER_241_899 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_905 ();
 DECAPx6_ASAP7_75t_R FILLER_241_911 ();
 DECAPx10_ASAP7_75t_R FILLER_241_927 ();
 DECAPx10_ASAP7_75t_R FILLER_241_949 ();
 DECAPx6_ASAP7_75t_R FILLER_241_971 ();
 DECAPx2_ASAP7_75t_R FILLER_241_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_991 ();
 DECAPx1_ASAP7_75t_R FILLER_241_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_999 ();
 DECAPx4_ASAP7_75t_R FILLER_241_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_241_1038 ();
 FILLER_ASAP7_75t_R FILLER_241_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_241_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_241_1361 ();
 FILLER_ASAP7_75t_R FILLER_241_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_242_2 ();
 DECAPx10_ASAP7_75t_R FILLER_242_24 ();
 DECAPx4_ASAP7_75t_R FILLER_242_46 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_56 ();
 DECAPx1_ASAP7_75t_R FILLER_242_65 ();
 FILLER_ASAP7_75t_R FILLER_242_95 ();
 DECAPx6_ASAP7_75t_R FILLER_242_123 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_137 ();
 DECAPx4_ASAP7_75t_R FILLER_242_148 ();
 FILLER_ASAP7_75t_R FILLER_242_158 ();
 FILLER_ASAP7_75t_R FILLER_242_163 ();
 DECAPx1_ASAP7_75t_R FILLER_242_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_175 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_182 ();
 DECAPx6_ASAP7_75t_R FILLER_242_188 ();
 FILLER_ASAP7_75t_R FILLER_242_202 ();
 DECAPx6_ASAP7_75t_R FILLER_242_210 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_232 ();
 FILLER_ASAP7_75t_R FILLER_242_241 ();
 DECAPx6_ASAP7_75t_R FILLER_242_249 ();
 FILLER_ASAP7_75t_R FILLER_242_263 ();
 DECAPx6_ASAP7_75t_R FILLER_242_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_285 ();
 FILLER_ASAP7_75t_R FILLER_242_294 ();
 DECAPx2_ASAP7_75t_R FILLER_242_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_308 ();
 DECAPx4_ASAP7_75t_R FILLER_242_335 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_345 ();
 DECAPx2_ASAP7_75t_R FILLER_242_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_360 ();
 DECAPx1_ASAP7_75t_R FILLER_242_364 ();
 DECAPx6_ASAP7_75t_R FILLER_242_374 ();
 DECAPx2_ASAP7_75t_R FILLER_242_388 ();
 FILLER_ASAP7_75t_R FILLER_242_400 ();
 DECAPx10_ASAP7_75t_R FILLER_242_405 ();
 DECAPx2_ASAP7_75t_R FILLER_242_427 ();
 FILLER_ASAP7_75t_R FILLER_242_433 ();
 DECAPx6_ASAP7_75t_R FILLER_242_443 ();
 DECAPx1_ASAP7_75t_R FILLER_242_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_461 ();
 DECAPx1_ASAP7_75t_R FILLER_242_464 ();
 FILLER_ASAP7_75t_R FILLER_242_471 ();
 DECAPx10_ASAP7_75t_R FILLER_242_479 ();
 DECAPx1_ASAP7_75t_R FILLER_242_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_505 ();
 DECAPx4_ASAP7_75t_R FILLER_242_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_522 ();
 DECAPx1_ASAP7_75t_R FILLER_242_529 ();
 DECAPx2_ASAP7_75t_R FILLER_242_536 ();
 DECAPx4_ASAP7_75t_R FILLER_242_545 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_555 ();
 FILLER_ASAP7_75t_R FILLER_242_564 ();
 FILLER_ASAP7_75t_R FILLER_242_572 ();
 DECAPx1_ASAP7_75t_R FILLER_242_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_587 ();
 DECAPx1_ASAP7_75t_R FILLER_242_594 ();
 DECAPx10_ASAP7_75t_R FILLER_242_601 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_623 ();
 DECAPx6_ASAP7_75t_R FILLER_242_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_643 ();
 DECAPx4_ASAP7_75t_R FILLER_242_658 ();
 FILLER_ASAP7_75t_R FILLER_242_682 ();
 DECAPx4_ASAP7_75t_R FILLER_242_693 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_703 ();
 DECAPx6_ASAP7_75t_R FILLER_242_720 ();
 DECAPx6_ASAP7_75t_R FILLER_242_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_757 ();
 DECAPx4_ASAP7_75t_R FILLER_242_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_777 ();
 DECAPx4_ASAP7_75t_R FILLER_242_787 ();
 FILLER_ASAP7_75t_R FILLER_242_797 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_805 ();
 DECAPx4_ASAP7_75t_R FILLER_242_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_824 ();
 DECAPx6_ASAP7_75t_R FILLER_242_839 ();
 FILLER_ASAP7_75t_R FILLER_242_853 ();
 DECAPx4_ASAP7_75t_R FILLER_242_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_871 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_875 ();
 FILLER_ASAP7_75t_R FILLER_242_881 ();
 DECAPx2_ASAP7_75t_R FILLER_242_886 ();
 FILLER_ASAP7_75t_R FILLER_242_892 ();
 DECAPx1_ASAP7_75t_R FILLER_242_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_901 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_905 ();
 DECAPx6_ASAP7_75t_R FILLER_242_922 ();
 DECAPx1_ASAP7_75t_R FILLER_242_936 ();
 FILLER_ASAP7_75t_R FILLER_242_954 ();
 FILLER_ASAP7_75t_R FILLER_242_959 ();
 FILLER_ASAP7_75t_R FILLER_242_964 ();
 FILLER_ASAP7_75t_R FILLER_242_969 ();
 DECAPx1_ASAP7_75t_R FILLER_242_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_978 ();
 FILLER_ASAP7_75t_R FILLER_242_993 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_1009 ();
 FILLER_ASAP7_75t_R FILLER_242_1018 ();
 FILLER_ASAP7_75t_R FILLER_242_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_242_1031 ();
 FILLER_ASAP7_75t_R FILLER_242_1037 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_242_1348 ();
 DECAPx2_ASAP7_75t_R FILLER_242_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_243_2 ();
 DECAPx2_ASAP7_75t_R FILLER_243_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_30 ();
 FILLER_ASAP7_75t_R FILLER_243_37 ();
 DECAPx4_ASAP7_75t_R FILLER_243_42 ();
 DECAPx1_ASAP7_75t_R FILLER_243_58 ();
 DECAPx4_ASAP7_75t_R FILLER_243_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_75 ();
 DECAPx1_ASAP7_75t_R FILLER_243_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_86 ();
 DECAPx4_ASAP7_75t_R FILLER_243_90 ();
 FILLER_ASAP7_75t_R FILLER_243_100 ();
 FILLER_ASAP7_75t_R FILLER_243_108 ();
 FILLER_ASAP7_75t_R FILLER_243_113 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_121 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_130 ();
 DECAPx2_ASAP7_75t_R FILLER_243_136 ();
 FILLER_ASAP7_75t_R FILLER_243_148 ();
 DECAPx1_ASAP7_75t_R FILLER_243_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_160 ();
 DECAPx2_ASAP7_75t_R FILLER_243_187 ();
 FILLER_ASAP7_75t_R FILLER_243_193 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_221 ();
 DECAPx2_ASAP7_75t_R FILLER_243_232 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_238 ();
 DECAPx2_ASAP7_75t_R FILLER_243_249 ();
 FILLER_ASAP7_75t_R FILLER_243_255 ();
 FILLER_ASAP7_75t_R FILLER_243_283 ();
 DECAPx6_ASAP7_75t_R FILLER_243_288 ();
 DECAPx2_ASAP7_75t_R FILLER_243_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_308 ();
 DECAPx10_ASAP7_75t_R FILLER_243_315 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_337 ();
 FILLER_ASAP7_75t_R FILLER_243_346 ();
 DECAPx2_ASAP7_75t_R FILLER_243_354 ();
 FILLER_ASAP7_75t_R FILLER_243_360 ();
 FILLER_ASAP7_75t_R FILLER_243_368 ();
 DECAPx10_ASAP7_75t_R FILLER_243_378 ();
 DECAPx6_ASAP7_75t_R FILLER_243_400 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_414 ();
 DECAPx1_ASAP7_75t_R FILLER_243_423 ();
 FILLER_ASAP7_75t_R FILLER_243_433 ();
 DECAPx4_ASAP7_75t_R FILLER_243_441 ();
 DECAPx2_ASAP7_75t_R FILLER_243_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_483 ();
 DECAPx2_ASAP7_75t_R FILLER_243_492 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_498 ();
 DECAPx10_ASAP7_75t_R FILLER_243_527 ();
 DECAPx10_ASAP7_75t_R FILLER_243_555 ();
 DECAPx4_ASAP7_75t_R FILLER_243_577 ();
 FILLER_ASAP7_75t_R FILLER_243_587 ();
 DECAPx6_ASAP7_75t_R FILLER_243_595 ();
 DECAPx10_ASAP7_75t_R FILLER_243_615 ();
 DECAPx2_ASAP7_75t_R FILLER_243_637 ();
 FILLER_ASAP7_75t_R FILLER_243_643 ();
 DECAPx2_ASAP7_75t_R FILLER_243_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_657 ();
 DECAPx2_ASAP7_75t_R FILLER_243_661 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_667 ();
 FILLER_ASAP7_75t_R FILLER_243_676 ();
 DECAPx4_ASAP7_75t_R FILLER_243_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_691 ();
 DECAPx1_ASAP7_75t_R FILLER_243_706 ();
 DECAPx2_ASAP7_75t_R FILLER_243_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_730 ();
 DECAPx10_ASAP7_75t_R FILLER_243_734 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_756 ();
 DECAPx10_ASAP7_75t_R FILLER_243_765 ();
 DECAPx6_ASAP7_75t_R FILLER_243_787 ();
 DECAPx2_ASAP7_75t_R FILLER_243_801 ();
 DECAPx2_ASAP7_75t_R FILLER_243_816 ();
 FILLER_ASAP7_75t_R FILLER_243_822 ();
 FILLER_ASAP7_75t_R FILLER_243_830 ();
 FILLER_ASAP7_75t_R FILLER_243_838 ();
 DECAPx10_ASAP7_75t_R FILLER_243_854 ();
 DECAPx2_ASAP7_75t_R FILLER_243_876 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_882 ();
 FILLER_ASAP7_75t_R FILLER_243_899 ();
 DECAPx1_ASAP7_75t_R FILLER_243_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_919 ();
 FILLER_ASAP7_75t_R FILLER_243_923 ();
 FILLER_ASAP7_75t_R FILLER_243_927 ();
 FILLER_ASAP7_75t_R FILLER_243_932 ();
 FILLER_ASAP7_75t_R FILLER_243_948 ();
 DECAPx1_ASAP7_75t_R FILLER_243_953 ();
 FILLER_ASAP7_75t_R FILLER_243_971 ();
 FILLER_ASAP7_75t_R FILLER_243_987 ();
 FILLER_ASAP7_75t_R FILLER_243_992 ();
 DECAPx4_ASAP7_75t_R FILLER_243_997 ();
 FILLER_ASAP7_75t_R FILLER_243_1007 ();
 DECAPx4_ASAP7_75t_R FILLER_243_1023 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_1033 ();
 FILLER_ASAP7_75t_R FILLER_243_1042 ();
 DECAPx1_ASAP7_75t_R FILLER_243_1047 ();
 FILLER_ASAP7_75t_R FILLER_243_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_243_1345 ();
 DECAPx4_ASAP7_75t_R FILLER_243_1367 ();
 DECAPx10_ASAP7_75t_R FILLER_244_2 ();
 DECAPx10_ASAP7_75t_R FILLER_244_50 ();
 DECAPx1_ASAP7_75t_R FILLER_244_72 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_82 ();
 FILLER_ASAP7_75t_R FILLER_244_92 ();
 DECAPx4_ASAP7_75t_R FILLER_244_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_107 ();
 FILLER_ASAP7_75t_R FILLER_244_134 ();
 DECAPx2_ASAP7_75t_R FILLER_244_139 ();
 FILLER_ASAP7_75t_R FILLER_244_145 ();
 DECAPx4_ASAP7_75t_R FILLER_244_153 ();
 DECAPx2_ASAP7_75t_R FILLER_244_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_175 ();
 DECAPx4_ASAP7_75t_R FILLER_244_179 ();
 DECAPx1_ASAP7_75t_R FILLER_244_195 ();
 DECAPx1_ASAP7_75t_R FILLER_244_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_209 ();
 FILLER_ASAP7_75t_R FILLER_244_213 ();
 DECAPx1_ASAP7_75t_R FILLER_244_218 ();
 FILLER_ASAP7_75t_R FILLER_244_228 ();
 DECAPx2_ASAP7_75t_R FILLER_244_236 ();
 DECAPx4_ASAP7_75t_R FILLER_244_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_260 ();
 DECAPx1_ASAP7_75t_R FILLER_244_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_271 ();
 DECAPx6_ASAP7_75t_R FILLER_244_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_289 ();
 DECAPx6_ASAP7_75t_R FILLER_244_298 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_312 ();
 DECAPx6_ASAP7_75t_R FILLER_244_321 ();
 FILLER_ASAP7_75t_R FILLER_244_335 ();
 FILLER_ASAP7_75t_R FILLER_244_363 ();
 FILLER_ASAP7_75t_R FILLER_244_368 ();
 DECAPx2_ASAP7_75t_R FILLER_244_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_384 ();
 DECAPx4_ASAP7_75t_R FILLER_244_391 ();
 DECAPx2_ASAP7_75t_R FILLER_244_407 ();
 FILLER_ASAP7_75t_R FILLER_244_413 ();
 DECAPx4_ASAP7_75t_R FILLER_244_441 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_451 ();
 FILLER_ASAP7_75t_R FILLER_244_460 ();
 FILLER_ASAP7_75t_R FILLER_244_464 ();
 DECAPx1_ASAP7_75t_R FILLER_244_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_476 ();
 DECAPx2_ASAP7_75t_R FILLER_244_480 ();
 DECAPx2_ASAP7_75t_R FILLER_244_494 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_500 ();
 DECAPx1_ASAP7_75t_R FILLER_244_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_513 ();
 FILLER_ASAP7_75t_R FILLER_244_517 ();
 FILLER_ASAP7_75t_R FILLER_244_525 ();
 DECAPx2_ASAP7_75t_R FILLER_244_535 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_541 ();
 DECAPx4_ASAP7_75t_R FILLER_244_570 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_580 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_609 ();
 FILLER_ASAP7_75t_R FILLER_244_620 ();
 DECAPx6_ASAP7_75t_R FILLER_244_628 ();
 FILLER_ASAP7_75t_R FILLER_244_642 ();
 FILLER_ASAP7_75t_R FILLER_244_650 ();
 DECAPx4_ASAP7_75t_R FILLER_244_655 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_665 ();
 DECAPx6_ASAP7_75t_R FILLER_244_674 ();
 DECAPx1_ASAP7_75t_R FILLER_244_688 ();
 DECAPx2_ASAP7_75t_R FILLER_244_695 ();
 DECAPx10_ASAP7_75t_R FILLER_244_704 ();
 DECAPx4_ASAP7_75t_R FILLER_244_726 ();
 DECAPx1_ASAP7_75t_R FILLER_244_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_743 ();
 DECAPx1_ASAP7_75t_R FILLER_244_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_757 ();
 DECAPx6_ASAP7_75t_R FILLER_244_761 ();
 DECAPx1_ASAP7_75t_R FILLER_244_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_779 ();
 DECAPx2_ASAP7_75t_R FILLER_244_794 ();
 DECAPx10_ASAP7_75t_R FILLER_244_814 ();
 DECAPx2_ASAP7_75t_R FILLER_244_836 ();
 FILLER_ASAP7_75t_R FILLER_244_842 ();
 DECAPx6_ASAP7_75t_R FILLER_244_847 ();
 DECAPx2_ASAP7_75t_R FILLER_244_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_867 ();
 FILLER_ASAP7_75t_R FILLER_244_871 ();
 FILLER_ASAP7_75t_R FILLER_244_887 ();
 DECAPx6_ASAP7_75t_R FILLER_244_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_906 ();
 DECAPx2_ASAP7_75t_R FILLER_244_910 ();
 FILLER_ASAP7_75t_R FILLER_244_930 ();
 DECAPx4_ASAP7_75t_R FILLER_244_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_956 ();
 DECAPx4_ASAP7_75t_R FILLER_244_971 ();
 FILLER_ASAP7_75t_R FILLER_244_981 ();
 DECAPx4_ASAP7_75t_R FILLER_244_986 ();
 FILLER_ASAP7_75t_R FILLER_244_996 ();
 DECAPx2_ASAP7_75t_R FILLER_244_1001 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_244_1016 ();
 DECAPx1_ASAP7_75t_R FILLER_244_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1142 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_244_1340 ();
 DECAPx6_ASAP7_75t_R FILLER_244_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_245_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_16 ();
 FILLER_ASAP7_75t_R FILLER_245_25 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_33 ();
 DECAPx2_ASAP7_75t_R FILLER_245_39 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_45 ();
 DECAPx6_ASAP7_75t_R FILLER_245_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_70 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_97 ();
 DECAPx1_ASAP7_75t_R FILLER_245_138 ();
 DECAPx6_ASAP7_75t_R FILLER_245_168 ();
 FILLER_ASAP7_75t_R FILLER_245_182 ();
 DECAPx4_ASAP7_75t_R FILLER_245_210 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_220 ();
 DECAPx4_ASAP7_75t_R FILLER_245_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_239 ();
 FILLER_ASAP7_75t_R FILLER_245_246 ();
 DECAPx6_ASAP7_75t_R FILLER_245_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_268 ();
 DECAPx6_ASAP7_75t_R FILLER_245_275 ();
 FILLER_ASAP7_75t_R FILLER_245_289 ();
 DECAPx2_ASAP7_75t_R FILLER_245_299 ();
 FILLER_ASAP7_75t_R FILLER_245_305 ();
 DECAPx6_ASAP7_75t_R FILLER_245_333 ();
 DECAPx1_ASAP7_75t_R FILLER_245_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_351 ();
 DECAPx6_ASAP7_75t_R FILLER_245_355 ();
 FILLER_ASAP7_75t_R FILLER_245_375 ();
 FILLER_ASAP7_75t_R FILLER_245_383 ();
 FILLER_ASAP7_75t_R FILLER_245_391 ();
 FILLER_ASAP7_75t_R FILLER_245_419 ();
 DECAPx2_ASAP7_75t_R FILLER_245_424 ();
 DECAPx1_ASAP7_75t_R FILLER_245_433 ();
 DECAPx6_ASAP7_75t_R FILLER_245_445 ();
 DECAPx2_ASAP7_75t_R FILLER_245_459 ();
 DECAPx6_ASAP7_75t_R FILLER_245_468 ();
 FILLER_ASAP7_75t_R FILLER_245_482 ();
 FILLER_ASAP7_75t_R FILLER_245_490 ();
 DECAPx10_ASAP7_75t_R FILLER_245_498 ();
 DECAPx2_ASAP7_75t_R FILLER_245_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_526 ();
 FILLER_ASAP7_75t_R FILLER_245_535 ();
 DECAPx1_ASAP7_75t_R FILLER_245_543 ();
 DECAPx2_ASAP7_75t_R FILLER_245_553 ();
 DECAPx2_ASAP7_75t_R FILLER_245_562 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_568 ();
 DECAPx2_ASAP7_75t_R FILLER_245_577 ();
 FILLER_ASAP7_75t_R FILLER_245_583 ();
 DECAPx2_ASAP7_75t_R FILLER_245_591 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_597 ();
 FILLER_ASAP7_75t_R FILLER_245_603 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_608 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_619 ();
 DECAPx4_ASAP7_75t_R FILLER_245_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_638 ();
 FILLER_ASAP7_75t_R FILLER_245_653 ();
 DECAPx2_ASAP7_75t_R FILLER_245_661 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_667 ();
 DECAPx2_ASAP7_75t_R FILLER_245_673 ();
 FILLER_ASAP7_75t_R FILLER_245_679 ();
 DECAPx2_ASAP7_75t_R FILLER_245_695 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_715 ();
 FILLER_ASAP7_75t_R FILLER_245_721 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_737 ();
 DECAPx2_ASAP7_75t_R FILLER_245_754 ();
 FILLER_ASAP7_75t_R FILLER_245_774 ();
 DECAPx2_ASAP7_75t_R FILLER_245_779 ();
 FILLER_ASAP7_75t_R FILLER_245_785 ();
 FILLER_ASAP7_75t_R FILLER_245_790 ();
 DECAPx6_ASAP7_75t_R FILLER_245_795 ();
 DECAPx2_ASAP7_75t_R FILLER_245_812 ();
 DECAPx4_ASAP7_75t_R FILLER_245_821 ();
 DECAPx1_ASAP7_75t_R FILLER_245_834 ();
 DECAPx4_ASAP7_75t_R FILLER_245_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_862 ();
 DECAPx2_ASAP7_75t_R FILLER_245_866 ();
 FILLER_ASAP7_75t_R FILLER_245_872 ();
 DECAPx10_ASAP7_75t_R FILLER_245_877 ();
 FILLER_ASAP7_75t_R FILLER_245_899 ();
 DECAPx6_ASAP7_75t_R FILLER_245_904 ();
 DECAPx2_ASAP7_75t_R FILLER_245_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_924 ();
 DECAPx4_ASAP7_75t_R FILLER_245_927 ();
 DECAPx10_ASAP7_75t_R FILLER_245_940 ();
 DECAPx6_ASAP7_75t_R FILLER_245_962 ();
 DECAPx6_ASAP7_75t_R FILLER_245_979 ();
 DECAPx1_ASAP7_75t_R FILLER_245_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_997 ();
 DECAPx6_ASAP7_75t_R FILLER_245_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_245_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_1021 ();
 DECAPx6_ASAP7_75t_R FILLER_245_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1155 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1177 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1199 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1221 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_245_1353 ();
 FILLER_ASAP7_75t_R FILLER_245_1375 ();
 DECAPx2_ASAP7_75t_R FILLER_246_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_8 ();
 DECAPx2_ASAP7_75t_R FILLER_246_35 ();
 FILLER_ASAP7_75t_R FILLER_246_47 ();
 DECAPx4_ASAP7_75t_R FILLER_246_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_67 ();
 FILLER_ASAP7_75t_R FILLER_246_74 ();
 FILLER_ASAP7_75t_R FILLER_246_83 ();
 FILLER_ASAP7_75t_R FILLER_246_92 ();
 FILLER_ASAP7_75t_R FILLER_246_100 ();
 FILLER_ASAP7_75t_R FILLER_246_117 ();
 DECAPx4_ASAP7_75t_R FILLER_246_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_135 ();
 FILLER_ASAP7_75t_R FILLER_246_158 ();
 DECAPx4_ASAP7_75t_R FILLER_246_163 ();
 FILLER_ASAP7_75t_R FILLER_246_173 ();
 DECAPx6_ASAP7_75t_R FILLER_246_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_195 ();
 FILLER_ASAP7_75t_R FILLER_246_202 ();
 DECAPx1_ASAP7_75t_R FILLER_246_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_211 ();
 DECAPx10_ASAP7_75t_R FILLER_246_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_260 ();
 FILLER_ASAP7_75t_R FILLER_246_287 ();
 FILLER_ASAP7_75t_R FILLER_246_295 ();
 DECAPx2_ASAP7_75t_R FILLER_246_303 ();
 DECAPx2_ASAP7_75t_R FILLER_246_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_321 ();
 FILLER_ASAP7_75t_R FILLER_246_325 ();
 DECAPx4_ASAP7_75t_R FILLER_246_333 ();
 FILLER_ASAP7_75t_R FILLER_246_343 ();
 DECAPx10_ASAP7_75t_R FILLER_246_351 ();
 DECAPx6_ASAP7_75t_R FILLER_246_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_395 ();
 DECAPx2_ASAP7_75t_R FILLER_246_402 ();
 DECAPx4_ASAP7_75t_R FILLER_246_411 ();
 DECAPx2_ASAP7_75t_R FILLER_246_429 ();
 FILLER_ASAP7_75t_R FILLER_246_435 ();
 DECAPx2_ASAP7_75t_R FILLER_246_443 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_246_449 ();
 DECAPx1_ASAP7_75t_R FILLER_246_458 ();
 DECAPx1_ASAP7_75t_R FILLER_246_464 ();
 FILLER_ASAP7_75t_R FILLER_246_474 ();
 DECAPx6_ASAP7_75t_R FILLER_246_482 ();
 DECAPx1_ASAP7_75t_R FILLER_246_496 ();
 FILLER_ASAP7_75t_R FILLER_246_506 ();
 DECAPx2_ASAP7_75t_R FILLER_246_514 ();
 FILLER_ASAP7_75t_R FILLER_246_523 ();
 DECAPx10_ASAP7_75t_R FILLER_246_531 ();
 DECAPx6_ASAP7_75t_R FILLER_246_553 ();
 FILLER_ASAP7_75t_R FILLER_246_567 ();
 DECAPx6_ASAP7_75t_R FILLER_246_595 ();
 DECAPx2_ASAP7_75t_R FILLER_246_615 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_246_621 ();
 DECAPx6_ASAP7_75t_R FILLER_246_630 ();
 DECAPx4_ASAP7_75t_R FILLER_246_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_660 ();
 FILLER_ASAP7_75t_R FILLER_246_675 ();
 DECAPx2_ASAP7_75t_R FILLER_246_680 ();
 DECAPx4_ASAP7_75t_R FILLER_246_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_710 ();
 DECAPx4_ASAP7_75t_R FILLER_246_714 ();
 FILLER_ASAP7_75t_R FILLER_246_724 ();
 DECAPx10_ASAP7_75t_R FILLER_246_729 ();
 DECAPx2_ASAP7_75t_R FILLER_246_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_760 ();
 DECAPx4_ASAP7_75t_R FILLER_246_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_774 ();
 DECAPx2_ASAP7_75t_R FILLER_246_789 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_246_795 ();
 DECAPx6_ASAP7_75t_R FILLER_246_812 ();
 FILLER_ASAP7_75t_R FILLER_246_826 ();
 DECAPx2_ASAP7_75t_R FILLER_246_831 ();
 FILLER_ASAP7_75t_R FILLER_246_840 ();
 DECAPx2_ASAP7_75t_R FILLER_246_845 ();
 FILLER_ASAP7_75t_R FILLER_246_865 ();
 DECAPx6_ASAP7_75t_R FILLER_246_881 ();
 DECAPx1_ASAP7_75t_R FILLER_246_895 ();
 DECAPx10_ASAP7_75t_R FILLER_246_902 ();
 DECAPx1_ASAP7_75t_R FILLER_246_924 ();
 DECAPx1_ASAP7_75t_R FILLER_246_931 ();
 DECAPx10_ASAP7_75t_R FILLER_246_941 ();
 DECAPx4_ASAP7_75t_R FILLER_246_963 ();
 FILLER_ASAP7_75t_R FILLER_246_973 ();
 FILLER_ASAP7_75t_R FILLER_246_981 ();
 DECAPx6_ASAP7_75t_R FILLER_246_989 ();
 DECAPx2_ASAP7_75t_R FILLER_246_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_1009 ();
 DECAPx6_ASAP7_75t_R FILLER_246_1013 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_246_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_246_1341 ();
 DECAPx6_ASAP7_75t_R FILLER_246_1363 ();
 DECAPx4_ASAP7_75t_R FILLER_247_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_12 ();
 DECAPx1_ASAP7_75t_R FILLER_247_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_23 ();
 DECAPx6_ASAP7_75t_R FILLER_247_27 ();
 DECAPx2_ASAP7_75t_R FILLER_247_41 ();
 FILLER_ASAP7_75t_R FILLER_247_53 ();
 DECAPx6_ASAP7_75t_R FILLER_247_61 ();
 DECAPx1_ASAP7_75t_R FILLER_247_81 ();
 FILLER_ASAP7_75t_R FILLER_247_92 ();
 DECAPx2_ASAP7_75t_R FILLER_247_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_107 ();
 FILLER_ASAP7_75t_R FILLER_247_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_142 ();
 DECAPx4_ASAP7_75t_R FILLER_247_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_161 ();
 DECAPx10_ASAP7_75t_R FILLER_247_188 ();
 DECAPx2_ASAP7_75t_R FILLER_247_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_216 ();
 DECAPx1_ASAP7_75t_R FILLER_247_223 ();
 DECAPx4_ASAP7_75t_R FILLER_247_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_240 ();
 FILLER_ASAP7_75t_R FILLER_247_244 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_252 ();
 DECAPx2_ASAP7_75t_R FILLER_247_258 ();
 DECAPx1_ASAP7_75t_R FILLER_247_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_274 ();
 DECAPx10_ASAP7_75t_R FILLER_247_278 ();
 DECAPx1_ASAP7_75t_R FILLER_247_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_304 ();
 DECAPx2_ASAP7_75t_R FILLER_247_311 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_317 ();
 FILLER_ASAP7_75t_R FILLER_247_326 ();
 FILLER_ASAP7_75t_R FILLER_247_336 ();
 DECAPx4_ASAP7_75t_R FILLER_247_344 ();
 DECAPx4_ASAP7_75t_R FILLER_247_360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_370 ();
 DECAPx6_ASAP7_75t_R FILLER_247_381 ();
 FILLER_ASAP7_75t_R FILLER_247_395 ();
 DECAPx4_ASAP7_75t_R FILLER_247_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_413 ();
 DECAPx2_ASAP7_75t_R FILLER_247_417 ();
 FILLER_ASAP7_75t_R FILLER_247_423 ();
 DECAPx2_ASAP7_75t_R FILLER_247_433 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_439 ();
 DECAPx6_ASAP7_75t_R FILLER_247_448 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_462 ();
 DECAPx1_ASAP7_75t_R FILLER_247_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_495 ();
 DECAPx6_ASAP7_75t_R FILLER_247_522 ();
 FILLER_ASAP7_75t_R FILLER_247_542 ();
 DECAPx2_ASAP7_75t_R FILLER_247_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_556 ();
 DECAPx2_ASAP7_75t_R FILLER_247_563 ();
 DECAPx2_ASAP7_75t_R FILLER_247_575 ();
 FILLER_ASAP7_75t_R FILLER_247_581 ();
 DECAPx10_ASAP7_75t_R FILLER_247_586 ();
 DECAPx2_ASAP7_75t_R FILLER_247_608 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_614 ();
 DECAPx6_ASAP7_75t_R FILLER_247_625 ();
 DECAPx2_ASAP7_75t_R FILLER_247_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_645 ();
 DECAPx6_ASAP7_75t_R FILLER_247_649 ();
 DECAPx1_ASAP7_75t_R FILLER_247_663 ();
 FILLER_ASAP7_75t_R FILLER_247_676 ();
 FILLER_ASAP7_75t_R FILLER_247_681 ();
 DECAPx10_ASAP7_75t_R FILLER_247_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_708 ();
 DECAPx2_ASAP7_75t_R FILLER_247_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_729 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_733 ();
 DECAPx6_ASAP7_75t_R FILLER_247_750 ();
 DECAPx2_ASAP7_75t_R FILLER_247_764 ();
 FILLER_ASAP7_75t_R FILLER_247_784 ();
 FILLER_ASAP7_75t_R FILLER_247_789 ();
 DECAPx2_ASAP7_75t_R FILLER_247_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_800 ();
 FILLER_ASAP7_75t_R FILLER_247_815 ();
 FILLER_ASAP7_75t_R FILLER_247_820 ();
 FILLER_ASAP7_75t_R FILLER_247_825 ();
 FILLER_ASAP7_75t_R FILLER_247_841 ();
 FILLER_ASAP7_75t_R FILLER_247_857 ();
 FILLER_ASAP7_75t_R FILLER_247_862 ();
 DECAPx6_ASAP7_75t_R FILLER_247_867 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_881 ();
 DECAPx4_ASAP7_75t_R FILLER_247_887 ();
 FILLER_ASAP7_75t_R FILLER_247_911 ();
 FILLER_ASAP7_75t_R FILLER_247_916 ();
 DECAPx1_ASAP7_75t_R FILLER_247_921 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_927 ();
 DECAPx1_ASAP7_75t_R FILLER_247_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_948 ();
 FILLER_ASAP7_75t_R FILLER_247_952 ();
 FILLER_ASAP7_75t_R FILLER_247_960 ();
 DECAPx1_ASAP7_75t_R FILLER_247_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_972 ();
 DECAPx4_ASAP7_75t_R FILLER_247_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_997 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_247_1021 ();
 FILLER_ASAP7_75t_R FILLER_247_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_247_1351 ();
 DECAPx1_ASAP7_75t_R FILLER_247_1373 ();
 DECAPx10_ASAP7_75t_R FILLER_248_2 ();
 DECAPx6_ASAP7_75t_R FILLER_248_24 ();
 DECAPx1_ASAP7_75t_R FILLER_248_38 ();
 DECAPx1_ASAP7_75t_R FILLER_248_50 ();
 DECAPx2_ASAP7_75t_R FILLER_248_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_66 ();
 FILLER_ASAP7_75t_R FILLER_248_73 ();
 DECAPx1_ASAP7_75t_R FILLER_248_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_87 ();
 FILLER_ASAP7_75t_R FILLER_248_96 ();
 DECAPx4_ASAP7_75t_R FILLER_248_104 ();
 FILLER_ASAP7_75t_R FILLER_248_114 ();
 DECAPx2_ASAP7_75t_R FILLER_248_122 ();
 FILLER_ASAP7_75t_R FILLER_248_134 ();
 FILLER_ASAP7_75t_R FILLER_248_144 ();
 DECAPx6_ASAP7_75t_R FILLER_248_152 ();
 FILLER_ASAP7_75t_R FILLER_248_166 ();
 FILLER_ASAP7_75t_R FILLER_248_174 ();
 DECAPx6_ASAP7_75t_R FILLER_248_179 ();
 DECAPx1_ASAP7_75t_R FILLER_248_193 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_203 ();
 DECAPx10_ASAP7_75t_R FILLER_248_209 ();
 DECAPx2_ASAP7_75t_R FILLER_248_231 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_237 ();
 DECAPx1_ASAP7_75t_R FILLER_248_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_270 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_277 ();
 FILLER_ASAP7_75t_R FILLER_248_286 ();
 DECAPx1_ASAP7_75t_R FILLER_248_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_295 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_322 ();
 DECAPx4_ASAP7_75t_R FILLER_248_333 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_343 ();
 FILLER_ASAP7_75t_R FILLER_248_372 ();
 DECAPx2_ASAP7_75t_R FILLER_248_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_386 ();
 FILLER_ASAP7_75t_R FILLER_248_413 ();
 FILLER_ASAP7_75t_R FILLER_248_421 ();
 DECAPx2_ASAP7_75t_R FILLER_248_429 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_435 ();
 FILLER_ASAP7_75t_R FILLER_248_444 ();
 FILLER_ASAP7_75t_R FILLER_248_453 ();
 DECAPx1_ASAP7_75t_R FILLER_248_458 ();
 DECAPx6_ASAP7_75t_R FILLER_248_464 ();
 FILLER_ASAP7_75t_R FILLER_248_478 ();
 DECAPx2_ASAP7_75t_R FILLER_248_483 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_489 ();
 DECAPx4_ASAP7_75t_R FILLER_248_498 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_508 ();
 DECAPx4_ASAP7_75t_R FILLER_248_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_524 ();
 FILLER_ASAP7_75t_R FILLER_248_528 ();
 DECAPx2_ASAP7_75t_R FILLER_248_538 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_544 ();
 DECAPx1_ASAP7_75t_R FILLER_248_573 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_603 ();
 FILLER_ASAP7_75t_R FILLER_248_609 ();
 FILLER_ASAP7_75t_R FILLER_248_617 ();
 DECAPx6_ASAP7_75t_R FILLER_248_627 ();
 FILLER_ASAP7_75t_R FILLER_248_641 ();
 DECAPx10_ASAP7_75t_R FILLER_248_657 ();
 DECAPx6_ASAP7_75t_R FILLER_248_679 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_693 ();
 DECAPx1_ASAP7_75t_R FILLER_248_702 ();
 DECAPx2_ASAP7_75t_R FILLER_248_709 ();
 FILLER_ASAP7_75t_R FILLER_248_715 ();
 FILLER_ASAP7_75t_R FILLER_248_731 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_747 ();
 FILLER_ASAP7_75t_R FILLER_248_764 ();
 FILLER_ASAP7_75t_R FILLER_248_769 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_785 ();
 DECAPx4_ASAP7_75t_R FILLER_248_791 ();
 FILLER_ASAP7_75t_R FILLER_248_801 ();
 FILLER_ASAP7_75t_R FILLER_248_817 ();
 FILLER_ASAP7_75t_R FILLER_248_822 ();
 DECAPx10_ASAP7_75t_R FILLER_248_827 ();
 DECAPx10_ASAP7_75t_R FILLER_248_849 ();
 FILLER_ASAP7_75t_R FILLER_248_871 ();
 FILLER_ASAP7_75t_R FILLER_248_887 ();
 DECAPx6_ASAP7_75t_R FILLER_248_903 ();
 DECAPx2_ASAP7_75t_R FILLER_248_945 ();
 DECAPx4_ASAP7_75t_R FILLER_248_965 ();
 FILLER_ASAP7_75t_R FILLER_248_975 ();
 DECAPx4_ASAP7_75t_R FILLER_248_983 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_993 ();
 FILLER_ASAP7_75t_R FILLER_248_1010 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_1018 ();
 FILLER_ASAP7_75t_R FILLER_248_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_248_1348 ();
 DECAPx2_ASAP7_75t_R FILLER_248_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_249_2 ();
 DECAPx1_ASAP7_75t_R FILLER_249_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_20 ();
 DECAPx2_ASAP7_75t_R FILLER_249_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_33 ();
 FILLER_ASAP7_75t_R FILLER_249_40 ();
 DECAPx6_ASAP7_75t_R FILLER_249_50 ();
 DECAPx2_ASAP7_75t_R FILLER_249_70 ();
 FILLER_ASAP7_75t_R FILLER_249_82 ();
 DECAPx1_ASAP7_75t_R FILLER_249_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_91 ();
 DECAPx2_ASAP7_75t_R FILLER_249_98 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_249_104 ();
 FILLER_ASAP7_75t_R FILLER_249_113 ();
 FILLER_ASAP7_75t_R FILLER_249_121 ();
 DECAPx2_ASAP7_75t_R FILLER_249_126 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_249_132 ();
 DECAPx4_ASAP7_75t_R FILLER_249_143 ();
 FILLER_ASAP7_75t_R FILLER_249_153 ();
 DECAPx6_ASAP7_75t_R FILLER_249_161 ();
 DECAPx4_ASAP7_75t_R FILLER_249_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_191 ();
 FILLER_ASAP7_75t_R FILLER_249_218 ();
 DECAPx6_ASAP7_75t_R FILLER_249_223 ();
 DECAPx2_ASAP7_75t_R FILLER_249_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_243 ();
 DECAPx2_ASAP7_75t_R FILLER_249_250 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_249_256 ();
 FILLER_ASAP7_75t_R FILLER_249_266 ();
 DECAPx1_ASAP7_75t_R FILLER_249_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_298 ();
 DECAPx2_ASAP7_75t_R FILLER_249_305 ();
 DECAPx2_ASAP7_75t_R FILLER_249_314 ();
 DECAPx2_ASAP7_75t_R FILLER_249_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_329 ();
 DECAPx1_ASAP7_75t_R FILLER_249_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_340 ();
 FILLER_ASAP7_75t_R FILLER_249_347 ();
 DECAPx2_ASAP7_75t_R FILLER_249_355 ();
 DECAPx1_ASAP7_75t_R FILLER_249_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_368 ();
 DECAPx6_ASAP7_75t_R FILLER_249_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_389 ();
 DECAPx2_ASAP7_75t_R FILLER_249_396 ();
 DECAPx2_ASAP7_75t_R FILLER_249_405 ();
 DECAPx6_ASAP7_75t_R FILLER_249_417 ();
 FILLER_ASAP7_75t_R FILLER_249_437 ();
 FILLER_ASAP7_75t_R FILLER_249_465 ();
 DECAPx4_ASAP7_75t_R FILLER_249_473 ();
 FILLER_ASAP7_75t_R FILLER_249_483 ();
 DECAPx4_ASAP7_75t_R FILLER_249_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_521 ();
 FILLER_ASAP7_75t_R FILLER_249_528 ();
 DECAPx6_ASAP7_75t_R FILLER_249_538 ();
 DECAPx1_ASAP7_75t_R FILLER_249_558 ();
 DECAPx4_ASAP7_75t_R FILLER_249_565 ();
 FILLER_ASAP7_75t_R FILLER_249_581 ();
 FILLER_ASAP7_75t_R FILLER_249_589 ();
 FILLER_ASAP7_75t_R FILLER_249_617 ();
 DECAPx10_ASAP7_75t_R FILLER_249_625 ();
 FILLER_ASAP7_75t_R FILLER_249_661 ();
 FILLER_ASAP7_75t_R FILLER_249_669 ();
 FILLER_ASAP7_75t_R FILLER_249_677 ();
 DECAPx1_ASAP7_75t_R FILLER_249_682 ();
 FILLER_ASAP7_75t_R FILLER_249_692 ();
 DECAPx4_ASAP7_75t_R FILLER_249_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_718 ();
 DECAPx2_ASAP7_75t_R FILLER_249_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_728 ();
 DECAPx6_ASAP7_75t_R FILLER_249_732 ();
 DECAPx1_ASAP7_75t_R FILLER_249_746 ();
 DECAPx10_ASAP7_75t_R FILLER_249_753 ();
 DECAPx6_ASAP7_75t_R FILLER_249_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_789 ();
 DECAPx10_ASAP7_75t_R FILLER_249_796 ();
 DECAPx6_ASAP7_75t_R FILLER_249_818 ();
 FILLER_ASAP7_75t_R FILLER_249_832 ();
 DECAPx6_ASAP7_75t_R FILLER_249_837 ();
 DECAPx2_ASAP7_75t_R FILLER_249_851 ();
 FILLER_ASAP7_75t_R FILLER_249_860 ();
 DECAPx4_ASAP7_75t_R FILLER_249_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_875 ();
 DECAPx4_ASAP7_75t_R FILLER_249_879 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_249_889 ();
 FILLER_ASAP7_75t_R FILLER_249_898 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_249_906 ();
 FILLER_ASAP7_75t_R FILLER_249_923 ();
 DECAPx2_ASAP7_75t_R FILLER_249_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_933 ();
 FILLER_ASAP7_75t_R FILLER_249_940 ();
 DECAPx2_ASAP7_75t_R FILLER_249_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_954 ();
 FILLER_ASAP7_75t_R FILLER_249_961 ();
 DECAPx6_ASAP7_75t_R FILLER_249_966 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_249_980 ();
 FILLER_ASAP7_75t_R FILLER_249_986 ();
 DECAPx2_ASAP7_75t_R FILLER_249_991 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_249_997 ();
 FILLER_ASAP7_75t_R FILLER_249_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_249_1011 ();
 DECAPx1_ASAP7_75t_R FILLER_249_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_249_1344 ();
 DECAPx4_ASAP7_75t_R FILLER_249_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_1376 ();
 DECAPx4_ASAP7_75t_R FILLER_250_2 ();
 FILLER_ASAP7_75t_R FILLER_250_38 ();
 DECAPx2_ASAP7_75t_R FILLER_250_46 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_52 ();
 DECAPx6_ASAP7_75t_R FILLER_250_81 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_95 ();
 FILLER_ASAP7_75t_R FILLER_250_124 ();
 DECAPx6_ASAP7_75t_R FILLER_250_129 ();
 DECAPx4_ASAP7_75t_R FILLER_250_149 ();
 DECAPx2_ASAP7_75t_R FILLER_250_165 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_171 ();
 FILLER_ASAP7_75t_R FILLER_250_182 ();
 DECAPx1_ASAP7_75t_R FILLER_250_190 ();
 FILLER_ASAP7_75t_R FILLER_250_200 ();
 DECAPx2_ASAP7_75t_R FILLER_250_208 ();
 FILLER_ASAP7_75t_R FILLER_250_214 ();
 FILLER_ASAP7_75t_R FILLER_250_222 ();
 FILLER_ASAP7_75t_R FILLER_250_232 ();
 DECAPx2_ASAP7_75t_R FILLER_250_240 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_252 ();
 FILLER_ASAP7_75t_R FILLER_250_262 ();
 FILLER_ASAP7_75t_R FILLER_250_271 ();
 FILLER_ASAP7_75t_R FILLER_250_280 ();
 FILLER_ASAP7_75t_R FILLER_250_289 ();
 DECAPx10_ASAP7_75t_R FILLER_250_294 ();
 DECAPx10_ASAP7_75t_R FILLER_250_316 ();
 DECAPx10_ASAP7_75t_R FILLER_250_338 ();
 DECAPx10_ASAP7_75t_R FILLER_250_360 ();
 DECAPx6_ASAP7_75t_R FILLER_250_382 ();
 DECAPx2_ASAP7_75t_R FILLER_250_396 ();
 DECAPx2_ASAP7_75t_R FILLER_250_428 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_434 ();
 FILLER_ASAP7_75t_R FILLER_250_444 ();
 DECAPx2_ASAP7_75t_R FILLER_250_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_459 ();
 FILLER_ASAP7_75t_R FILLER_250_464 ();
 DECAPx6_ASAP7_75t_R FILLER_250_474 ();
 DECAPx1_ASAP7_75t_R FILLER_250_494 ();
 FILLER_ASAP7_75t_R FILLER_250_501 ();
 FILLER_ASAP7_75t_R FILLER_250_509 ();
 DECAPx4_ASAP7_75t_R FILLER_250_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_527 ();
 DECAPx10_ASAP7_75t_R FILLER_250_534 ();
 DECAPx1_ASAP7_75t_R FILLER_250_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_560 ();
 DECAPx4_ASAP7_75t_R FILLER_250_567 ();
 DECAPx2_ASAP7_75t_R FILLER_250_583 ();
 FILLER_ASAP7_75t_R FILLER_250_592 ();
 DECAPx2_ASAP7_75t_R FILLER_250_600 ();
 DECAPx10_ASAP7_75t_R FILLER_250_609 ();
 DECAPx6_ASAP7_75t_R FILLER_250_631 ();
 DECAPx2_ASAP7_75t_R FILLER_250_645 ();
 DECAPx4_ASAP7_75t_R FILLER_250_657 ();
 DECAPx6_ASAP7_75t_R FILLER_250_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_695 ();
 DECAPx1_ASAP7_75t_R FILLER_250_702 ();
 DECAPx2_ASAP7_75t_R FILLER_250_709 ();
 DECAPx10_ASAP7_75t_R FILLER_250_718 ();
 DECAPx4_ASAP7_75t_R FILLER_250_740 ();
 DECAPx10_ASAP7_75t_R FILLER_250_756 ();
 DECAPx6_ASAP7_75t_R FILLER_250_778 ();
 DECAPx4_ASAP7_75t_R FILLER_250_798 ();
 FILLER_ASAP7_75t_R FILLER_250_808 ();
 DECAPx6_ASAP7_75t_R FILLER_250_813 ();
 DECAPx4_ASAP7_75t_R FILLER_250_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_851 ();
 FILLER_ASAP7_75t_R FILLER_250_866 ();
 DECAPx4_ASAP7_75t_R FILLER_250_882 ();
 FILLER_ASAP7_75t_R FILLER_250_892 ();
 DECAPx6_ASAP7_75t_R FILLER_250_900 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_914 ();
 DECAPx10_ASAP7_75t_R FILLER_250_943 ();
 DECAPx6_ASAP7_75t_R FILLER_250_965 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_979 ();
 DECAPx10_ASAP7_75t_R FILLER_250_996 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1040 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1128 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1238 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_250_1348 ();
 DECAPx2_ASAP7_75t_R FILLER_250_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_251_2 ();
 DECAPx1_ASAP7_75t_R FILLER_251_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_26 ();
 DECAPx10_ASAP7_75t_R FILLER_251_30 ();
 DECAPx2_ASAP7_75t_R FILLER_251_52 ();
 DECAPx1_ASAP7_75t_R FILLER_251_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_68 ();
 DECAPx10_ASAP7_75t_R FILLER_251_72 ();
 FILLER_ASAP7_75t_R FILLER_251_124 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_251_129 ();
 FILLER_ASAP7_75t_R FILLER_251_138 ();
 FILLER_ASAP7_75t_R FILLER_251_162 ();
 DECAPx1_ASAP7_75t_R FILLER_251_170 ();
 DECAPx2_ASAP7_75t_R FILLER_251_182 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_251_188 ();
 FILLER_ASAP7_75t_R FILLER_251_217 ();
 FILLER_ASAP7_75t_R FILLER_251_227 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_251_251 ();
 DECAPx1_ASAP7_75t_R FILLER_251_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_264 ();
 DECAPx6_ASAP7_75t_R FILLER_251_273 ();
 DECAPx1_ASAP7_75t_R FILLER_251_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_291 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_251_298 ();
 DECAPx2_ASAP7_75t_R FILLER_251_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_310 ();
 DECAPx2_ASAP7_75t_R FILLER_251_319 ();
 FILLER_ASAP7_75t_R FILLER_251_325 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_251_335 ();
 DECAPx6_ASAP7_75t_R FILLER_251_344 ();
 DECAPx4_ASAP7_75t_R FILLER_251_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_374 ();
 FILLER_ASAP7_75t_R FILLER_251_383 ();
 FILLER_ASAP7_75t_R FILLER_251_391 ();
 DECAPx1_ASAP7_75t_R FILLER_251_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_403 ();
 DECAPx2_ASAP7_75t_R FILLER_251_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_416 ();
 DECAPx4_ASAP7_75t_R FILLER_251_420 ();
 FILLER_ASAP7_75t_R FILLER_251_436 ();
 FILLER_ASAP7_75t_R FILLER_251_444 ();
 DECAPx1_ASAP7_75t_R FILLER_251_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_457 ();
 DECAPx4_ASAP7_75t_R FILLER_251_466 ();
 FILLER_ASAP7_75t_R FILLER_251_476 ();
 DECAPx4_ASAP7_75t_R FILLER_251_486 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_251_496 ();
 DECAPx6_ASAP7_75t_R FILLER_251_525 ();
 FILLER_ASAP7_75t_R FILLER_251_545 ();
 FILLER_ASAP7_75t_R FILLER_251_553 ();
 FILLER_ASAP7_75t_R FILLER_251_561 ();
 FILLER_ASAP7_75t_R FILLER_251_571 ();
 DECAPx10_ASAP7_75t_R FILLER_251_579 ();
 DECAPx4_ASAP7_75t_R FILLER_251_601 ();
 FILLER_ASAP7_75t_R FILLER_251_619 ();
 FILLER_ASAP7_75t_R FILLER_251_627 ();
 DECAPx6_ASAP7_75t_R FILLER_251_635 ();
 FILLER_ASAP7_75t_R FILLER_251_655 ();
 DECAPx4_ASAP7_75t_R FILLER_251_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_670 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_251_677 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_251_683 ();
 DECAPx6_ASAP7_75t_R FILLER_251_689 ();
 DECAPx1_ASAP7_75t_R FILLER_251_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_707 ();
 DECAPx2_ASAP7_75t_R FILLER_251_722 ();
 FILLER_ASAP7_75t_R FILLER_251_742 ();
 DECAPx1_ASAP7_75t_R FILLER_251_747 ();
 DECAPx1_ASAP7_75t_R FILLER_251_757 ();
 FILLER_ASAP7_75t_R FILLER_251_764 ();
 FILLER_ASAP7_75t_R FILLER_251_780 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_251_785 ();
 FILLER_ASAP7_75t_R FILLER_251_802 ();
 DECAPx4_ASAP7_75t_R FILLER_251_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_828 ();
 DECAPx2_ASAP7_75t_R FILLER_251_832 ();
 FILLER_ASAP7_75t_R FILLER_251_838 ();
 DECAPx2_ASAP7_75t_R FILLER_251_843 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_251_849 ();
 DECAPx6_ASAP7_75t_R FILLER_251_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_869 ();
 FILLER_ASAP7_75t_R FILLER_251_876 ();
 DECAPx10_ASAP7_75t_R FILLER_251_884 ();
 DECAPx2_ASAP7_75t_R FILLER_251_906 ();
 FILLER_ASAP7_75t_R FILLER_251_923 ();
 DECAPx2_ASAP7_75t_R FILLER_251_927 ();
 FILLER_ASAP7_75t_R FILLER_251_936 ();
 FILLER_ASAP7_75t_R FILLER_251_941 ();
 DECAPx1_ASAP7_75t_R FILLER_251_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_950 ();
 FILLER_ASAP7_75t_R FILLER_251_957 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_251_965 ();
 DECAPx6_ASAP7_75t_R FILLER_251_971 ();
 DECAPx6_ASAP7_75t_R FILLER_251_988 ();
 DECAPx2_ASAP7_75t_R FILLER_251_1002 ();
 FILLER_ASAP7_75t_R FILLER_251_1011 ();
 FILLER_ASAP7_75t_R FILLER_251_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1024 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1178 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_251_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_1376 ();
 DECAPx6_ASAP7_75t_R FILLER_252_2 ();
 DECAPx2_ASAP7_75t_R FILLER_252_16 ();
 DECAPx1_ASAP7_75t_R FILLER_252_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_32 ();
 FILLER_ASAP7_75t_R FILLER_252_39 ();
 DECAPx10_ASAP7_75t_R FILLER_252_44 ();
 DECAPx4_ASAP7_75t_R FILLER_252_66 ();
 DECAPx1_ASAP7_75t_R FILLER_252_84 ();
 DECAPx6_ASAP7_75t_R FILLER_252_96 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_110 ();
 FILLER_ASAP7_75t_R FILLER_252_135 ();
 FILLER_ASAP7_75t_R FILLER_252_145 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_153 ();
 DECAPx4_ASAP7_75t_R FILLER_252_164 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_174 ();
 DECAPx6_ASAP7_75t_R FILLER_252_180 ();
 DECAPx1_ASAP7_75t_R FILLER_252_194 ();
 FILLER_ASAP7_75t_R FILLER_252_204 ();
 DECAPx4_ASAP7_75t_R FILLER_252_209 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_225 ();
 FILLER_ASAP7_75t_R FILLER_252_236 ();
 FILLER_ASAP7_75t_R FILLER_252_244 ();
 FILLER_ASAP7_75t_R FILLER_252_252 ();
 DECAPx1_ASAP7_75t_R FILLER_252_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_264 ();
 DECAPx6_ASAP7_75t_R FILLER_252_273 ();
 FILLER_ASAP7_75t_R FILLER_252_313 ();
 DECAPx1_ASAP7_75t_R FILLER_252_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_327 ();
 DECAPx2_ASAP7_75t_R FILLER_252_336 ();
 FILLER_ASAP7_75t_R FILLER_252_348 ();
 FILLER_ASAP7_75t_R FILLER_252_376 ();
 DECAPx1_ASAP7_75t_R FILLER_252_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_390 ();
 DECAPx6_ASAP7_75t_R FILLER_252_399 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_413 ();
 DECAPx2_ASAP7_75t_R FILLER_252_422 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_428 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_434 ();
 FILLER_ASAP7_75t_R FILLER_252_445 ();
 DECAPx2_ASAP7_75t_R FILLER_252_454 ();
 FILLER_ASAP7_75t_R FILLER_252_460 ();
 FILLER_ASAP7_75t_R FILLER_252_464 ();
 DECAPx2_ASAP7_75t_R FILLER_252_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_480 ();
 DECAPx10_ASAP7_75t_R FILLER_252_487 ();
 DECAPx1_ASAP7_75t_R FILLER_252_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_513 ();
 DECAPx2_ASAP7_75t_R FILLER_252_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_523 ();
 DECAPx2_ASAP7_75t_R FILLER_252_532 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_538 ();
 DECAPx4_ASAP7_75t_R FILLER_252_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_557 ();
 FILLER_ASAP7_75t_R FILLER_252_566 ();
 DECAPx6_ASAP7_75t_R FILLER_252_574 ();
 FILLER_ASAP7_75t_R FILLER_252_588 ();
 DECAPx4_ASAP7_75t_R FILLER_252_596 ();
 DECAPx1_ASAP7_75t_R FILLER_252_609 ();
 DECAPx2_ASAP7_75t_R FILLER_252_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_627 ();
 FILLER_ASAP7_75t_R FILLER_252_636 ();
 DECAPx10_ASAP7_75t_R FILLER_252_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_668 ();
 DECAPx6_ASAP7_75t_R FILLER_252_675 ();
 FILLER_ASAP7_75t_R FILLER_252_689 ();
 DECAPx1_ASAP7_75t_R FILLER_252_694 ();
 DECAPx4_ASAP7_75t_R FILLER_252_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_711 ();
 FILLER_ASAP7_75t_R FILLER_252_715 ();
 DECAPx2_ASAP7_75t_R FILLER_252_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_737 ();
 DECAPx2_ASAP7_75t_R FILLER_252_741 ();
 DECAPx4_ASAP7_75t_R FILLER_252_761 ();
 FILLER_ASAP7_75t_R FILLER_252_771 ();
 FILLER_ASAP7_75t_R FILLER_252_776 ();
 DECAPx4_ASAP7_75t_R FILLER_252_781 ();
 DECAPx2_ASAP7_75t_R FILLER_252_797 ();
 DECAPx2_ASAP7_75t_R FILLER_252_806 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_812 ();
 DECAPx1_ASAP7_75t_R FILLER_252_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_822 ();
 FILLER_ASAP7_75t_R FILLER_252_829 ();
 DECAPx1_ASAP7_75t_R FILLER_252_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_841 ();
 DECAPx6_ASAP7_75t_R FILLER_252_856 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_870 ();
 DECAPx2_ASAP7_75t_R FILLER_252_879 ();
 FILLER_ASAP7_75t_R FILLER_252_885 ();
 FILLER_ASAP7_75t_R FILLER_252_890 ();
 FILLER_ASAP7_75t_R FILLER_252_895 ();
 FILLER_ASAP7_75t_R FILLER_252_911 ();
 DECAPx2_ASAP7_75t_R FILLER_252_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_922 ();
 DECAPx1_ASAP7_75t_R FILLER_252_929 ();
 FILLER_ASAP7_75t_R FILLER_252_947 ();
 FILLER_ASAP7_75t_R FILLER_252_963 ();
 FILLER_ASAP7_75t_R FILLER_252_979 ();
 DECAPx2_ASAP7_75t_R FILLER_252_984 ();
 FILLER_ASAP7_75t_R FILLER_252_996 ();
 DECAPx2_ASAP7_75t_R FILLER_252_1001 ();
 FILLER_ASAP7_75t_R FILLER_252_1007 ();
 FILLER_ASAP7_75t_R FILLER_252_1023 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_252_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_252_1361 ();
 FILLER_ASAP7_75t_R FILLER_252_1375 ();
 DECAPx6_ASAP7_75t_R FILLER_253_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_16 ();
 DECAPx2_ASAP7_75t_R FILLER_253_45 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_51 ();
 DECAPx4_ASAP7_75t_R FILLER_253_60 ();
 FILLER_ASAP7_75t_R FILLER_253_70 ();
 FILLER_ASAP7_75t_R FILLER_253_75 ();
 DECAPx2_ASAP7_75t_R FILLER_253_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_89 ();
 DECAPx1_ASAP7_75t_R FILLER_253_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_100 ();
 DECAPx2_ASAP7_75t_R FILLER_253_127 ();
 FILLER_ASAP7_75t_R FILLER_253_133 ();
 DECAPx1_ASAP7_75t_R FILLER_253_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_147 ();
 FILLER_ASAP7_75t_R FILLER_253_154 ();
 DECAPx2_ASAP7_75t_R FILLER_253_164 ();
 DECAPx1_ASAP7_75t_R FILLER_253_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_200 ();
 DECAPx6_ASAP7_75t_R FILLER_253_207 ();
 DECAPx2_ASAP7_75t_R FILLER_253_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_227 ();
 DECAPx4_ASAP7_75t_R FILLER_253_236 ();
 DECAPx4_ASAP7_75t_R FILLER_253_254 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_264 ();
 FILLER_ASAP7_75t_R FILLER_253_273 ();
 DECAPx2_ASAP7_75t_R FILLER_253_281 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_287 ();
 DECAPx4_ASAP7_75t_R FILLER_253_296 ();
 FILLER_ASAP7_75t_R FILLER_253_306 ();
 FILLER_ASAP7_75t_R FILLER_253_314 ();
 DECAPx1_ASAP7_75t_R FILLER_253_322 ();
 DECAPx2_ASAP7_75t_R FILLER_253_332 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_338 ();
 DECAPx1_ASAP7_75t_R FILLER_253_349 ();
 DECAPx2_ASAP7_75t_R FILLER_253_359 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_368 ();
 FILLER_ASAP7_75t_R FILLER_253_377 ();
 DECAPx2_ASAP7_75t_R FILLER_253_385 ();
 DECAPx2_ASAP7_75t_R FILLER_253_399 ();
 FILLER_ASAP7_75t_R FILLER_253_405 ();
 DECAPx1_ASAP7_75t_R FILLER_253_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_437 ();
 DECAPx2_ASAP7_75t_R FILLER_253_446 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_452 ();
 FILLER_ASAP7_75t_R FILLER_253_463 ();
 DECAPx2_ASAP7_75t_R FILLER_253_471 ();
 FILLER_ASAP7_75t_R FILLER_253_483 ();
 DECAPx4_ASAP7_75t_R FILLER_253_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_501 ();
 DECAPx2_ASAP7_75t_R FILLER_253_508 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_514 ();
 FILLER_ASAP7_75t_R FILLER_253_523 ();
 DECAPx1_ASAP7_75t_R FILLER_253_533 ();
 DECAPx10_ASAP7_75t_R FILLER_253_545 ();
 DECAPx1_ASAP7_75t_R FILLER_253_567 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_579 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_608 ();
 DECAPx6_ASAP7_75t_R FILLER_253_617 ();
 FILLER_ASAP7_75t_R FILLER_253_637 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_645 ();
 FILLER_ASAP7_75t_R FILLER_253_654 ();
 DECAPx6_ASAP7_75t_R FILLER_253_659 ();
 DECAPx2_ASAP7_75t_R FILLER_253_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_679 ();
 FILLER_ASAP7_75t_R FILLER_253_694 ();
 FILLER_ASAP7_75t_R FILLER_253_705 ();
 DECAPx10_ASAP7_75t_R FILLER_253_710 ();
 DECAPx2_ASAP7_75t_R FILLER_253_732 ();
 DECAPx4_ASAP7_75t_R FILLER_253_741 ();
 DECAPx4_ASAP7_75t_R FILLER_253_757 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_767 ();
 FILLER_ASAP7_75t_R FILLER_253_784 ();
 DECAPx4_ASAP7_75t_R FILLER_253_800 ();
 DECAPx2_ASAP7_75t_R FILLER_253_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_819 ();
 DECAPx4_ASAP7_75t_R FILLER_253_834 ();
 FILLER_ASAP7_75t_R FILLER_253_850 ();
 DECAPx4_ASAP7_75t_R FILLER_253_858 ();
 DECAPx6_ASAP7_75t_R FILLER_253_871 ();
 DECAPx2_ASAP7_75t_R FILLER_253_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_891 ();
 DECAPx4_ASAP7_75t_R FILLER_253_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_916 ();
 FILLER_ASAP7_75t_R FILLER_253_923 ();
 FILLER_ASAP7_75t_R FILLER_253_927 ();
 DECAPx1_ASAP7_75t_R FILLER_253_943 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_950 ();
 DECAPx2_ASAP7_75t_R FILLER_253_959 ();
 DECAPx6_ASAP7_75t_R FILLER_253_968 ();
 DECAPx1_ASAP7_75t_R FILLER_253_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_986 ();
 FILLER_ASAP7_75t_R FILLER_253_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_253_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_253_1351 ();
 DECAPx1_ASAP7_75t_R FILLER_253_1373 ();
 DECAPx10_ASAP7_75t_R FILLER_254_2 ();
 DECAPx2_ASAP7_75t_R FILLER_254_24 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_254_30 ();
 DECAPx4_ASAP7_75t_R FILLER_254_36 ();
 DECAPx2_ASAP7_75t_R FILLER_254_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_78 ();
 FILLER_ASAP7_75t_R FILLER_254_85 ();
 DECAPx4_ASAP7_75t_R FILLER_254_93 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_254_103 ();
 FILLER_ASAP7_75t_R FILLER_254_112 ();
 FILLER_ASAP7_75t_R FILLER_254_120 ();
 DECAPx1_ASAP7_75t_R FILLER_254_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_129 ();
 DECAPx1_ASAP7_75t_R FILLER_254_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_137 ();
 DECAPx2_ASAP7_75t_R FILLER_254_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_150 ();
 DECAPx1_ASAP7_75t_R FILLER_254_154 ();
 DECAPx1_ASAP7_75t_R FILLER_254_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_168 ();
 FILLER_ASAP7_75t_R FILLER_254_175 ();
 DECAPx2_ASAP7_75t_R FILLER_254_183 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_254_189 ();
 FILLER_ASAP7_75t_R FILLER_254_218 ();
 DECAPx1_ASAP7_75t_R FILLER_254_223 ();
 FILLER_ASAP7_75t_R FILLER_254_233 ();
 DECAPx2_ASAP7_75t_R FILLER_254_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_247 ();
 DECAPx4_ASAP7_75t_R FILLER_254_256 ();
 FILLER_ASAP7_75t_R FILLER_254_266 ();
 DECAPx10_ASAP7_75t_R FILLER_254_294 ();
 DECAPx4_ASAP7_75t_R FILLER_254_316 ();
 DECAPx2_ASAP7_75t_R FILLER_254_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_338 ();
 DECAPx4_ASAP7_75t_R FILLER_254_347 ();
 DECAPx1_ASAP7_75t_R FILLER_254_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_367 ();
 DECAPx6_ASAP7_75t_R FILLER_254_374 ();
 DECAPx1_ASAP7_75t_R FILLER_254_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_392 ();
 FILLER_ASAP7_75t_R FILLER_254_399 ();
 DECAPx1_ASAP7_75t_R FILLER_254_407 ();
 DECAPx1_ASAP7_75t_R FILLER_254_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_421 ();
 DECAPx2_ASAP7_75t_R FILLER_254_425 ();
 FILLER_ASAP7_75t_R FILLER_254_437 ();
 DECAPx2_ASAP7_75t_R FILLER_254_445 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_254_451 ();
 FILLER_ASAP7_75t_R FILLER_254_460 ();
 FILLER_ASAP7_75t_R FILLER_254_464 ();
 DECAPx2_ASAP7_75t_R FILLER_254_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_480 ();
 FILLER_ASAP7_75t_R FILLER_254_507 ();
 DECAPx2_ASAP7_75t_R FILLER_254_515 ();
 DECAPx4_ASAP7_75t_R FILLER_254_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_537 ();
 DECAPx6_ASAP7_75t_R FILLER_254_546 ();
 DECAPx1_ASAP7_75t_R FILLER_254_560 ();
 FILLER_ASAP7_75t_R FILLER_254_570 ();
 DECAPx2_ASAP7_75t_R FILLER_254_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_586 ();
 DECAPx1_ASAP7_75t_R FILLER_254_593 ();
 DECAPx2_ASAP7_75t_R FILLER_254_600 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_254_606 ();
 DECAPx10_ASAP7_75t_R FILLER_254_615 ();
 DECAPx1_ASAP7_75t_R FILLER_254_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_641 ();
 DECAPx1_ASAP7_75t_R FILLER_254_656 ();
 DECAPx10_ASAP7_75t_R FILLER_254_674 ();
 DECAPx10_ASAP7_75t_R FILLER_254_696 ();
 DECAPx2_ASAP7_75t_R FILLER_254_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_724 ();
 DECAPx10_ASAP7_75t_R FILLER_254_728 ();
 FILLER_ASAP7_75t_R FILLER_254_750 ();
 FILLER_ASAP7_75t_R FILLER_254_755 ();
 DECAPx10_ASAP7_75t_R FILLER_254_760 ();
 DECAPx10_ASAP7_75t_R FILLER_254_782 ();
 DECAPx6_ASAP7_75t_R FILLER_254_804 ();
 DECAPx2_ASAP7_75t_R FILLER_254_818 ();
 DECAPx6_ASAP7_75t_R FILLER_254_830 ();
 FILLER_ASAP7_75t_R FILLER_254_844 ();
 DECAPx1_ASAP7_75t_R FILLER_254_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_856 ();
 FILLER_ASAP7_75t_R FILLER_254_860 ();
 FILLER_ASAP7_75t_R FILLER_254_876 ();
 FILLER_ASAP7_75t_R FILLER_254_892 ();
 DECAPx2_ASAP7_75t_R FILLER_254_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_903 ();
 FILLER_ASAP7_75t_R FILLER_254_907 ();
 DECAPx2_ASAP7_75t_R FILLER_254_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_924 ();
 DECAPx10_ASAP7_75t_R FILLER_254_931 ();
 DECAPx6_ASAP7_75t_R FILLER_254_953 ();
 FILLER_ASAP7_75t_R FILLER_254_970 ();
 DECAPx6_ASAP7_75t_R FILLER_254_975 ();
 DECAPx1_ASAP7_75t_R FILLER_254_989 ();
 DECAPx10_ASAP7_75t_R FILLER_254_999 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1065 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_254_1351 ();
 DECAPx1_ASAP7_75t_R FILLER_254_1373 ();
 DECAPx10_ASAP7_75t_R FILLER_255_2 ();
 DECAPx10_ASAP7_75t_R FILLER_255_24 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_46 ();
 DECAPx2_ASAP7_75t_R FILLER_255_55 ();
 DECAPx4_ASAP7_75t_R FILLER_255_64 ();
 DECAPx4_ASAP7_75t_R FILLER_255_100 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_110 ();
 DECAPx2_ASAP7_75t_R FILLER_255_119 ();
 FILLER_ASAP7_75t_R FILLER_255_125 ();
 DECAPx1_ASAP7_75t_R FILLER_255_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_157 ();
 DECAPx6_ASAP7_75t_R FILLER_255_164 ();
 DECAPx2_ASAP7_75t_R FILLER_255_178 ();
 DECAPx2_ASAP7_75t_R FILLER_255_187 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_193 ();
 DECAPx1_ASAP7_75t_R FILLER_255_202 ();
 DECAPx10_ASAP7_75t_R FILLER_255_209 ();
 DECAPx6_ASAP7_75t_R FILLER_255_231 ();
 DECAPx1_ASAP7_75t_R FILLER_255_245 ();
 FILLER_ASAP7_75t_R FILLER_255_255 ();
 DECAPx2_ASAP7_75t_R FILLER_255_263 ();
 FILLER_ASAP7_75t_R FILLER_255_269 ();
 FILLER_ASAP7_75t_R FILLER_255_277 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_285 ();
 FILLER_ASAP7_75t_R FILLER_255_314 ();
 FILLER_ASAP7_75t_R FILLER_255_319 ();
 DECAPx6_ASAP7_75t_R FILLER_255_327 ();
 FILLER_ASAP7_75t_R FILLER_255_341 ();
 DECAPx1_ASAP7_75t_R FILLER_255_349 ();
 FILLER_ASAP7_75t_R FILLER_255_379 ();
 DECAPx2_ASAP7_75t_R FILLER_255_384 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_390 ();
 DECAPx10_ASAP7_75t_R FILLER_255_396 ();
 DECAPx4_ASAP7_75t_R FILLER_255_424 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_434 ();
 FILLER_ASAP7_75t_R FILLER_255_443 ();
 DECAPx2_ASAP7_75t_R FILLER_255_448 ();
 DECAPx1_ASAP7_75t_R FILLER_255_460 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_467 ();
 DECAPx2_ASAP7_75t_R FILLER_255_476 ();
 FILLER_ASAP7_75t_R FILLER_255_482 ();
 DECAPx1_ASAP7_75t_R FILLER_255_490 ();
 FILLER_ASAP7_75t_R FILLER_255_497 ();
 DECAPx4_ASAP7_75t_R FILLER_255_525 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_535 ();
 FILLER_ASAP7_75t_R FILLER_255_544 ();
 DECAPx2_ASAP7_75t_R FILLER_255_552 ();
 FILLER_ASAP7_75t_R FILLER_255_564 ();
 DECAPx2_ASAP7_75t_R FILLER_255_569 ();
 DECAPx10_ASAP7_75t_R FILLER_255_581 ();
 DECAPx4_ASAP7_75t_R FILLER_255_603 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_613 ();
 FILLER_ASAP7_75t_R FILLER_255_622 ();
 FILLER_ASAP7_75t_R FILLER_255_630 ();
 DECAPx4_ASAP7_75t_R FILLER_255_635 ();
 FILLER_ASAP7_75t_R FILLER_255_645 ();
 FILLER_ASAP7_75t_R FILLER_255_653 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_661 ();
 FILLER_ASAP7_75t_R FILLER_255_667 ();
 DECAPx2_ASAP7_75t_R FILLER_255_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_681 ();
 DECAPx6_ASAP7_75t_R FILLER_255_685 ();
 DECAPx2_ASAP7_75t_R FILLER_255_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_711 ();
 DECAPx6_ASAP7_75t_R FILLER_255_726 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_740 ();
 DECAPx10_ASAP7_75t_R FILLER_255_757 ();
 DECAPx4_ASAP7_75t_R FILLER_255_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_789 ();
 DECAPx2_ASAP7_75t_R FILLER_255_793 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_799 ();
 FILLER_ASAP7_75t_R FILLER_255_816 ();
 DECAPx10_ASAP7_75t_R FILLER_255_821 ();
 DECAPx10_ASAP7_75t_R FILLER_255_843 ();
 DECAPx6_ASAP7_75t_R FILLER_255_865 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_879 ();
 DECAPx6_ASAP7_75t_R FILLER_255_885 ();
 DECAPx2_ASAP7_75t_R FILLER_255_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_905 ();
 FILLER_ASAP7_75t_R FILLER_255_915 ();
 DECAPx1_ASAP7_75t_R FILLER_255_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_924 ();
 DECAPx6_ASAP7_75t_R FILLER_255_927 ();
 FILLER_ASAP7_75t_R FILLER_255_941 ();
 FILLER_ASAP7_75t_R FILLER_255_946 ();
 DECAPx2_ASAP7_75t_R FILLER_255_951 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_957 ();
 DECAPx1_ASAP7_75t_R FILLER_255_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_978 ();
 DECAPx10_ASAP7_75t_R FILLER_255_993 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_255_1345 ();
 DECAPx4_ASAP7_75t_R FILLER_255_1367 ();
 DECAPx10_ASAP7_75t_R FILLER_256_2 ();
 DECAPx10_ASAP7_75t_R FILLER_256_24 ();
 DECAPx10_ASAP7_75t_R FILLER_256_46 ();
 DECAPx6_ASAP7_75t_R FILLER_256_68 ();
 DECAPx2_ASAP7_75t_R FILLER_256_82 ();
 DECAPx4_ASAP7_75t_R FILLER_256_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_101 ();
 DECAPx1_ASAP7_75t_R FILLER_256_128 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_138 ();
 FILLER_ASAP7_75t_R FILLER_256_144 ();
 DECAPx10_ASAP7_75t_R FILLER_256_172 ();
 DECAPx6_ASAP7_75t_R FILLER_256_194 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_208 ();
 FILLER_ASAP7_75t_R FILLER_256_217 ();
 DECAPx10_ASAP7_75t_R FILLER_256_225 ();
 DECAPx10_ASAP7_75t_R FILLER_256_247 ();
 DECAPx4_ASAP7_75t_R FILLER_256_269 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_279 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_285 ();
 FILLER_ASAP7_75t_R FILLER_256_294 ();
 DECAPx2_ASAP7_75t_R FILLER_256_302 ();
 FILLER_ASAP7_75t_R FILLER_256_308 ();
 DECAPx1_ASAP7_75t_R FILLER_256_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_340 ();
 DECAPx6_ASAP7_75t_R FILLER_256_347 ();
 DECAPx2_ASAP7_75t_R FILLER_256_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_367 ();
 DECAPx6_ASAP7_75t_R FILLER_256_371 ();
 DECAPx2_ASAP7_75t_R FILLER_256_385 ();
 FILLER_ASAP7_75t_R FILLER_256_397 ();
 DECAPx2_ASAP7_75t_R FILLER_256_402 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_408 ();
 DECAPx6_ASAP7_75t_R FILLER_256_437 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_451 ();
 DECAPx1_ASAP7_75t_R FILLER_256_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_461 ();
 DECAPx6_ASAP7_75t_R FILLER_256_464 ();
 DECAPx1_ASAP7_75t_R FILLER_256_478 ();
 DECAPx10_ASAP7_75t_R FILLER_256_488 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_510 ();
 DECAPx10_ASAP7_75t_R FILLER_256_516 ();
 DECAPx1_ASAP7_75t_R FILLER_256_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_542 ();
 DECAPx6_ASAP7_75t_R FILLER_256_569 ();
 DECAPx2_ASAP7_75t_R FILLER_256_583 ();
 FILLER_ASAP7_75t_R FILLER_256_595 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_603 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_609 ();
 DECAPx6_ASAP7_75t_R FILLER_256_638 ();
 FILLER_ASAP7_75t_R FILLER_256_652 ();
 FILLER_ASAP7_75t_R FILLER_256_660 ();
 DECAPx1_ASAP7_75t_R FILLER_256_676 ();
 FILLER_ASAP7_75t_R FILLER_256_694 ();
 DECAPx4_ASAP7_75t_R FILLER_256_710 ();
 FILLER_ASAP7_75t_R FILLER_256_734 ();
 DECAPx1_ASAP7_75t_R FILLER_256_742 ();
 DECAPx1_ASAP7_75t_R FILLER_256_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_759 ();
 DECAPx1_ASAP7_75t_R FILLER_256_763 ();
 FILLER_ASAP7_75t_R FILLER_256_777 ();
 FILLER_ASAP7_75t_R FILLER_256_783 ();
 FILLER_ASAP7_75t_R FILLER_256_788 ();
 DECAPx1_ASAP7_75t_R FILLER_256_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_803 ();
 FILLER_ASAP7_75t_R FILLER_256_818 ();
 FILLER_ASAP7_75t_R FILLER_256_823 ();
 DECAPx2_ASAP7_75t_R FILLER_256_828 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_834 ();
 FILLER_ASAP7_75t_R FILLER_256_851 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_856 ();
 DECAPx4_ASAP7_75t_R FILLER_256_862 ();
 FILLER_ASAP7_75t_R FILLER_256_872 ();
 FILLER_ASAP7_75t_R FILLER_256_877 ();
 DECAPx1_ASAP7_75t_R FILLER_256_888 ();
 FILLER_ASAP7_75t_R FILLER_256_906 ();
 DECAPx10_ASAP7_75t_R FILLER_256_911 ();
 DECAPx1_ASAP7_75t_R FILLER_256_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_937 ();
 FILLER_ASAP7_75t_R FILLER_256_952 ();
 DECAPx1_ASAP7_75t_R FILLER_256_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_972 ();
 DECAPx10_ASAP7_75t_R FILLER_256_987 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_256_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_256_1361 ();
 FILLER_ASAP7_75t_R FILLER_256_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_257_2 ();
 DECAPx10_ASAP7_75t_R FILLER_257_24 ();
 DECAPx10_ASAP7_75t_R FILLER_257_46 ();
 DECAPx10_ASAP7_75t_R FILLER_257_68 ();
 DECAPx6_ASAP7_75t_R FILLER_257_90 ();
 FILLER_ASAP7_75t_R FILLER_257_104 ();
 DECAPx1_ASAP7_75t_R FILLER_257_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_116 ();
 DECAPx10_ASAP7_75t_R FILLER_257_120 ();
 DECAPx4_ASAP7_75t_R FILLER_257_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_152 ();
 FILLER_ASAP7_75t_R FILLER_257_159 ();
 DECAPx10_ASAP7_75t_R FILLER_257_164 ();
 DECAPx6_ASAP7_75t_R FILLER_257_186 ();
 DECAPx2_ASAP7_75t_R FILLER_257_200 ();
 DECAPx4_ASAP7_75t_R FILLER_257_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_242 ();
 DECAPx1_ASAP7_75t_R FILLER_257_246 ();
 DECAPx2_ASAP7_75t_R FILLER_257_256 ();
 FILLER_ASAP7_75t_R FILLER_257_262 ();
 FILLER_ASAP7_75t_R FILLER_257_267 ();
 DECAPx10_ASAP7_75t_R FILLER_257_275 ();
 DECAPx1_ASAP7_75t_R FILLER_257_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_301 ();
 DECAPx2_ASAP7_75t_R FILLER_257_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_311 ();
 DECAPx2_ASAP7_75t_R FILLER_257_318 ();
 DECAPx4_ASAP7_75t_R FILLER_257_327 ();
 DECAPx10_ASAP7_75t_R FILLER_257_340 ();
 DECAPx4_ASAP7_75t_R FILLER_257_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_372 ();
 DECAPx2_ASAP7_75t_R FILLER_257_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_382 ();
 DECAPx1_ASAP7_75t_R FILLER_257_409 ();
 DECAPx2_ASAP7_75t_R FILLER_257_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_425 ();
 DECAPx10_ASAP7_75t_R FILLER_257_429 ();
 DECAPx6_ASAP7_75t_R FILLER_257_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_491 ();
 FILLER_ASAP7_75t_R FILLER_257_518 ();
 DECAPx4_ASAP7_75t_R FILLER_257_523 ();
 DECAPx6_ASAP7_75t_R FILLER_257_536 ();
 DECAPx1_ASAP7_75t_R FILLER_257_550 ();
 FILLER_ASAP7_75t_R FILLER_257_560 ();
 DECAPx1_ASAP7_75t_R FILLER_257_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_569 ();
 DECAPx2_ASAP7_75t_R FILLER_257_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_579 ();
 DECAPx2_ASAP7_75t_R FILLER_257_586 ();
 DECAPx2_ASAP7_75t_R FILLER_257_618 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_257_624 ();
 DECAPx10_ASAP7_75t_R FILLER_257_630 ();
 DECAPx4_ASAP7_75t_R FILLER_257_652 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_257_662 ();
 DECAPx6_ASAP7_75t_R FILLER_257_671 ();
 DECAPx2_ASAP7_75t_R FILLER_257_685 ();
 DECAPx2_ASAP7_75t_R FILLER_257_694 ();
 FILLER_ASAP7_75t_R FILLER_257_706 ();
 DECAPx2_ASAP7_75t_R FILLER_257_714 ();
 FILLER_ASAP7_75t_R FILLER_257_723 ();
 DECAPx1_ASAP7_75t_R FILLER_257_739 ();
 FILLER_ASAP7_75t_R FILLER_257_746 ();
 DECAPx1_ASAP7_75t_R FILLER_257_762 ();
 FILLER_ASAP7_75t_R FILLER_257_772 ();
 FILLER_ASAP7_75t_R FILLER_257_780 ();
 DECAPx4_ASAP7_75t_R FILLER_257_788 ();
 FILLER_ASAP7_75t_R FILLER_257_798 ();
 DECAPx6_ASAP7_75t_R FILLER_257_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_817 ();
 FILLER_ASAP7_75t_R FILLER_257_832 ();
 DECAPx10_ASAP7_75t_R FILLER_257_848 ();
 DECAPx2_ASAP7_75t_R FILLER_257_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_876 ();
 DECAPx4_ASAP7_75t_R FILLER_257_891 ();
 FILLER_ASAP7_75t_R FILLER_257_901 ();
 FILLER_ASAP7_75t_R FILLER_257_906 ();
 DECAPx6_ASAP7_75t_R FILLER_257_911 ();
 FILLER_ASAP7_75t_R FILLER_257_927 ();
 DECAPx2_ASAP7_75t_R FILLER_257_932 ();
 FILLER_ASAP7_75t_R FILLER_257_943 ();
 DECAPx10_ASAP7_75t_R FILLER_257_948 ();
 DECAPx4_ASAP7_75t_R FILLER_257_970 ();
 FILLER_ASAP7_75t_R FILLER_257_980 ();
 FILLER_ASAP7_75t_R FILLER_257_986 ();
 DECAPx10_ASAP7_75t_R FILLER_257_991 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1013 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1057 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_257_1343 ();
 DECAPx4_ASAP7_75t_R FILLER_257_1365 ();
 FILLER_ASAP7_75t_R FILLER_257_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_258_2 ();
 DECAPx10_ASAP7_75t_R FILLER_258_24 ();
 DECAPx10_ASAP7_75t_R FILLER_258_46 ();
 DECAPx10_ASAP7_75t_R FILLER_258_68 ();
 DECAPx10_ASAP7_75t_R FILLER_258_90 ();
 DECAPx10_ASAP7_75t_R FILLER_258_112 ();
 DECAPx10_ASAP7_75t_R FILLER_258_134 ();
 DECAPx10_ASAP7_75t_R FILLER_258_156 ();
 DECAPx10_ASAP7_75t_R FILLER_258_178 ();
 DECAPx6_ASAP7_75t_R FILLER_258_200 ();
 DECAPx2_ASAP7_75t_R FILLER_258_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_220 ();
 FILLER_ASAP7_75t_R FILLER_258_224 ();
 FILLER_ASAP7_75t_R FILLER_258_232 ();
 FILLER_ASAP7_75t_R FILLER_258_260 ();
 DECAPx2_ASAP7_75t_R FILLER_258_288 ();
 DECAPx6_ASAP7_75t_R FILLER_258_300 ();
 DECAPx2_ASAP7_75t_R FILLER_258_314 ();
 DECAPx1_ASAP7_75t_R FILLER_258_323 ();
 DECAPx1_ASAP7_75t_R FILLER_258_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_337 ();
 DECAPx1_ASAP7_75t_R FILLER_258_364 ();
 DECAPx4_ASAP7_75t_R FILLER_258_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_384 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_258_391 ();
 DECAPx4_ASAP7_75t_R FILLER_258_400 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_258_410 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_258_439 ();
 DECAPx1_ASAP7_75t_R FILLER_258_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_452 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_258_459 ();
 FILLER_ASAP7_75t_R FILLER_258_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_258_472 ();
 DECAPx2_ASAP7_75t_R FILLER_258_481 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_258_487 ();
 FILLER_ASAP7_75t_R FILLER_258_496 ();
 DECAPx1_ASAP7_75t_R FILLER_258_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_508 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_258_535 ();
 DECAPx6_ASAP7_75t_R FILLER_258_544 ();
 DECAPx1_ASAP7_75t_R FILLER_258_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_562 ();
 DECAPx2_ASAP7_75t_R FILLER_258_569 ();
 DECAPx10_ASAP7_75t_R FILLER_258_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_623 ();
 DECAPx10_ASAP7_75t_R FILLER_258_630 ();
 DECAPx2_ASAP7_75t_R FILLER_258_652 ();
 DECAPx6_ASAP7_75t_R FILLER_258_664 ();
 FILLER_ASAP7_75t_R FILLER_258_678 ();
 DECAPx10_ASAP7_75t_R FILLER_258_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_708 ();
 DECAPx6_ASAP7_75t_R FILLER_258_712 ();
 DECAPx1_ASAP7_75t_R FILLER_258_726 ();
 DECAPx10_ASAP7_75t_R FILLER_258_736 ();
 DECAPx2_ASAP7_75t_R FILLER_258_758 ();
 FILLER_ASAP7_75t_R FILLER_258_778 ();
 FILLER_ASAP7_75t_R FILLER_258_794 ();
 DECAPx2_ASAP7_75t_R FILLER_258_810 ();
 DECAPx4_ASAP7_75t_R FILLER_258_825 ();
 FILLER_ASAP7_75t_R FILLER_258_838 ();
 DECAPx2_ASAP7_75t_R FILLER_258_843 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_258_849 ();
 FILLER_ASAP7_75t_R FILLER_258_866 ();
 FILLER_ASAP7_75t_R FILLER_258_872 ();
 DECAPx10_ASAP7_75t_R FILLER_258_878 ();
 DECAPx2_ASAP7_75t_R FILLER_258_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_906 ();
 DECAPx2_ASAP7_75t_R FILLER_258_910 ();
 DECAPx4_ASAP7_75t_R FILLER_258_919 ();
 DECAPx10_ASAP7_75t_R FILLER_258_943 ();
 DECAPx10_ASAP7_75t_R FILLER_258_965 ();
 DECAPx10_ASAP7_75t_R FILLER_258_987 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1031 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1053 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_258_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_258_1361 ();
 FILLER_ASAP7_75t_R FILLER_258_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_259_2 ();
 DECAPx10_ASAP7_75t_R FILLER_259_24 ();
 DECAPx10_ASAP7_75t_R FILLER_259_46 ();
 DECAPx10_ASAP7_75t_R FILLER_259_68 ();
 DECAPx10_ASAP7_75t_R FILLER_259_90 ();
 DECAPx10_ASAP7_75t_R FILLER_259_112 ();
 DECAPx10_ASAP7_75t_R FILLER_259_134 ();
 DECAPx10_ASAP7_75t_R FILLER_259_156 ();
 DECAPx10_ASAP7_75t_R FILLER_259_178 ();
 DECAPx6_ASAP7_75t_R FILLER_259_200 ();
 DECAPx1_ASAP7_75t_R FILLER_259_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_218 ();
 FILLER_ASAP7_75t_R FILLER_259_245 ();
 FILLER_ASAP7_75t_R FILLER_259_253 ();
 DECAPx2_ASAP7_75t_R FILLER_259_258 ();
 FILLER_ASAP7_75t_R FILLER_259_264 ();
 DECAPx1_ASAP7_75t_R FILLER_259_272 ();
 DECAPx2_ASAP7_75t_R FILLER_259_279 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_259_285 ();
 FILLER_ASAP7_75t_R FILLER_259_314 ();
 FILLER_ASAP7_75t_R FILLER_259_342 ();
 FILLER_ASAP7_75t_R FILLER_259_350 ();
 FILLER_ASAP7_75t_R FILLER_259_378 ();
 DECAPx1_ASAP7_75t_R FILLER_259_406 ();
 FILLER_ASAP7_75t_R FILLER_259_416 ();
 DECAPx2_ASAP7_75t_R FILLER_259_424 ();
 FILLER_ASAP7_75t_R FILLER_259_430 ();
 DECAPx2_ASAP7_75t_R FILLER_259_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_259_468 ();
 DECAPx2_ASAP7_75t_R FILLER_259_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_503 ();
 FILLER_ASAP7_75t_R FILLER_259_507 ();
 FILLER_ASAP7_75t_R FILLER_259_515 ();
 FILLER_ASAP7_75t_R FILLER_259_523 ();
 FILLER_ASAP7_75t_R FILLER_259_551 ();
 FILLER_ASAP7_75t_R FILLER_259_579 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_259_587 ();
 DECAPx10_ASAP7_75t_R FILLER_259_593 ();
 DECAPx2_ASAP7_75t_R FILLER_259_641 ();
 FILLER_ASAP7_75t_R FILLER_259_647 ();
 FILLER_ASAP7_75t_R FILLER_259_655 ();
 DECAPx2_ASAP7_75t_R FILLER_259_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_677 ();
 DECAPx4_ASAP7_75t_R FILLER_259_692 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_259_702 ();
 DECAPx6_ASAP7_75t_R FILLER_259_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_725 ();
 DECAPx4_ASAP7_75t_R FILLER_259_732 ();
 FILLER_ASAP7_75t_R FILLER_259_742 ();
 DECAPx10_ASAP7_75t_R FILLER_259_747 ();
 DECAPx6_ASAP7_75t_R FILLER_259_769 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_259_783 ();
 DECAPx2_ASAP7_75t_R FILLER_259_789 ();
 FILLER_ASAP7_75t_R FILLER_259_795 ();
 DECAPx6_ASAP7_75t_R FILLER_259_803 ();
 DECAPx2_ASAP7_75t_R FILLER_259_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_823 ();
 DECAPx10_ASAP7_75t_R FILLER_259_827 ();
 DECAPx10_ASAP7_75t_R FILLER_259_858 ();
 FILLER_ASAP7_75t_R FILLER_259_880 ();
 FILLER_ASAP7_75t_R FILLER_259_896 ();
 DECAPx2_ASAP7_75t_R FILLER_259_901 ();
 DECAPx1_ASAP7_75t_R FILLER_259_921 ();
 DECAPx2_ASAP7_75t_R FILLER_259_927 ();
 DECAPx2_ASAP7_75t_R FILLER_259_936 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_259_945 ();
 FILLER_ASAP7_75t_R FILLER_259_958 ();
 DECAPx2_ASAP7_75t_R FILLER_259_966 ();
 FILLER_ASAP7_75t_R FILLER_259_972 ();
 DECAPx10_ASAP7_75t_R FILLER_259_988 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1010 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1142 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_259_1340 ();
 DECAPx6_ASAP7_75t_R FILLER_259_1362 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_260_2 ();
 DECAPx10_ASAP7_75t_R FILLER_260_24 ();
 DECAPx10_ASAP7_75t_R FILLER_260_46 ();
 DECAPx10_ASAP7_75t_R FILLER_260_68 ();
 DECAPx10_ASAP7_75t_R FILLER_260_90 ();
 DECAPx10_ASAP7_75t_R FILLER_260_112 ();
 DECAPx10_ASAP7_75t_R FILLER_260_134 ();
 DECAPx10_ASAP7_75t_R FILLER_260_156 ();
 DECAPx10_ASAP7_75t_R FILLER_260_178 ();
 DECAPx10_ASAP7_75t_R FILLER_260_200 ();
 FILLER_ASAP7_75t_R FILLER_260_222 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_260_230 ();
 DECAPx10_ASAP7_75t_R FILLER_260_236 ();
 DECAPx10_ASAP7_75t_R FILLER_260_258 ();
 DECAPx6_ASAP7_75t_R FILLER_260_280 ();
 DECAPx1_ASAP7_75t_R FILLER_260_294 ();
 FILLER_ASAP7_75t_R FILLER_260_304 ();
 DECAPx4_ASAP7_75t_R FILLER_260_309 ();
 DECAPx1_ASAP7_75t_R FILLER_260_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_329 ();
 DECAPx2_ASAP7_75t_R FILLER_260_333 ();
 FILLER_ASAP7_75t_R FILLER_260_339 ();
 DECAPx2_ASAP7_75t_R FILLER_260_347 ();
 FILLER_ASAP7_75t_R FILLER_260_356 ();
 DECAPx2_ASAP7_75t_R FILLER_260_364 ();
 DECAPx4_ASAP7_75t_R FILLER_260_373 ();
 DECAPx2_ASAP7_75t_R FILLER_260_389 ();
 DECAPx10_ASAP7_75t_R FILLER_260_398 ();
 DECAPx2_ASAP7_75t_R FILLER_260_420 ();
 FILLER_ASAP7_75t_R FILLER_260_426 ();
 DECAPx1_ASAP7_75t_R FILLER_260_431 ();
 DECAPx2_ASAP7_75t_R FILLER_260_441 ();
 DECAPx4_ASAP7_75t_R FILLER_260_450 ();
 FILLER_ASAP7_75t_R FILLER_260_460 ();
 DECAPx2_ASAP7_75t_R FILLER_260_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_260_470 ();
 DECAPx2_ASAP7_75t_R FILLER_260_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_485 ();
 DECAPx10_ASAP7_75t_R FILLER_260_489 ();
 DECAPx4_ASAP7_75t_R FILLER_260_511 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_260_521 ();
 DECAPx2_ASAP7_75t_R FILLER_260_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_533 ();
 DECAPx1_ASAP7_75t_R FILLER_260_540 ();
 DECAPx4_ASAP7_75t_R FILLER_260_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_557 ();
 DECAPx1_ASAP7_75t_R FILLER_260_564 ();
 DECAPx10_ASAP7_75t_R FILLER_260_571 ();
 DECAPx10_ASAP7_75t_R FILLER_260_593 ();
 DECAPx1_ASAP7_75t_R FILLER_260_615 ();
 DECAPx1_ASAP7_75t_R FILLER_260_625 ();
 DECAPx10_ASAP7_75t_R FILLER_260_632 ();
 DECAPx1_ASAP7_75t_R FILLER_260_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_658 ();
 DECAPx6_ASAP7_75t_R FILLER_260_665 ();
 FILLER_ASAP7_75t_R FILLER_260_685 ();
 DECAPx4_ASAP7_75t_R FILLER_260_693 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_260_703 ();
 FILLER_ASAP7_75t_R FILLER_260_720 ();
 DECAPx2_ASAP7_75t_R FILLER_260_725 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_260_731 ();
 FILLER_ASAP7_75t_R FILLER_260_748 ();
 DECAPx10_ASAP7_75t_R FILLER_260_753 ();
 DECAPx6_ASAP7_75t_R FILLER_260_775 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_260_789 ();
 DECAPx4_ASAP7_75t_R FILLER_260_806 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_260_816 ();
 FILLER_ASAP7_75t_R FILLER_260_825 ();
 DECAPx2_ASAP7_75t_R FILLER_260_833 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_260_849 ();
 FILLER_ASAP7_75t_R FILLER_260_858 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_260_863 ();
 DECAPx1_ASAP7_75t_R FILLER_260_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_876 ();
 DECAPx10_ASAP7_75t_R FILLER_260_883 ();
 DECAPx4_ASAP7_75t_R FILLER_260_905 ();
 FILLER_ASAP7_75t_R FILLER_260_915 ();
 DECAPx4_ASAP7_75t_R FILLER_260_920 ();
 FILLER_ASAP7_75t_R FILLER_260_936 ();
 DECAPx1_ASAP7_75t_R FILLER_260_944 ();
 FILLER_ASAP7_75t_R FILLER_260_962 ();
 FILLER_ASAP7_75t_R FILLER_260_978 ();
 DECAPx10_ASAP7_75t_R FILLER_260_986 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1008 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1184 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_260_1338 ();
 DECAPx6_ASAP7_75t_R FILLER_260_1360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_260_1374 ();
 DECAPx10_ASAP7_75t_R FILLER_261_2 ();
 DECAPx10_ASAP7_75t_R FILLER_261_24 ();
 DECAPx10_ASAP7_75t_R FILLER_261_46 ();
 DECAPx10_ASAP7_75t_R FILLER_261_68 ();
 DECAPx10_ASAP7_75t_R FILLER_261_90 ();
 DECAPx10_ASAP7_75t_R FILLER_261_112 ();
 DECAPx10_ASAP7_75t_R FILLER_261_134 ();
 DECAPx10_ASAP7_75t_R FILLER_261_156 ();
 DECAPx10_ASAP7_75t_R FILLER_261_178 ();
 DECAPx10_ASAP7_75t_R FILLER_261_200 ();
 DECAPx10_ASAP7_75t_R FILLER_261_222 ();
 DECAPx10_ASAP7_75t_R FILLER_261_244 ();
 DECAPx10_ASAP7_75t_R FILLER_261_266 ();
 DECAPx10_ASAP7_75t_R FILLER_261_288 ();
 DECAPx10_ASAP7_75t_R FILLER_261_310 ();
 DECAPx10_ASAP7_75t_R FILLER_261_332 ();
 DECAPx10_ASAP7_75t_R FILLER_261_354 ();
 DECAPx10_ASAP7_75t_R FILLER_261_376 ();
 DECAPx10_ASAP7_75t_R FILLER_261_398 ();
 DECAPx10_ASAP7_75t_R FILLER_261_420 ();
 DECAPx10_ASAP7_75t_R FILLER_261_442 ();
 DECAPx10_ASAP7_75t_R FILLER_261_464 ();
 DECAPx10_ASAP7_75t_R FILLER_261_486 ();
 DECAPx10_ASAP7_75t_R FILLER_261_508 ();
 DECAPx10_ASAP7_75t_R FILLER_261_530 ();
 DECAPx10_ASAP7_75t_R FILLER_261_552 ();
 DECAPx10_ASAP7_75t_R FILLER_261_574 ();
 DECAPx10_ASAP7_75t_R FILLER_261_596 ();
 DECAPx10_ASAP7_75t_R FILLER_261_618 ();
 DECAPx10_ASAP7_75t_R FILLER_261_640 ();
 DECAPx10_ASAP7_75t_R FILLER_261_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_684 ();
 FILLER_ASAP7_75t_R FILLER_261_691 ();
 DECAPx2_ASAP7_75t_R FILLER_261_696 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_261_702 ();
 FILLER_ASAP7_75t_R FILLER_261_711 ();
 DECAPx2_ASAP7_75t_R FILLER_261_727 ();
 DECAPx4_ASAP7_75t_R FILLER_261_736 ();
 DECAPx1_ASAP7_75t_R FILLER_261_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_753 ();
 FILLER_ASAP7_75t_R FILLER_261_760 ();
 FILLER_ASAP7_75t_R FILLER_261_768 ();
 DECAPx6_ASAP7_75t_R FILLER_261_773 ();
 DECAPx2_ASAP7_75t_R FILLER_261_787 ();
 FILLER_ASAP7_75t_R FILLER_261_799 ();
 DECAPx4_ASAP7_75t_R FILLER_261_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_817 ();
 DECAPx6_ASAP7_75t_R FILLER_261_832 ();
 DECAPx1_ASAP7_75t_R FILLER_261_846 ();
 DECAPx4_ASAP7_75t_R FILLER_261_864 ();
 FILLER_ASAP7_75t_R FILLER_261_874 ();
 FILLER_ASAP7_75t_R FILLER_261_890 ();
 DECAPx6_ASAP7_75t_R FILLER_261_895 ();
 DECAPx1_ASAP7_75t_R FILLER_261_909 ();
 DECAPx2_ASAP7_75t_R FILLER_261_916 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_261_922 ();
 FILLER_ASAP7_75t_R FILLER_261_927 ();
 DECAPx2_ASAP7_75t_R FILLER_261_943 ();
 FILLER_ASAP7_75t_R FILLER_261_949 ();
 FILLER_ASAP7_75t_R FILLER_261_957 ();
 DECAPx1_ASAP7_75t_R FILLER_261_965 ();
 FILLER_ASAP7_75t_R FILLER_261_975 ();
 FILLER_ASAP7_75t_R FILLER_261_980 ();
 DECAPx10_ASAP7_75t_R FILLER_261_985 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1007 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1029 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1051 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_261_1337 ();
 DECAPx4_ASAP7_75t_R FILLER_261_1359 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_261_1374 ();
 DECAPx10_ASAP7_75t_R FILLER_262_2 ();
 DECAPx10_ASAP7_75t_R FILLER_262_24 ();
 DECAPx10_ASAP7_75t_R FILLER_262_46 ();
 DECAPx10_ASAP7_75t_R FILLER_262_68 ();
 DECAPx10_ASAP7_75t_R FILLER_262_90 ();
 DECAPx10_ASAP7_75t_R FILLER_262_112 ();
 DECAPx10_ASAP7_75t_R FILLER_262_134 ();
 DECAPx10_ASAP7_75t_R FILLER_262_156 ();
 DECAPx10_ASAP7_75t_R FILLER_262_178 ();
 DECAPx10_ASAP7_75t_R FILLER_262_200 ();
 DECAPx10_ASAP7_75t_R FILLER_262_222 ();
 DECAPx10_ASAP7_75t_R FILLER_262_244 ();
 DECAPx10_ASAP7_75t_R FILLER_262_266 ();
 DECAPx10_ASAP7_75t_R FILLER_262_288 ();
 DECAPx10_ASAP7_75t_R FILLER_262_310 ();
 DECAPx10_ASAP7_75t_R FILLER_262_332 ();
 DECAPx10_ASAP7_75t_R FILLER_262_354 ();
 DECAPx10_ASAP7_75t_R FILLER_262_376 ();
 DECAPx10_ASAP7_75t_R FILLER_262_398 ();
 DECAPx10_ASAP7_75t_R FILLER_262_420 ();
 DECAPx6_ASAP7_75t_R FILLER_262_442 ();
 DECAPx2_ASAP7_75t_R FILLER_262_456 ();
 DECAPx10_ASAP7_75t_R FILLER_262_464 ();
 DECAPx10_ASAP7_75t_R FILLER_262_486 ();
 DECAPx10_ASAP7_75t_R FILLER_262_508 ();
 DECAPx10_ASAP7_75t_R FILLER_262_530 ();
 DECAPx10_ASAP7_75t_R FILLER_262_552 ();
 DECAPx10_ASAP7_75t_R FILLER_262_574 ();
 DECAPx10_ASAP7_75t_R FILLER_262_596 ();
 DECAPx10_ASAP7_75t_R FILLER_262_618 ();
 DECAPx10_ASAP7_75t_R FILLER_262_640 ();
 DECAPx6_ASAP7_75t_R FILLER_262_662 ();
 DECAPx2_ASAP7_75t_R FILLER_262_676 ();
 FILLER_ASAP7_75t_R FILLER_262_696 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_262_701 ();
 DECAPx10_ASAP7_75t_R FILLER_262_710 ();
 DECAPx6_ASAP7_75t_R FILLER_262_732 ();
 DECAPx1_ASAP7_75t_R FILLER_262_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_750 ();
 DECAPx4_ASAP7_75t_R FILLER_262_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_775 ();
 FILLER_ASAP7_75t_R FILLER_262_782 ();
 DECAPx6_ASAP7_75t_R FILLER_262_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_801 ();
 DECAPx6_ASAP7_75t_R FILLER_262_805 ();
 DECAPx1_ASAP7_75t_R FILLER_262_819 ();
 DECAPx10_ASAP7_75t_R FILLER_262_829 ();
 DECAPx1_ASAP7_75t_R FILLER_262_851 ();
 DECAPx6_ASAP7_75t_R FILLER_262_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_875 ();
 FILLER_ASAP7_75t_R FILLER_262_882 ();
 DECAPx4_ASAP7_75t_R FILLER_262_887 ();
 DECAPx4_ASAP7_75t_R FILLER_262_900 ();
 FILLER_ASAP7_75t_R FILLER_262_916 ();
 DECAPx2_ASAP7_75t_R FILLER_262_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_930 ();
 DECAPx10_ASAP7_75t_R FILLER_262_937 ();
 DECAPx10_ASAP7_75t_R FILLER_262_959 ();
 DECAPx10_ASAP7_75t_R FILLER_262_981 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1157 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1179 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_262_1333 ();
 DECAPx2_ASAP7_75t_R FILLER_262_1355 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_262_1361 ();
 FILLER_ASAP7_75t_R FILLER_262_1367 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_262_1374 ();
 DECAPx10_ASAP7_75t_R FILLER_263_2 ();
 DECAPx10_ASAP7_75t_R FILLER_263_24 ();
 DECAPx10_ASAP7_75t_R FILLER_263_46 ();
 DECAPx10_ASAP7_75t_R FILLER_263_68 ();
 DECAPx10_ASAP7_75t_R FILLER_263_90 ();
 DECAPx10_ASAP7_75t_R FILLER_263_112 ();
 DECAPx10_ASAP7_75t_R FILLER_263_134 ();
 DECAPx10_ASAP7_75t_R FILLER_263_156 ();
 DECAPx10_ASAP7_75t_R FILLER_263_178 ();
 DECAPx10_ASAP7_75t_R FILLER_263_200 ();
 DECAPx10_ASAP7_75t_R FILLER_263_222 ();
 DECAPx10_ASAP7_75t_R FILLER_263_244 ();
 DECAPx10_ASAP7_75t_R FILLER_263_266 ();
 DECAPx10_ASAP7_75t_R FILLER_263_288 ();
 DECAPx10_ASAP7_75t_R FILLER_263_310 ();
 DECAPx10_ASAP7_75t_R FILLER_263_332 ();
 DECAPx10_ASAP7_75t_R FILLER_263_354 ();
 DECAPx10_ASAP7_75t_R FILLER_263_376 ();
 DECAPx10_ASAP7_75t_R FILLER_263_398 ();
 DECAPx10_ASAP7_75t_R FILLER_263_420 ();
 DECAPx10_ASAP7_75t_R FILLER_263_442 ();
 DECAPx10_ASAP7_75t_R FILLER_263_464 ();
 DECAPx10_ASAP7_75t_R FILLER_263_486 ();
 DECAPx10_ASAP7_75t_R FILLER_263_508 ();
 DECAPx10_ASAP7_75t_R FILLER_263_530 ();
 DECAPx10_ASAP7_75t_R FILLER_263_552 ();
 DECAPx10_ASAP7_75t_R FILLER_263_574 ();
 DECAPx10_ASAP7_75t_R FILLER_263_596 ();
 DECAPx10_ASAP7_75t_R FILLER_263_618 ();
 DECAPx10_ASAP7_75t_R FILLER_263_640 ();
 DECAPx6_ASAP7_75t_R FILLER_263_662 ();
 FILLER_ASAP7_75t_R FILLER_263_676 ();
 FILLER_ASAP7_75t_R FILLER_263_684 ();
 DECAPx10_ASAP7_75t_R FILLER_263_692 ();
 DECAPx2_ASAP7_75t_R FILLER_263_714 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_263_720 ();
 FILLER_ASAP7_75t_R FILLER_263_726 ();
 FILLER_ASAP7_75t_R FILLER_263_734 ();
 DECAPx4_ASAP7_75t_R FILLER_263_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_752 ();
 FILLER_ASAP7_75t_R FILLER_263_767 ();
 DECAPx1_ASAP7_75t_R FILLER_263_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_776 ();
 DECAPx2_ASAP7_75t_R FILLER_263_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_789 ();
 FILLER_ASAP7_75t_R FILLER_263_804 ();
 DECAPx2_ASAP7_75t_R FILLER_263_812 ();
 FILLER_ASAP7_75t_R FILLER_263_818 ();
 FILLER_ASAP7_75t_R FILLER_263_823 ();
 DECAPx2_ASAP7_75t_R FILLER_263_828 ();
 FILLER_ASAP7_75t_R FILLER_263_837 ();
 DECAPx1_ASAP7_75t_R FILLER_263_845 ();
 DECAPx2_ASAP7_75t_R FILLER_263_852 ();
 DECAPx6_ASAP7_75t_R FILLER_263_861 ();
 DECAPx4_ASAP7_75t_R FILLER_263_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_891 ();
 FILLER_ASAP7_75t_R FILLER_263_895 ();
 DECAPx2_ASAP7_75t_R FILLER_263_900 ();
 DECAPx1_ASAP7_75t_R FILLER_263_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_924 ();
 DECAPx10_ASAP7_75t_R FILLER_263_927 ();
 DECAPx10_ASAP7_75t_R FILLER_263_949 ();
 DECAPx10_ASAP7_75t_R FILLER_263_971 ();
 DECAPx10_ASAP7_75t_R FILLER_263_993 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_263_1323 ();
 DECAPx6_ASAP7_75t_R FILLER_263_1345 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_263_1359 ();
 FILLER_ASAP7_75t_R FILLER_263_1367 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_263_1374 ();
 DECAPx10_ASAP7_75t_R FILLER_264_2 ();
 DECAPx10_ASAP7_75t_R FILLER_264_24 ();
 DECAPx10_ASAP7_75t_R FILLER_264_46 ();
 DECAPx10_ASAP7_75t_R FILLER_264_68 ();
 DECAPx10_ASAP7_75t_R FILLER_264_90 ();
 DECAPx10_ASAP7_75t_R FILLER_264_112 ();
 DECAPx10_ASAP7_75t_R FILLER_264_134 ();
 DECAPx10_ASAP7_75t_R FILLER_264_156 ();
 DECAPx10_ASAP7_75t_R FILLER_264_178 ();
 DECAPx10_ASAP7_75t_R FILLER_264_200 ();
 DECAPx10_ASAP7_75t_R FILLER_264_222 ();
 DECAPx10_ASAP7_75t_R FILLER_264_244 ();
 DECAPx10_ASAP7_75t_R FILLER_264_266 ();
 DECAPx10_ASAP7_75t_R FILLER_264_288 ();
 DECAPx10_ASAP7_75t_R FILLER_264_310 ();
 DECAPx10_ASAP7_75t_R FILLER_264_332 ();
 DECAPx10_ASAP7_75t_R FILLER_264_354 ();
 DECAPx10_ASAP7_75t_R FILLER_264_376 ();
 DECAPx10_ASAP7_75t_R FILLER_264_398 ();
 DECAPx10_ASAP7_75t_R FILLER_264_420 ();
 DECAPx6_ASAP7_75t_R FILLER_264_442 ();
 DECAPx2_ASAP7_75t_R FILLER_264_456 ();
 DECAPx10_ASAP7_75t_R FILLER_264_464 ();
 DECAPx10_ASAP7_75t_R FILLER_264_486 ();
 DECAPx10_ASAP7_75t_R FILLER_264_508 ();
 DECAPx10_ASAP7_75t_R FILLER_264_530 ();
 DECAPx10_ASAP7_75t_R FILLER_264_552 ();
 DECAPx10_ASAP7_75t_R FILLER_264_574 ();
 DECAPx10_ASAP7_75t_R FILLER_264_596 ();
 DECAPx10_ASAP7_75t_R FILLER_264_618 ();
 DECAPx10_ASAP7_75t_R FILLER_264_640 ();
 DECAPx10_ASAP7_75t_R FILLER_264_662 ();
 DECAPx10_ASAP7_75t_R FILLER_264_684 ();
 DECAPx6_ASAP7_75t_R FILLER_264_706 ();
 DECAPx2_ASAP7_75t_R FILLER_264_720 ();
 FILLER_ASAP7_75t_R FILLER_264_740 ();
 DECAPx2_ASAP7_75t_R FILLER_264_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_751 ();
 DECAPx6_ASAP7_75t_R FILLER_264_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_772 ();
 FILLER_ASAP7_75t_R FILLER_264_787 ();
 DECAPx1_ASAP7_75t_R FILLER_264_792 ();
 FILLER_ASAP7_75t_R FILLER_264_802 ();
 FILLER_ASAP7_75t_R FILLER_264_810 ();
 DECAPx1_ASAP7_75t_R FILLER_264_815 ();
 DECAPx1_ASAP7_75t_R FILLER_264_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_837 ();
 DECAPx2_ASAP7_75t_R FILLER_264_844 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_264_850 ();
 FILLER_ASAP7_75t_R FILLER_264_867 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_264_872 ();
 DECAPx2_ASAP7_75t_R FILLER_264_881 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_264_887 ();
 DECAPx2_ASAP7_75t_R FILLER_264_904 ();
 DECAPx10_ASAP7_75t_R FILLER_264_916 ();
 DECAPx10_ASAP7_75t_R FILLER_264_938 ();
 DECAPx10_ASAP7_75t_R FILLER_264_960 ();
 DECAPx10_ASAP7_75t_R FILLER_264_982 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1048 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1070 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1158 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1180 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_264_1334 ();
 DECAPx2_ASAP7_75t_R FILLER_264_1356 ();
 FILLER_ASAP7_75t_R FILLER_264_1362 ();
 FILLER_ASAP7_75t_R FILLER_264_1367 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_264_1374 ();
 DECAPx10_ASAP7_75t_R FILLER_265_2 ();
 DECAPx10_ASAP7_75t_R FILLER_265_24 ();
 DECAPx10_ASAP7_75t_R FILLER_265_46 ();
 DECAPx10_ASAP7_75t_R FILLER_265_68 ();
 DECAPx10_ASAP7_75t_R FILLER_265_90 ();
 DECAPx10_ASAP7_75t_R FILLER_265_112 ();
 DECAPx10_ASAP7_75t_R FILLER_265_134 ();
 DECAPx10_ASAP7_75t_R FILLER_265_156 ();
 DECAPx10_ASAP7_75t_R FILLER_265_178 ();
 DECAPx10_ASAP7_75t_R FILLER_265_200 ();
 DECAPx10_ASAP7_75t_R FILLER_265_222 ();
 DECAPx10_ASAP7_75t_R FILLER_265_244 ();
 DECAPx10_ASAP7_75t_R FILLER_265_266 ();
 DECAPx10_ASAP7_75t_R FILLER_265_288 ();
 DECAPx10_ASAP7_75t_R FILLER_265_310 ();
 DECAPx10_ASAP7_75t_R FILLER_265_332 ();
 DECAPx10_ASAP7_75t_R FILLER_265_354 ();
 DECAPx10_ASAP7_75t_R FILLER_265_376 ();
 DECAPx10_ASAP7_75t_R FILLER_265_398 ();
 DECAPx10_ASAP7_75t_R FILLER_265_420 ();
 DECAPx10_ASAP7_75t_R FILLER_265_442 ();
 DECAPx10_ASAP7_75t_R FILLER_265_464 ();
 DECAPx10_ASAP7_75t_R FILLER_265_486 ();
 DECAPx10_ASAP7_75t_R FILLER_265_508 ();
 DECAPx10_ASAP7_75t_R FILLER_265_530 ();
 DECAPx10_ASAP7_75t_R FILLER_265_552 ();
 DECAPx10_ASAP7_75t_R FILLER_265_574 ();
 DECAPx10_ASAP7_75t_R FILLER_265_596 ();
 DECAPx10_ASAP7_75t_R FILLER_265_618 ();
 DECAPx10_ASAP7_75t_R FILLER_265_640 ();
 DECAPx10_ASAP7_75t_R FILLER_265_662 ();
 DECAPx10_ASAP7_75t_R FILLER_265_684 ();
 DECAPx10_ASAP7_75t_R FILLER_265_706 ();
 FILLER_ASAP7_75t_R FILLER_265_728 ();
 DECAPx10_ASAP7_75t_R FILLER_265_736 ();
 DECAPx6_ASAP7_75t_R FILLER_265_758 ();
 DECAPx1_ASAP7_75t_R FILLER_265_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_776 ();
 DECAPx6_ASAP7_75t_R FILLER_265_783 ();
 DECAPx1_ASAP7_75t_R FILLER_265_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_801 ();
 FILLER_ASAP7_75t_R FILLER_265_816 ();
 DECAPx2_ASAP7_75t_R FILLER_265_821 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_265_827 ();
 FILLER_ASAP7_75t_R FILLER_265_833 ();
 DECAPx1_ASAP7_75t_R FILLER_265_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_853 ();
 DECAPx2_ASAP7_75t_R FILLER_265_857 ();
 FILLER_ASAP7_75t_R FILLER_265_863 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_265_868 ();
 DECAPx2_ASAP7_75t_R FILLER_265_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_891 ();
 DECAPx4_ASAP7_75t_R FILLER_265_895 ();
 DECAPx6_ASAP7_75t_R FILLER_265_908 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_265_922 ();
 DECAPx10_ASAP7_75t_R FILLER_265_927 ();
 DECAPx10_ASAP7_75t_R FILLER_265_949 ();
 DECAPx10_ASAP7_75t_R FILLER_265_971 ();
 DECAPx10_ASAP7_75t_R FILLER_265_993 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_265_1323 ();
 DECAPx6_ASAP7_75t_R FILLER_265_1345 ();
 DECAPx2_ASAP7_75t_R FILLER_265_1359 ();
 FILLER_ASAP7_75t_R FILLER_265_1368 ();
 DECAPx1_ASAP7_75t_R FILLER_265_1373 ();
 DECAPx10_ASAP7_75t_R FILLER_266_2 ();
 DECAPx10_ASAP7_75t_R FILLER_266_24 ();
 DECAPx10_ASAP7_75t_R FILLER_266_46 ();
 DECAPx10_ASAP7_75t_R FILLER_266_68 ();
 DECAPx10_ASAP7_75t_R FILLER_266_90 ();
 DECAPx10_ASAP7_75t_R FILLER_266_112 ();
 DECAPx10_ASAP7_75t_R FILLER_266_134 ();
 DECAPx10_ASAP7_75t_R FILLER_266_156 ();
 DECAPx10_ASAP7_75t_R FILLER_266_178 ();
 DECAPx10_ASAP7_75t_R FILLER_266_200 ();
 DECAPx10_ASAP7_75t_R FILLER_266_222 ();
 DECAPx10_ASAP7_75t_R FILLER_266_244 ();
 DECAPx10_ASAP7_75t_R FILLER_266_266 ();
 DECAPx10_ASAP7_75t_R FILLER_266_288 ();
 DECAPx10_ASAP7_75t_R FILLER_266_310 ();
 DECAPx10_ASAP7_75t_R FILLER_266_332 ();
 DECAPx10_ASAP7_75t_R FILLER_266_354 ();
 DECAPx10_ASAP7_75t_R FILLER_266_376 ();
 DECAPx10_ASAP7_75t_R FILLER_266_398 ();
 DECAPx10_ASAP7_75t_R FILLER_266_420 ();
 DECAPx6_ASAP7_75t_R FILLER_266_442 ();
 DECAPx2_ASAP7_75t_R FILLER_266_456 ();
 DECAPx10_ASAP7_75t_R FILLER_266_464 ();
 DECAPx10_ASAP7_75t_R FILLER_266_486 ();
 DECAPx10_ASAP7_75t_R FILLER_266_508 ();
 DECAPx10_ASAP7_75t_R FILLER_266_530 ();
 DECAPx10_ASAP7_75t_R FILLER_266_552 ();
 DECAPx10_ASAP7_75t_R FILLER_266_574 ();
 DECAPx10_ASAP7_75t_R FILLER_266_596 ();
 DECAPx10_ASAP7_75t_R FILLER_266_618 ();
 DECAPx10_ASAP7_75t_R FILLER_266_640 ();
 DECAPx10_ASAP7_75t_R FILLER_266_662 ();
 DECAPx10_ASAP7_75t_R FILLER_266_684 ();
 DECAPx10_ASAP7_75t_R FILLER_266_706 ();
 DECAPx10_ASAP7_75t_R FILLER_266_728 ();
 DECAPx10_ASAP7_75t_R FILLER_266_750 ();
 DECAPx10_ASAP7_75t_R FILLER_266_772 ();
 DECAPx10_ASAP7_75t_R FILLER_266_794 ();
 DECAPx10_ASAP7_75t_R FILLER_266_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_838 ();
 DECAPx10_ASAP7_75t_R FILLER_266_845 ();
 DECAPx2_ASAP7_75t_R FILLER_266_867 ();
 DECAPx10_ASAP7_75t_R FILLER_266_879 ();
 DECAPx10_ASAP7_75t_R FILLER_266_901 ();
 DECAPx10_ASAP7_75t_R FILLER_266_923 ();
 DECAPx10_ASAP7_75t_R FILLER_266_945 ();
 DECAPx10_ASAP7_75t_R FILLER_266_967 ();
 DECAPx10_ASAP7_75t_R FILLER_266_989 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1033 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1055 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_266_1341 ();
 DECAPx2_ASAP7_75t_R FILLER_266_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_1369 ();
 DECAPx1_ASAP7_75t_R FILLER_266_1373 ();
 DECAPx10_ASAP7_75t_R FILLER_267_2 ();
 DECAPx10_ASAP7_75t_R FILLER_267_24 ();
 DECAPx10_ASAP7_75t_R FILLER_267_46 ();
 DECAPx10_ASAP7_75t_R FILLER_267_68 ();
 DECAPx10_ASAP7_75t_R FILLER_267_90 ();
 DECAPx10_ASAP7_75t_R FILLER_267_112 ();
 DECAPx10_ASAP7_75t_R FILLER_267_134 ();
 DECAPx10_ASAP7_75t_R FILLER_267_156 ();
 DECAPx10_ASAP7_75t_R FILLER_267_178 ();
 DECAPx10_ASAP7_75t_R FILLER_267_200 ();
 DECAPx10_ASAP7_75t_R FILLER_267_222 ();
 DECAPx10_ASAP7_75t_R FILLER_267_244 ();
 DECAPx10_ASAP7_75t_R FILLER_267_266 ();
 DECAPx10_ASAP7_75t_R FILLER_267_288 ();
 DECAPx10_ASAP7_75t_R FILLER_267_310 ();
 DECAPx10_ASAP7_75t_R FILLER_267_332 ();
 DECAPx10_ASAP7_75t_R FILLER_267_354 ();
 DECAPx10_ASAP7_75t_R FILLER_267_376 ();
 DECAPx10_ASAP7_75t_R FILLER_267_398 ();
 DECAPx10_ASAP7_75t_R FILLER_267_420 ();
 DECAPx10_ASAP7_75t_R FILLER_267_442 ();
 DECAPx10_ASAP7_75t_R FILLER_267_464 ();
 DECAPx10_ASAP7_75t_R FILLER_267_486 ();
 DECAPx10_ASAP7_75t_R FILLER_267_508 ();
 DECAPx10_ASAP7_75t_R FILLER_267_530 ();
 DECAPx10_ASAP7_75t_R FILLER_267_552 ();
 DECAPx10_ASAP7_75t_R FILLER_267_574 ();
 DECAPx10_ASAP7_75t_R FILLER_267_596 ();
 DECAPx10_ASAP7_75t_R FILLER_267_618 ();
 DECAPx10_ASAP7_75t_R FILLER_267_640 ();
 DECAPx10_ASAP7_75t_R FILLER_267_662 ();
 DECAPx10_ASAP7_75t_R FILLER_267_684 ();
 DECAPx10_ASAP7_75t_R FILLER_267_706 ();
 DECAPx10_ASAP7_75t_R FILLER_267_728 ();
 DECAPx10_ASAP7_75t_R FILLER_267_750 ();
 DECAPx10_ASAP7_75t_R FILLER_267_772 ();
 DECAPx10_ASAP7_75t_R FILLER_267_794 ();
 DECAPx10_ASAP7_75t_R FILLER_267_816 ();
 DECAPx10_ASAP7_75t_R FILLER_267_838 ();
 DECAPx10_ASAP7_75t_R FILLER_267_860 ();
 DECAPx10_ASAP7_75t_R FILLER_267_882 ();
 DECAPx6_ASAP7_75t_R FILLER_267_904 ();
 DECAPx2_ASAP7_75t_R FILLER_267_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_924 ();
 DECAPx10_ASAP7_75t_R FILLER_267_927 ();
 DECAPx10_ASAP7_75t_R FILLER_267_949 ();
 DECAPx10_ASAP7_75t_R FILLER_267_971 ();
 DECAPx10_ASAP7_75t_R FILLER_267_993 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_267_1345 ();
 DECAPx1_ASAP7_75t_R FILLER_267_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_1371 ();
 FILLER_ASAP7_75t_R FILLER_267_1375 ();
 DECAPx10_ASAP7_75t_R FILLER_268_2 ();
 DECAPx10_ASAP7_75t_R FILLER_268_24 ();
 DECAPx10_ASAP7_75t_R FILLER_268_46 ();
 DECAPx10_ASAP7_75t_R FILLER_268_68 ();
 DECAPx10_ASAP7_75t_R FILLER_268_90 ();
 DECAPx10_ASAP7_75t_R FILLER_268_112 ();
 DECAPx10_ASAP7_75t_R FILLER_268_134 ();
 DECAPx10_ASAP7_75t_R FILLER_268_156 ();
 DECAPx10_ASAP7_75t_R FILLER_268_178 ();
 DECAPx10_ASAP7_75t_R FILLER_268_200 ();
 DECAPx10_ASAP7_75t_R FILLER_268_222 ();
 DECAPx10_ASAP7_75t_R FILLER_268_244 ();
 DECAPx10_ASAP7_75t_R FILLER_268_266 ();
 DECAPx10_ASAP7_75t_R FILLER_268_288 ();
 DECAPx10_ASAP7_75t_R FILLER_268_310 ();
 DECAPx10_ASAP7_75t_R FILLER_268_332 ();
 DECAPx10_ASAP7_75t_R FILLER_268_354 ();
 DECAPx10_ASAP7_75t_R FILLER_268_376 ();
 DECAPx10_ASAP7_75t_R FILLER_268_398 ();
 DECAPx10_ASAP7_75t_R FILLER_268_420 ();
 DECAPx6_ASAP7_75t_R FILLER_268_442 ();
 DECAPx2_ASAP7_75t_R FILLER_268_456 ();
 DECAPx10_ASAP7_75t_R FILLER_268_464 ();
 DECAPx10_ASAP7_75t_R FILLER_268_486 ();
 DECAPx10_ASAP7_75t_R FILLER_268_508 ();
 DECAPx10_ASAP7_75t_R FILLER_268_530 ();
 DECAPx10_ASAP7_75t_R FILLER_268_552 ();
 DECAPx10_ASAP7_75t_R FILLER_268_574 ();
 DECAPx10_ASAP7_75t_R FILLER_268_596 ();
 DECAPx10_ASAP7_75t_R FILLER_268_618 ();
 DECAPx10_ASAP7_75t_R FILLER_268_640 ();
 DECAPx10_ASAP7_75t_R FILLER_268_662 ();
 DECAPx10_ASAP7_75t_R FILLER_268_684 ();
 DECAPx10_ASAP7_75t_R FILLER_268_706 ();
 DECAPx10_ASAP7_75t_R FILLER_268_728 ();
 DECAPx10_ASAP7_75t_R FILLER_268_750 ();
 DECAPx10_ASAP7_75t_R FILLER_268_772 ();
 DECAPx10_ASAP7_75t_R FILLER_268_794 ();
 DECAPx10_ASAP7_75t_R FILLER_268_816 ();
 DECAPx10_ASAP7_75t_R FILLER_268_838 ();
 DECAPx10_ASAP7_75t_R FILLER_268_860 ();
 DECAPx10_ASAP7_75t_R FILLER_268_882 ();
 DECAPx10_ASAP7_75t_R FILLER_268_904 ();
 DECAPx10_ASAP7_75t_R FILLER_268_926 ();
 DECAPx10_ASAP7_75t_R FILLER_268_948 ();
 DECAPx10_ASAP7_75t_R FILLER_268_970 ();
 DECAPx10_ASAP7_75t_R FILLER_268_992 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_268_1344 ();
 DECAPx4_ASAP7_75t_R FILLER_268_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_269_2 ();
 DECAPx10_ASAP7_75t_R FILLER_269_24 ();
 DECAPx10_ASAP7_75t_R FILLER_269_46 ();
 DECAPx10_ASAP7_75t_R FILLER_269_68 ();
 DECAPx10_ASAP7_75t_R FILLER_269_90 ();
 DECAPx10_ASAP7_75t_R FILLER_269_112 ();
 DECAPx10_ASAP7_75t_R FILLER_269_134 ();
 DECAPx10_ASAP7_75t_R FILLER_269_156 ();
 DECAPx10_ASAP7_75t_R FILLER_269_178 ();
 DECAPx10_ASAP7_75t_R FILLER_269_200 ();
 DECAPx10_ASAP7_75t_R FILLER_269_222 ();
 DECAPx10_ASAP7_75t_R FILLER_269_244 ();
 DECAPx10_ASAP7_75t_R FILLER_269_266 ();
 DECAPx10_ASAP7_75t_R FILLER_269_288 ();
 DECAPx10_ASAP7_75t_R FILLER_269_310 ();
 DECAPx10_ASAP7_75t_R FILLER_269_332 ();
 DECAPx10_ASAP7_75t_R FILLER_269_354 ();
 DECAPx10_ASAP7_75t_R FILLER_269_376 ();
 DECAPx10_ASAP7_75t_R FILLER_269_398 ();
 DECAPx10_ASAP7_75t_R FILLER_269_420 ();
 DECAPx10_ASAP7_75t_R FILLER_269_442 ();
 DECAPx10_ASAP7_75t_R FILLER_269_464 ();
 DECAPx10_ASAP7_75t_R FILLER_269_486 ();
 DECAPx10_ASAP7_75t_R FILLER_269_508 ();
 DECAPx10_ASAP7_75t_R FILLER_269_530 ();
 DECAPx10_ASAP7_75t_R FILLER_269_552 ();
 DECAPx10_ASAP7_75t_R FILLER_269_574 ();
 DECAPx10_ASAP7_75t_R FILLER_269_596 ();
 DECAPx10_ASAP7_75t_R FILLER_269_618 ();
 DECAPx10_ASAP7_75t_R FILLER_269_640 ();
 DECAPx10_ASAP7_75t_R FILLER_269_662 ();
 DECAPx10_ASAP7_75t_R FILLER_269_684 ();
 DECAPx10_ASAP7_75t_R FILLER_269_706 ();
 DECAPx10_ASAP7_75t_R FILLER_269_728 ();
 DECAPx10_ASAP7_75t_R FILLER_269_750 ();
 DECAPx10_ASAP7_75t_R FILLER_269_772 ();
 DECAPx10_ASAP7_75t_R FILLER_269_794 ();
 DECAPx10_ASAP7_75t_R FILLER_269_816 ();
 DECAPx10_ASAP7_75t_R FILLER_269_838 ();
 DECAPx10_ASAP7_75t_R FILLER_269_860 ();
 DECAPx10_ASAP7_75t_R FILLER_269_882 ();
 DECAPx6_ASAP7_75t_R FILLER_269_904 ();
 DECAPx2_ASAP7_75t_R FILLER_269_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_924 ();
 DECAPx10_ASAP7_75t_R FILLER_269_927 ();
 DECAPx10_ASAP7_75t_R FILLER_269_949 ();
 DECAPx10_ASAP7_75t_R FILLER_269_971 ();
 DECAPx10_ASAP7_75t_R FILLER_269_993 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_269_1345 ();
 DECAPx4_ASAP7_75t_R FILLER_269_1367 ();
 DECAPx10_ASAP7_75t_R FILLER_270_2 ();
 DECAPx10_ASAP7_75t_R FILLER_270_24 ();
 DECAPx10_ASAP7_75t_R FILLER_270_46 ();
 DECAPx10_ASAP7_75t_R FILLER_270_68 ();
 DECAPx10_ASAP7_75t_R FILLER_270_90 ();
 DECAPx10_ASAP7_75t_R FILLER_270_112 ();
 DECAPx10_ASAP7_75t_R FILLER_270_134 ();
 DECAPx10_ASAP7_75t_R FILLER_270_156 ();
 DECAPx10_ASAP7_75t_R FILLER_270_178 ();
 DECAPx10_ASAP7_75t_R FILLER_270_200 ();
 DECAPx10_ASAP7_75t_R FILLER_270_222 ();
 DECAPx10_ASAP7_75t_R FILLER_270_244 ();
 DECAPx10_ASAP7_75t_R FILLER_270_266 ();
 DECAPx10_ASAP7_75t_R FILLER_270_288 ();
 DECAPx10_ASAP7_75t_R FILLER_270_310 ();
 DECAPx10_ASAP7_75t_R FILLER_270_332 ();
 DECAPx10_ASAP7_75t_R FILLER_270_354 ();
 DECAPx10_ASAP7_75t_R FILLER_270_376 ();
 DECAPx10_ASAP7_75t_R FILLER_270_398 ();
 DECAPx10_ASAP7_75t_R FILLER_270_420 ();
 DECAPx6_ASAP7_75t_R FILLER_270_442 ();
 DECAPx2_ASAP7_75t_R FILLER_270_456 ();
 DECAPx10_ASAP7_75t_R FILLER_270_464 ();
 DECAPx10_ASAP7_75t_R FILLER_270_486 ();
 DECAPx10_ASAP7_75t_R FILLER_270_508 ();
 DECAPx10_ASAP7_75t_R FILLER_270_530 ();
 DECAPx10_ASAP7_75t_R FILLER_270_552 ();
 DECAPx10_ASAP7_75t_R FILLER_270_574 ();
 DECAPx10_ASAP7_75t_R FILLER_270_596 ();
 DECAPx10_ASAP7_75t_R FILLER_270_618 ();
 DECAPx10_ASAP7_75t_R FILLER_270_640 ();
 DECAPx10_ASAP7_75t_R FILLER_270_662 ();
 DECAPx10_ASAP7_75t_R FILLER_270_684 ();
 DECAPx10_ASAP7_75t_R FILLER_270_706 ();
 DECAPx10_ASAP7_75t_R FILLER_270_728 ();
 DECAPx10_ASAP7_75t_R FILLER_270_750 ();
 DECAPx10_ASAP7_75t_R FILLER_270_772 ();
 DECAPx10_ASAP7_75t_R FILLER_270_794 ();
 DECAPx10_ASAP7_75t_R FILLER_270_816 ();
 DECAPx10_ASAP7_75t_R FILLER_270_838 ();
 DECAPx10_ASAP7_75t_R FILLER_270_860 ();
 DECAPx10_ASAP7_75t_R FILLER_270_882 ();
 DECAPx10_ASAP7_75t_R FILLER_270_904 ();
 DECAPx10_ASAP7_75t_R FILLER_270_926 ();
 DECAPx10_ASAP7_75t_R FILLER_270_948 ();
 DECAPx10_ASAP7_75t_R FILLER_270_970 ();
 DECAPx10_ASAP7_75t_R FILLER_270_992 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_270_1344 ();
 DECAPx4_ASAP7_75t_R FILLER_270_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_271_2 ();
 DECAPx10_ASAP7_75t_R FILLER_271_24 ();
 DECAPx10_ASAP7_75t_R FILLER_271_46 ();
 DECAPx10_ASAP7_75t_R FILLER_271_68 ();
 DECAPx10_ASAP7_75t_R FILLER_271_90 ();
 DECAPx10_ASAP7_75t_R FILLER_271_112 ();
 DECAPx10_ASAP7_75t_R FILLER_271_134 ();
 DECAPx10_ASAP7_75t_R FILLER_271_156 ();
 DECAPx10_ASAP7_75t_R FILLER_271_178 ();
 DECAPx10_ASAP7_75t_R FILLER_271_200 ();
 DECAPx10_ASAP7_75t_R FILLER_271_222 ();
 DECAPx10_ASAP7_75t_R FILLER_271_244 ();
 DECAPx10_ASAP7_75t_R FILLER_271_266 ();
 DECAPx10_ASAP7_75t_R FILLER_271_288 ();
 DECAPx10_ASAP7_75t_R FILLER_271_310 ();
 DECAPx10_ASAP7_75t_R FILLER_271_332 ();
 DECAPx10_ASAP7_75t_R FILLER_271_354 ();
 DECAPx10_ASAP7_75t_R FILLER_271_376 ();
 DECAPx10_ASAP7_75t_R FILLER_271_398 ();
 DECAPx10_ASAP7_75t_R FILLER_271_420 ();
 DECAPx10_ASAP7_75t_R FILLER_271_442 ();
 DECAPx10_ASAP7_75t_R FILLER_271_464 ();
 DECAPx10_ASAP7_75t_R FILLER_271_486 ();
 DECAPx10_ASAP7_75t_R FILLER_271_508 ();
 DECAPx10_ASAP7_75t_R FILLER_271_530 ();
 DECAPx10_ASAP7_75t_R FILLER_271_552 ();
 DECAPx10_ASAP7_75t_R FILLER_271_574 ();
 DECAPx10_ASAP7_75t_R FILLER_271_596 ();
 DECAPx10_ASAP7_75t_R FILLER_271_618 ();
 DECAPx10_ASAP7_75t_R FILLER_271_640 ();
 DECAPx10_ASAP7_75t_R FILLER_271_662 ();
 DECAPx10_ASAP7_75t_R FILLER_271_684 ();
 DECAPx10_ASAP7_75t_R FILLER_271_706 ();
 DECAPx10_ASAP7_75t_R FILLER_271_728 ();
 DECAPx10_ASAP7_75t_R FILLER_271_750 ();
 DECAPx10_ASAP7_75t_R FILLER_271_772 ();
 DECAPx10_ASAP7_75t_R FILLER_271_794 ();
 DECAPx10_ASAP7_75t_R FILLER_271_816 ();
 DECAPx10_ASAP7_75t_R FILLER_271_838 ();
 DECAPx10_ASAP7_75t_R FILLER_271_860 ();
 DECAPx10_ASAP7_75t_R FILLER_271_882 ();
 DECAPx6_ASAP7_75t_R FILLER_271_904 ();
 DECAPx2_ASAP7_75t_R FILLER_271_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_924 ();
 DECAPx10_ASAP7_75t_R FILLER_271_927 ();
 DECAPx10_ASAP7_75t_R FILLER_271_949 ();
 DECAPx10_ASAP7_75t_R FILLER_271_971 ();
 DECAPx10_ASAP7_75t_R FILLER_271_993 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_271_1345 ();
 DECAPx4_ASAP7_75t_R FILLER_271_1367 ();
 DECAPx10_ASAP7_75t_R FILLER_272_2 ();
 DECAPx10_ASAP7_75t_R FILLER_272_24 ();
 DECAPx10_ASAP7_75t_R FILLER_272_46 ();
 DECAPx10_ASAP7_75t_R FILLER_272_68 ();
 DECAPx10_ASAP7_75t_R FILLER_272_90 ();
 DECAPx10_ASAP7_75t_R FILLER_272_112 ();
 DECAPx10_ASAP7_75t_R FILLER_272_134 ();
 DECAPx10_ASAP7_75t_R FILLER_272_156 ();
 DECAPx10_ASAP7_75t_R FILLER_272_178 ();
 DECAPx10_ASAP7_75t_R FILLER_272_200 ();
 DECAPx10_ASAP7_75t_R FILLER_272_222 ();
 DECAPx10_ASAP7_75t_R FILLER_272_244 ();
 DECAPx10_ASAP7_75t_R FILLER_272_266 ();
 DECAPx10_ASAP7_75t_R FILLER_272_288 ();
 DECAPx10_ASAP7_75t_R FILLER_272_310 ();
 DECAPx10_ASAP7_75t_R FILLER_272_332 ();
 DECAPx10_ASAP7_75t_R FILLER_272_354 ();
 DECAPx10_ASAP7_75t_R FILLER_272_376 ();
 DECAPx10_ASAP7_75t_R FILLER_272_398 ();
 DECAPx10_ASAP7_75t_R FILLER_272_420 ();
 DECAPx6_ASAP7_75t_R FILLER_272_442 ();
 DECAPx2_ASAP7_75t_R FILLER_272_456 ();
 DECAPx10_ASAP7_75t_R FILLER_272_464 ();
 DECAPx10_ASAP7_75t_R FILLER_272_486 ();
 DECAPx10_ASAP7_75t_R FILLER_272_508 ();
 DECAPx10_ASAP7_75t_R FILLER_272_530 ();
 DECAPx10_ASAP7_75t_R FILLER_272_552 ();
 DECAPx10_ASAP7_75t_R FILLER_272_574 ();
 DECAPx10_ASAP7_75t_R FILLER_272_596 ();
 DECAPx10_ASAP7_75t_R FILLER_272_618 ();
 DECAPx10_ASAP7_75t_R FILLER_272_640 ();
 DECAPx10_ASAP7_75t_R FILLER_272_662 ();
 DECAPx10_ASAP7_75t_R FILLER_272_684 ();
 DECAPx10_ASAP7_75t_R FILLER_272_706 ();
 DECAPx10_ASAP7_75t_R FILLER_272_728 ();
 DECAPx10_ASAP7_75t_R FILLER_272_750 ();
 DECAPx10_ASAP7_75t_R FILLER_272_772 ();
 DECAPx10_ASAP7_75t_R FILLER_272_794 ();
 DECAPx10_ASAP7_75t_R FILLER_272_816 ();
 DECAPx10_ASAP7_75t_R FILLER_272_838 ();
 DECAPx10_ASAP7_75t_R FILLER_272_860 ();
 DECAPx10_ASAP7_75t_R FILLER_272_882 ();
 DECAPx10_ASAP7_75t_R FILLER_272_904 ();
 DECAPx10_ASAP7_75t_R FILLER_272_926 ();
 DECAPx10_ASAP7_75t_R FILLER_272_948 ();
 DECAPx10_ASAP7_75t_R FILLER_272_970 ();
 DECAPx10_ASAP7_75t_R FILLER_272_992 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_272_1344 ();
 DECAPx4_ASAP7_75t_R FILLER_272_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_273_2 ();
 DECAPx10_ASAP7_75t_R FILLER_273_24 ();
 DECAPx10_ASAP7_75t_R FILLER_273_46 ();
 DECAPx10_ASAP7_75t_R FILLER_273_68 ();
 DECAPx10_ASAP7_75t_R FILLER_273_90 ();
 DECAPx10_ASAP7_75t_R FILLER_273_112 ();
 DECAPx10_ASAP7_75t_R FILLER_273_134 ();
 DECAPx10_ASAP7_75t_R FILLER_273_156 ();
 DECAPx10_ASAP7_75t_R FILLER_273_178 ();
 DECAPx10_ASAP7_75t_R FILLER_273_200 ();
 DECAPx10_ASAP7_75t_R FILLER_273_222 ();
 DECAPx10_ASAP7_75t_R FILLER_273_244 ();
 DECAPx10_ASAP7_75t_R FILLER_273_266 ();
 DECAPx10_ASAP7_75t_R FILLER_273_288 ();
 DECAPx10_ASAP7_75t_R FILLER_273_310 ();
 DECAPx10_ASAP7_75t_R FILLER_273_332 ();
 DECAPx10_ASAP7_75t_R FILLER_273_354 ();
 DECAPx10_ASAP7_75t_R FILLER_273_376 ();
 DECAPx10_ASAP7_75t_R FILLER_273_398 ();
 DECAPx10_ASAP7_75t_R FILLER_273_420 ();
 DECAPx10_ASAP7_75t_R FILLER_273_442 ();
 DECAPx10_ASAP7_75t_R FILLER_273_464 ();
 DECAPx10_ASAP7_75t_R FILLER_273_486 ();
 DECAPx10_ASAP7_75t_R FILLER_273_508 ();
 DECAPx10_ASAP7_75t_R FILLER_273_530 ();
 DECAPx10_ASAP7_75t_R FILLER_273_552 ();
 DECAPx10_ASAP7_75t_R FILLER_273_574 ();
 DECAPx10_ASAP7_75t_R FILLER_273_596 ();
 DECAPx2_ASAP7_75t_R FILLER_273_618 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_273_624 ();
 DECAPx4_ASAP7_75t_R FILLER_273_632 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_273_642 ();
 FILLER_ASAP7_75t_R FILLER_273_650 ();
 DECAPx4_ASAP7_75t_R FILLER_273_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_667 ();
 DECAPx10_ASAP7_75t_R FILLER_273_673 ();
 DECAPx10_ASAP7_75t_R FILLER_273_695 ();
 DECAPx10_ASAP7_75t_R FILLER_273_717 ();
 DECAPx10_ASAP7_75t_R FILLER_273_739 ();
 DECAPx10_ASAP7_75t_R FILLER_273_761 ();
 DECAPx10_ASAP7_75t_R FILLER_273_783 ();
 DECAPx10_ASAP7_75t_R FILLER_273_805 ();
 DECAPx10_ASAP7_75t_R FILLER_273_827 ();
 DECAPx10_ASAP7_75t_R FILLER_273_849 ();
 DECAPx10_ASAP7_75t_R FILLER_273_871 ();
 DECAPx10_ASAP7_75t_R FILLER_273_893 ();
 DECAPx4_ASAP7_75t_R FILLER_273_915 ();
 DECAPx10_ASAP7_75t_R FILLER_273_927 ();
 DECAPx10_ASAP7_75t_R FILLER_273_949 ();
 DECAPx10_ASAP7_75t_R FILLER_273_971 ();
 DECAPx10_ASAP7_75t_R FILLER_273_993 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_273_1345 ();
 DECAPx4_ASAP7_75t_R FILLER_273_1367 ();
 DECAPx10_ASAP7_75t_R FILLER_274_2 ();
 DECAPx10_ASAP7_75t_R FILLER_274_24 ();
 DECAPx10_ASAP7_75t_R FILLER_274_46 ();
 DECAPx10_ASAP7_75t_R FILLER_274_68 ();
 DECAPx10_ASAP7_75t_R FILLER_274_90 ();
 DECAPx10_ASAP7_75t_R FILLER_274_112 ();
 DECAPx10_ASAP7_75t_R FILLER_274_134 ();
 DECAPx10_ASAP7_75t_R FILLER_274_156 ();
 DECAPx10_ASAP7_75t_R FILLER_274_178 ();
 DECAPx10_ASAP7_75t_R FILLER_274_200 ();
 DECAPx10_ASAP7_75t_R FILLER_274_222 ();
 DECAPx10_ASAP7_75t_R FILLER_274_244 ();
 DECAPx10_ASAP7_75t_R FILLER_274_266 ();
 DECAPx10_ASAP7_75t_R FILLER_274_288 ();
 DECAPx10_ASAP7_75t_R FILLER_274_310 ();
 DECAPx10_ASAP7_75t_R FILLER_274_332 ();
 DECAPx10_ASAP7_75t_R FILLER_274_354 ();
 DECAPx10_ASAP7_75t_R FILLER_274_376 ();
 DECAPx10_ASAP7_75t_R FILLER_274_398 ();
 DECAPx10_ASAP7_75t_R FILLER_274_420 ();
 DECAPx6_ASAP7_75t_R FILLER_274_442 ();
 DECAPx2_ASAP7_75t_R FILLER_274_456 ();
 DECAPx10_ASAP7_75t_R FILLER_274_464 ();
 DECAPx10_ASAP7_75t_R FILLER_274_486 ();
 DECAPx10_ASAP7_75t_R FILLER_274_508 ();
 DECAPx10_ASAP7_75t_R FILLER_274_530 ();
 DECAPx10_ASAP7_75t_R FILLER_274_552 ();
 DECAPx10_ASAP7_75t_R FILLER_274_574 ();
 DECAPx10_ASAP7_75t_R FILLER_274_596 ();
 DECAPx2_ASAP7_75t_R FILLER_274_618 ();
 FILLER_ASAP7_75t_R FILLER_274_629 ();
 DECAPx2_ASAP7_75t_R FILLER_274_636 ();
 FILLER_ASAP7_75t_R FILLER_274_642 ();
 FILLER_ASAP7_75t_R FILLER_274_649 ();
 FILLER_ASAP7_75t_R FILLER_274_656 ();
 FILLER_ASAP7_75t_R FILLER_274_663 ();
 FILLER_ASAP7_75t_R FILLER_274_670 ();
 FILLER_ASAP7_75t_R FILLER_274_677 ();
 DECAPx10_ASAP7_75t_R FILLER_274_684 ();
 DECAPx10_ASAP7_75t_R FILLER_274_706 ();
 DECAPx6_ASAP7_75t_R FILLER_274_728 ();
 FILLER_ASAP7_75t_R FILLER_274_742 ();
 DECAPx6_ASAP7_75t_R FILLER_274_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_763 ();
 DECAPx10_ASAP7_75t_R FILLER_274_769 ();
 DECAPx10_ASAP7_75t_R FILLER_274_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_813 ();
 FILLER_ASAP7_75t_R FILLER_274_819 ();
 DECAPx2_ASAP7_75t_R FILLER_274_826 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_274_832 ();
 FILLER_ASAP7_75t_R FILLER_274_840 ();
 DECAPx10_ASAP7_75t_R FILLER_274_847 ();
 DECAPx10_ASAP7_75t_R FILLER_274_874 ();
 DECAPx10_ASAP7_75t_R FILLER_274_896 ();
 DECAPx2_ASAP7_75t_R FILLER_274_918 ();
 DECAPx10_ASAP7_75t_R FILLER_274_926 ();
 DECAPx2_ASAP7_75t_R FILLER_274_948 ();
 FILLER_ASAP7_75t_R FILLER_274_954 ();
 DECAPx10_ASAP7_75t_R FILLER_274_961 ();
 DECAPx10_ASAP7_75t_R FILLER_274_983 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1027 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1071 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1137 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1159 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_274_1335 ();
 DECAPx6_ASAP7_75t_R FILLER_274_1357 ();
 DECAPx2_ASAP7_75t_R FILLER_274_1371 ();
 assign alert_major_o = net450;
endmodule
